//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 1 1 0 1 0 0 1 0 0 0 1 1 1 1 0 0 0 1 0 0 0 0 0 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n791, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n876, new_n877,
    new_n879, new_n880, new_n881, new_n882, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980;
  INV_X1    g000(.A(KEYINPUT80), .ZN(new_n202));
  INV_X1    g001(.A(G141gat), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G148gat), .ZN(new_n204));
  INV_X1    g003(.A(G148gat), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT79), .B1(new_n205), .B2(G141gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT79), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n207), .A2(new_n203), .A3(G148gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n205), .A2(KEYINPUT80), .A3(G141gat), .ZN(new_n209));
  NAND4_X1  g008(.A1(new_n204), .A2(new_n206), .A3(new_n208), .A4(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT2), .ZN(new_n211));
  INV_X1    g010(.A(G155gat), .ZN(new_n212));
  INV_X1    g011(.A(G162gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n214), .B1(new_n212), .B2(new_n213), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n210), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n203), .A2(G148gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n205), .A2(G141gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n211), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  XOR2_X1   g019(.A(G155gat), .B(G162gat), .Z(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n216), .A2(new_n217), .A3(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT78), .B(KEYINPUT29), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT76), .ZN(new_n227));
  AND2_X1   g026(.A1(G197gat), .A2(G204gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(G197gat), .A2(G204gat), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT73), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G197gat), .ZN(new_n231));
  INV_X1    g030(.A(G204gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT73), .ZN(new_n234));
  NAND2_X1  g033(.A1(G197gat), .A2(G204gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n230), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G211gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(KEYINPUT75), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT75), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G211gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n239), .A2(new_n241), .A3(G218gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT74), .B(KEYINPUT22), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(G211gat), .B(G218gat), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n237), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n245), .B1(new_n237), .B2(new_n244), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n227), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n237), .A2(new_n244), .ZN(new_n249));
  INV_X1    g048(.A(new_n245), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n237), .A2(new_n244), .A3(new_n245), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n251), .A2(KEYINPUT76), .A3(new_n252), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n248), .A2(new_n253), .A3(KEYINPUT77), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT77), .B1(new_n248), .B2(new_n253), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n226), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n216), .A2(new_n222), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT29), .B1(new_n251), .B2(new_n252), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n257), .B1(new_n258), .B2(KEYINPUT3), .ZN(new_n259));
  NAND2_X1  g058(.A1(G228gat), .A2(G233gat), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n256), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n224), .B1(new_n251), .B2(new_n252), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n257), .B1(new_n263), .B2(KEYINPUT3), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n248), .A2(new_n253), .A3(new_n226), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT87), .B1(new_n266), .B2(new_n260), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT87), .ZN(new_n268));
  AOI211_X1 g067(.A(new_n268), .B(new_n261), .C1(new_n264), .C2(new_n265), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n262), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(G22gat), .ZN(new_n271));
  INV_X1    g070(.A(G22gat), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n262), .B(new_n272), .C1(new_n267), .C2(new_n269), .ZN(new_n273));
  XOR2_X1   g072(.A(G78gat), .B(G106gat), .Z(new_n274));
  XNOR2_X1  g073(.A(KEYINPUT31), .B(G50gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n271), .A2(KEYINPUT88), .A3(new_n273), .A4(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT88), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n273), .A2(new_n279), .ZN(new_n280));
  AOI22_X1  g079(.A1(new_n280), .A2(new_n276), .B1(new_n271), .B2(new_n273), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  AOI22_X1  g081(.A1(new_n215), .A2(new_n210), .B1(new_n220), .B2(new_n221), .ZN(new_n283));
  INV_X1    g082(.A(G120gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(G113gat), .ZN(new_n285));
  INV_X1    g084(.A(G113gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(G120gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G127gat), .B(G134gat), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT1), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G113gat), .B(G120gat), .ZN(new_n292));
  INV_X1    g091(.A(G134gat), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n293), .A2(G127gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(G127gat), .ZN(new_n295));
  OAI22_X1  g094(.A1(new_n292), .A2(KEYINPUT1), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n283), .A2(KEYINPUT4), .A3(new_n291), .A4(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT68), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n289), .B1(new_n290), .B2(new_n288), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n296), .A2(new_n291), .A3(KEYINPUT68), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n257), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n297), .B1(new_n303), .B2(KEYINPUT4), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n296), .A2(new_n291), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n305), .A2(new_n306), .A3(new_n223), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT81), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n305), .A2(KEYINPUT81), .A3(new_n306), .A4(new_n223), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n304), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(G225gat), .A2(G233gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(KEYINPUT89), .B(KEYINPUT39), .ZN(new_n313));
  OR3_X1    g112(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n315), .B(G29gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(G57gat), .B(G85gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n316), .B(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(KEYINPUT84), .B(G1gat), .ZN(new_n319));
  XOR2_X1   g118(.A(new_n318), .B(new_n319), .Z(new_n320));
  NAND3_X1  g119(.A1(new_n283), .A2(new_n291), .A3(new_n296), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n257), .A2(new_n306), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n321), .A2(new_n322), .A3(new_n312), .ZN(new_n323));
  OAI211_X1 g122(.A(KEYINPUT39), .B(new_n323), .C1(new_n311), .C2(new_n312), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n314), .A2(new_n320), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT40), .ZN(new_n326));
  OR2_X1    g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n312), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n328), .B1(new_n309), .B2(new_n310), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT4), .ZN(new_n330));
  OAI21_X1  g129(.A(KEYINPUT82), .B1(new_n303), .B2(new_n330), .ZN(new_n331));
  OR2_X1    g130(.A1(new_n321), .A2(KEYINPUT4), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n296), .A2(new_n291), .A3(KEYINPUT68), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT68), .B1(new_n296), .B2(new_n291), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n283), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT82), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n335), .A2(new_n336), .A3(KEYINPUT4), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n331), .A2(new_n332), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n329), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT5), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n321), .A2(new_n322), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n340), .B1(new_n341), .B2(new_n328), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n340), .B(new_n297), .C1(new_n303), .C2(KEYINPUT4), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n329), .A2(new_n345), .A3(KEYINPUT85), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT85), .B1(new_n329), .B2(new_n345), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n343), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n320), .ZN(new_n349));
  AOI22_X1  g148(.A1(new_n325), .A2(new_n326), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n248), .A2(new_n253), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT77), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n248), .A2(new_n253), .A3(KEYINPUT77), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NOR3_X1   g156(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT23), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(G169gat), .ZN(new_n360));
  INV_X1    g159(.A(G176gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n359), .A2(KEYINPUT66), .A3(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT66), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT23), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT65), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n367), .A2(new_n360), .A3(new_n361), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n366), .B1(new_n368), .B2(new_n356), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n365), .B1(new_n369), .B2(new_n362), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT24), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n371), .A2(G183gat), .A3(G190gat), .ZN(new_n372));
  NOR2_X1   g171(.A1(G169gat), .A2(G176gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(G183gat), .A2(G190gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT24), .ZN(new_n375));
  NOR2_X1   g174(.A1(G183gat), .A2(G190gat), .ZN(new_n376));
  OAI221_X1 g175(.A(new_n372), .B1(new_n373), .B2(KEYINPUT23), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n364), .A2(new_n370), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT25), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n363), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT26), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n383), .B1(new_n357), .B2(new_n358), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT28), .ZN(new_n386));
  OR2_X1    g185(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(KEYINPUT67), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT67), .ZN(new_n390));
  AND2_X1   g189(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n391));
  NOR2_X1   g190(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  AOI211_X1 g192(.A(new_n386), .B(G190gat), .C1(new_n389), .C2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n387), .A2(new_n388), .ZN(new_n395));
  INV_X1    g194(.A(G190gat), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT28), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n374), .B(new_n385), .C1(new_n394), .C2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(KEYINPUT64), .B(G169gat), .ZN(new_n399));
  NOR3_X1   g198(.A1(new_n399), .A2(new_n366), .A3(G176gat), .ZN(new_n400));
  OR2_X1    g199(.A1(new_n362), .A2(KEYINPUT25), .ZN(new_n401));
  NOR3_X1   g200(.A1(new_n400), .A2(new_n377), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n380), .A2(new_n398), .A3(new_n403), .ZN(new_n404));
  AND2_X1   g203(.A1(G226gat), .A2(G233gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n405), .B1(new_n404), .B2(new_n225), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n355), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n389), .A2(new_n393), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n410), .A2(KEYINPUT28), .A3(new_n396), .ZN(new_n411));
  INV_X1    g210(.A(new_n397), .ZN(new_n412));
  AOI22_X1  g211(.A1(new_n411), .A2(new_n412), .B1(new_n384), .B2(new_n382), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n402), .B1(new_n413), .B2(new_n374), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT29), .B1(new_n414), .B2(new_n380), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n406), .B(new_n351), .C1(new_n415), .C2(new_n405), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n409), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT30), .ZN(new_n419));
  XOR2_X1   g218(.A(G8gat), .B(G36gat), .Z(new_n420));
  XNOR2_X1  g219(.A(new_n420), .B(G64gat), .ZN(new_n421));
  INV_X1    g220(.A(G92gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n421), .B(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n418), .A2(new_n419), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n418), .A2(new_n424), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n419), .B1(new_n417), .B2(new_n423), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n327), .A2(new_n350), .A3(new_n425), .A4(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT37), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n254), .A2(new_n255), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n224), .B1(new_n414), .B2(new_n380), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n431), .B(new_n406), .C1(new_n405), .C2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n351), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT29), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n405), .B1(new_n404), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n434), .B1(new_n407), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n430), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  XOR2_X1   g237(.A(KEYINPUT90), .B(KEYINPUT38), .Z(new_n439));
  NOR3_X1   g238(.A1(new_n438), .A2(new_n424), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n409), .A2(new_n416), .A3(new_n430), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT91), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n409), .A2(new_n416), .A3(KEYINPUT91), .A4(new_n430), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n440), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n348), .A2(KEYINPUT6), .A3(new_n349), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n348), .A2(new_n349), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT6), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n343), .B(new_n320), .C1(new_n346), .C2(new_n347), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n446), .A2(new_n447), .A3(new_n451), .ZN(new_n452));
  AOI22_X1  g251(.A1(new_n443), .A2(new_n444), .B1(KEYINPUT37), .B2(new_n417), .ZN(new_n453));
  INV_X1    g252(.A(new_n439), .ZN(new_n454));
  AOI22_X1  g253(.A1(new_n453), .A2(new_n423), .B1(new_n426), .B2(new_n454), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n282), .B(new_n429), .C1(new_n452), .C2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n280), .A2(new_n276), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n271), .A2(new_n273), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n277), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n428), .A2(new_n425), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n450), .A2(KEYINPUT86), .A3(new_n449), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n329), .A2(new_n345), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT85), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n329), .A2(KEYINPUT85), .A3(new_n345), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n320), .B1(new_n467), .B2(new_n343), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n462), .A2(new_n468), .ZN(new_n469));
  AOI221_X4 g268(.A(new_n320), .B1(KEYINPUT86), .B2(new_n449), .C1(new_n467), .C2(new_n343), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n461), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT36), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n301), .A2(new_n302), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n404), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(G227gat), .A2(G233gat), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n380), .A2(new_n398), .A3(new_n473), .A4(new_n403), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT71), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT34), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(G15gat), .B(G43gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n481), .B(G71gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n482), .B(G99gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n475), .A2(new_n477), .ZN(new_n484));
  INV_X1    g283(.A(new_n476), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  XOR2_X1   g285(.A(KEYINPUT69), .B(KEYINPUT33), .Z(new_n487));
  INV_X1    g286(.A(KEYINPUT32), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n483), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n476), .B1(new_n475), .B2(new_n477), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT70), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n483), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(G99gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n482), .B(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT70), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n493), .A2(new_n496), .A3(new_n487), .ZN(new_n497));
  NOR3_X1   g296(.A1(new_n491), .A2(new_n488), .A3(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n480), .B1(new_n490), .B2(new_n498), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n475), .A2(KEYINPUT71), .A3(new_n476), .A4(new_n477), .ZN(new_n500));
  XOR2_X1   g299(.A(new_n500), .B(KEYINPUT72), .Z(new_n501));
  NAND2_X1  g300(.A1(new_n478), .A2(new_n479), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT34), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n497), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n486), .A2(KEYINPUT32), .A3(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n489), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n495), .B1(new_n491), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n504), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n499), .A2(new_n501), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n501), .B1(new_n499), .B2(new_n509), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n472), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n501), .ZN(new_n513));
  INV_X1    g312(.A(new_n509), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n504), .B1(new_n508), .B2(new_n506), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n499), .A2(new_n501), .A3(new_n509), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(KEYINPUT36), .A3(new_n517), .ZN(new_n518));
  AOI22_X1  g317(.A1(new_n460), .A2(new_n471), .B1(new_n512), .B2(new_n518), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n459), .A2(new_n516), .A3(new_n277), .A4(new_n517), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT35), .B1(new_n520), .B2(new_n471), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n510), .A2(new_n511), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n451), .A2(new_n447), .ZN(new_n523));
  XOR2_X1   g322(.A(KEYINPUT92), .B(KEYINPUT35), .Z(new_n524));
  AOI21_X1  g323(.A(new_n524), .B1(new_n428), .B2(new_n425), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n282), .A2(new_n522), .A3(new_n523), .A4(new_n525), .ZN(new_n526));
  AOI22_X1  g325(.A1(new_n456), .A2(new_n519), .B1(new_n521), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT10), .ZN(new_n528));
  NAND2_X1  g327(.A1(G85gat), .A2(G92gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  NAND2_X1  g329(.A1(G99gat), .A2(G106gat), .ZN(new_n531));
  INV_X1    g330(.A(G85gat), .ZN(new_n532));
  AOI22_X1  g331(.A1(KEYINPUT8), .A2(new_n531), .B1(new_n532), .B2(new_n422), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  XOR2_X1   g333(.A(G99gat), .B(G106gat), .Z(new_n535));
  NOR2_X1   g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n534), .A2(new_n535), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n536), .B1(new_n537), .B2(KEYINPUT103), .ZN(new_n538));
  XOR2_X1   g337(.A(G71gat), .B(G78gat), .Z(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT9), .ZN(new_n541));
  INV_X1    g340(.A(G71gat), .ZN(new_n542));
  INV_X1    g341(.A(G78gat), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(G57gat), .B(G64gat), .Z(new_n545));
  NAND3_X1  g344(.A1(new_n540), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n544), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(new_n539), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n538), .B(new_n550), .C1(KEYINPUT103), .C2(new_n535), .ZN(new_n551));
  OR2_X1    g350(.A1(new_n537), .A2(new_n536), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT102), .B1(new_n552), .B2(new_n549), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n549), .B(KEYINPUT102), .C1(new_n537), .C2(new_n536), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n528), .B(new_n551), .C1(new_n553), .C2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n552), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n557), .A2(new_n550), .A3(KEYINPUT10), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(G230gat), .ZN(new_n560));
  INV_X1    g359(.A(G233gat), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n551), .B1(new_n553), .B2(new_n555), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(new_n562), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G120gat), .B(G148gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT104), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(G176gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G204gat), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n567), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n564), .A2(new_n566), .A3(new_n571), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n573), .A2(KEYINPUT105), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(KEYINPUT105), .B1(new_n573), .B2(new_n574), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G43gat), .B(G50gat), .ZN(new_n579));
  INV_X1    g378(.A(G29gat), .ZN(new_n580));
  INV_X1    g379(.A(G36gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n582), .A2(KEYINPUT94), .A3(KEYINPUT14), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(KEYINPUT14), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n583), .B1(new_n584), .B2(KEYINPUT94), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n580), .A2(new_n581), .ZN(new_n586));
  OAI211_X1 g385(.A(KEYINPUT15), .B(new_n579), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n579), .A2(KEYINPUT15), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT95), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n579), .A2(KEYINPUT15), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n590), .A2(new_n584), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n587), .B1(new_n592), .B2(new_n586), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT17), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(G8gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(G15gat), .B(G22gat), .ZN(new_n597));
  OR2_X1    g396(.A1(new_n597), .A2(G1gat), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT96), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n596), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT16), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n597), .B1(new_n601), .B2(G1gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n600), .B(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n587), .B(KEYINPUT17), .C1(new_n592), .C2(new_n586), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n595), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G229gat), .A2(G233gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n604), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT18), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n607), .A2(KEYINPUT18), .A3(new_n608), .A4(new_n609), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n608), .B(KEYINPUT13), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n609), .B(KEYINPUT97), .ZN(new_n616));
  OR3_X1    g415(.A1(new_n593), .A2(KEYINPUT98), .A3(new_n604), .ZN(new_n617));
  OAI21_X1  g416(.A(KEYINPUT98), .B1(new_n593), .B2(new_n604), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n615), .B1(new_n616), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(KEYINPUT93), .B1(new_n614), .B2(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G113gat), .B(G141gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(G197gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT11), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(new_n360), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n625), .B(KEYINPUT12), .Z(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n621), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n615), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n617), .A2(new_n618), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT97), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n609), .B(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n629), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n633), .A2(new_n612), .A3(new_n613), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n634), .A2(KEYINPUT93), .A3(new_n626), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n628), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n578), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n527), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n550), .A2(KEYINPUT21), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n604), .A2(new_n639), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n604), .A2(new_n639), .ZN(new_n641));
  AND2_X1   g440(.A1(new_n550), .A2(KEYINPUT21), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g444(.A(G127gat), .B(G155gat), .Z(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g446(.A(G183gat), .B(G211gat), .Z(new_n648));
  NAND2_X1  g447(.A1(G231gat), .A2(G233gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g449(.A(KEYINPUT99), .B(KEYINPUT100), .Z(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n647), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g452(.A(G190gat), .B(G218gat), .Z(new_n654));
  NOR2_X1   g453(.A1(new_n654), .A2(KEYINPUT101), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n595), .A2(new_n552), .A3(new_n606), .ZN(new_n656));
  NAND3_X1  g455(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n593), .A2(new_n557), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n654), .A2(KEYINPUT101), .ZN(new_n660));
  AND3_X1   g459(.A1(new_n659), .A2(new_n213), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n213), .B1(new_n659), .B2(new_n660), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n655), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n659), .A2(new_n660), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(G162gat), .ZN(new_n665));
  INV_X1    g464(.A(new_n655), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n659), .A2(new_n213), .A3(new_n660), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(G134gat), .ZN(new_n670));
  AND3_X1   g469(.A1(new_n663), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n670), .B1(new_n663), .B2(new_n668), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n653), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n638), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n469), .A2(new_n470), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(G1gat), .ZN(G1324gat));
  INV_X1    g477(.A(KEYINPUT42), .ZN(new_n679));
  INV_X1    g478(.A(new_n461), .ZN(new_n680));
  NOR2_X1   g479(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n601), .A2(new_n596), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n675), .A2(new_n680), .A3(new_n682), .A4(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n638), .A2(new_n674), .ZN(new_n686));
  OAI21_X1  g485(.A(G8gat), .B1(new_n686), .B2(new_n461), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n679), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n686), .A2(new_n461), .A3(new_n683), .ZN(new_n689));
  AOI21_X1  g488(.A(KEYINPUT42), .B1(new_n689), .B2(new_n682), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT106), .ZN(G1325gat));
  AOI21_X1  g491(.A(G15gat), .B1(new_n675), .B2(new_n522), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n512), .A2(new_n518), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT107), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(G15gat), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n697), .B(KEYINPUT108), .Z(new_n698));
  AOI21_X1  g497(.A(new_n693), .B1(new_n698), .B2(new_n675), .ZN(G1326gat));
  NOR2_X1   g498(.A1(new_n686), .A2(new_n282), .ZN(new_n700));
  XOR2_X1   g499(.A(KEYINPUT43), .B(G22gat), .Z(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1327gat));
  NAND2_X1  g501(.A1(new_n663), .A2(new_n668), .ZN(new_n703));
  INV_X1    g502(.A(new_n670), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n663), .A2(new_n668), .A3(new_n670), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(KEYINPUT44), .B1(new_n527), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n521), .A2(new_n526), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n471), .A2(new_n460), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n456), .A2(new_n694), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n712), .A2(new_n713), .A3(new_n673), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n708), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n653), .ZN(new_n716));
  OAI21_X1  g515(.A(KEYINPUT110), .B1(new_n716), .B2(new_n637), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT110), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n653), .A2(new_n718), .A3(new_n578), .A4(new_n636), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n715), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n676), .ZN(new_n723));
  OAI21_X1  g522(.A(G29gat), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n712), .A2(new_n673), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n725), .A2(new_n716), .A3(new_n637), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n726), .A2(new_n580), .A3(new_n676), .ZN(new_n727));
  OR2_X1    g526(.A1(new_n727), .A2(KEYINPUT109), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT45), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(KEYINPUT109), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n729), .B1(new_n728), .B2(new_n730), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n724), .B1(new_n731), .B2(new_n732), .ZN(G1328gat));
  NAND3_X1  g532(.A1(new_n726), .A2(new_n581), .A3(new_n680), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n734), .A2(KEYINPUT46), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT111), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(KEYINPUT46), .ZN(new_n737));
  OAI21_X1  g536(.A(G36gat), .B1(new_n722), .B2(new_n461), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(G1329gat));
  INV_X1    g538(.A(KEYINPUT47), .ZN(new_n740));
  INV_X1    g539(.A(new_n694), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n713), .B1(new_n712), .B2(new_n673), .ZN(new_n742));
  AOI211_X1 g541(.A(KEYINPUT44), .B(new_n707), .C1(new_n709), .C2(new_n711), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n741), .B(new_n721), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT112), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT112), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n715), .A2(new_n746), .A3(new_n741), .A4(new_n721), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n745), .A2(G43gat), .A3(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n716), .A2(new_n637), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n522), .ZN(new_n751));
  NOR4_X1   g550(.A1(new_n725), .A2(new_n750), .A3(G43gat), .A4(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n740), .B1(new_n748), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n715), .A2(new_n696), .A3(new_n721), .ZN(new_n755));
  AOI211_X1 g554(.A(KEYINPUT47), .B(new_n752), .C1(new_n755), .C2(G43gat), .ZN(new_n756));
  OAI21_X1  g555(.A(KEYINPUT113), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT113), .ZN(new_n758));
  INV_X1    g557(.A(new_n756), .ZN(new_n759));
  INV_X1    g558(.A(G43gat), .ZN(new_n760));
  AOI211_X1 g559(.A(new_n694), .B(new_n720), .C1(new_n708), .C2(new_n714), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n760), .B1(new_n761), .B2(new_n746), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n752), .B1(new_n762), .B2(new_n745), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n758), .B(new_n759), .C1(new_n763), .C2(new_n740), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n757), .A2(new_n764), .ZN(G1330gat));
  OAI21_X1  g564(.A(G50gat), .B1(new_n722), .B2(new_n282), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT114), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT48), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(G50gat), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n726), .A2(new_n769), .A3(new_n460), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n768), .B(new_n771), .ZN(G1331gat));
  INV_X1    g571(.A(new_n636), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n674), .A2(new_n773), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n527), .A2(new_n774), .A3(new_n578), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n676), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n680), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n778), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n779));
  XOR2_X1   g578(.A(KEYINPUT49), .B(G64gat), .Z(new_n780));
  OAI21_X1  g579(.A(new_n779), .B1(new_n778), .B2(new_n780), .ZN(G1333gat));
  NAND3_X1  g580(.A1(new_n775), .A2(G71gat), .A3(new_n696), .ZN(new_n782));
  XOR2_X1   g581(.A(new_n782), .B(KEYINPUT115), .Z(new_n783));
  INV_X1    g582(.A(new_n775), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n542), .B1(new_n784), .B2(new_n751), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(KEYINPUT50), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT50), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n783), .A2(new_n788), .A3(new_n785), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n789), .ZN(G1334gat));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n460), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g591(.A1(new_n653), .A2(new_n773), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n725), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(KEYINPUT51), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT117), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n797), .B1(new_n725), .B2(new_n793), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n795), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n794), .A2(KEYINPUT117), .A3(KEYINPUT51), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n723), .A2(new_n578), .A3(G85gat), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n578), .ZN(new_n803));
  INV_X1    g602(.A(new_n793), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n715), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n805), .A2(KEYINPUT116), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n578), .B1(new_n708), .B2(new_n714), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n808), .B1(new_n809), .B2(new_n804), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n723), .B1(new_n807), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n802), .B1(new_n812), .B2(new_n532), .ZN(G1336gat));
  NOR3_X1   g612(.A1(new_n578), .A2(G92gat), .A3(new_n461), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n799), .A2(new_n800), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n816));
  OAI21_X1  g615(.A(G92gat), .B1(new_n805), .B2(new_n461), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n795), .A2(new_n819), .A3(new_n798), .ZN(new_n820));
  OAI211_X1 g619(.A(KEYINPUT118), .B(new_n797), .C1(new_n725), .C2(new_n793), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n820), .A2(new_n814), .A3(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n680), .B1(new_n806), .B2(new_n810), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n822), .B1(new_n823), .B2(G92gat), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n818), .B1(new_n824), .B2(new_n816), .ZN(G1337gat));
  NOR3_X1   g624(.A1(new_n751), .A2(new_n578), .A3(G99gat), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n799), .A2(new_n800), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n695), .B1(new_n807), .B2(new_n811), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n827), .B1(new_n828), .B2(new_n494), .ZN(G1338gat));
  NOR3_X1   g628(.A1(new_n578), .A2(new_n282), .A3(G106gat), .ZN(new_n830));
  XOR2_X1   g629(.A(new_n830), .B(KEYINPUT119), .Z(new_n831));
  NAND3_X1  g630(.A1(new_n799), .A2(new_n800), .A3(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n833));
  OAI21_X1  g632(.A(G106gat), .B1(new_n805), .B2(new_n282), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n820), .A2(new_n821), .A3(new_n831), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n460), .B1(new_n806), .B2(new_n810), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n836), .B1(new_n837), .B2(G106gat), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n835), .B1(new_n838), .B2(new_n833), .ZN(G1339gat));
  AOI21_X1  g638(.A(new_n562), .B1(new_n556), .B2(new_n558), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n571), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(KEYINPUT54), .B1(new_n559), .B2(new_n563), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n842), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT120), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n844), .A2(KEYINPUT120), .A3(new_n845), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n842), .B(KEYINPUT55), .C1(new_n840), .C2(new_n843), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n851), .A2(new_n574), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n850), .A2(new_n636), .A3(new_n852), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n634), .A2(new_n626), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n630), .A2(new_n632), .A3(new_n629), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n608), .B1(new_n607), .B2(new_n609), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n625), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n854), .B(new_n857), .C1(new_n576), .C2(new_n577), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n673), .B1(new_n853), .B2(new_n858), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n844), .A2(KEYINPUT120), .A3(new_n845), .ZN(new_n860));
  AOI21_X1  g659(.A(KEYINPUT120), .B1(new_n844), .B2(new_n845), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n852), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n854), .A2(new_n857), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n707), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n653), .B1(new_n859), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n674), .A2(new_n578), .A3(new_n773), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n723), .A2(new_n680), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n868), .A2(new_n520), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n636), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g672(.A1(new_n871), .A2(new_n803), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g674(.A1(new_n871), .A2(new_n716), .ZN(new_n876));
  NOR2_X1   g675(.A1(KEYINPUT121), .A2(G127gat), .ZN(new_n877));
  XOR2_X1   g676(.A(new_n876), .B(new_n877), .Z(G1342gat));
  NAND2_X1  g677(.A1(new_n871), .A2(new_n673), .ZN(new_n879));
  NOR2_X1   g678(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n880));
  AND2_X1   g679(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n882), .B1(new_n879), .B2(new_n880), .ZN(G1343gat));
  INV_X1    g682(.A(KEYINPUT123), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n870), .A2(new_n741), .ZN(new_n885));
  XOR2_X1   g684(.A(KEYINPUT122), .B(KEYINPUT57), .Z(new_n886));
  AOI21_X1  g685(.A(new_n886), .B1(new_n867), .B2(new_n460), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT57), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n636), .A2(new_n852), .A3(new_n846), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n673), .B1(new_n889), .B2(new_n858), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n653), .B1(new_n864), .B2(new_n890), .ZN(new_n891));
  AOI211_X1 g690(.A(new_n888), .B(new_n282), .C1(new_n891), .C2(new_n866), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n636), .B(new_n885), .C1(new_n887), .C2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n884), .B1(new_n893), .B2(G141gat), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n867), .A2(new_n460), .A3(new_n869), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n636), .A2(new_n203), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n895), .A2(new_n696), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n897), .B1(new_n893), .B2(G141gat), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n894), .A2(new_n898), .A3(KEYINPUT58), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT58), .ZN(new_n900));
  AOI221_X4 g699(.A(new_n897), .B1(new_n884), .B2(new_n900), .C1(G141gat), .C2(new_n893), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n899), .A2(new_n901), .ZN(G1344gat));
  NOR2_X1   g701(.A1(new_n895), .A2(new_n696), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n205), .A3(new_n803), .ZN(new_n904));
  INV_X1    g703(.A(new_n885), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n867), .A2(new_n460), .ZN(new_n906));
  INV_X1    g705(.A(new_n886), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n892), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n905), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AOI211_X1 g709(.A(KEYINPUT59), .B(new_n205), .C1(new_n910), .C2(new_n803), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT59), .ZN(new_n912));
  OAI21_X1  g711(.A(KEYINPUT124), .B1(new_n707), .B2(new_n862), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT124), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n673), .A2(new_n914), .A3(new_n852), .A4(new_n850), .ZN(new_n915));
  INV_X1    g714(.A(new_n863), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n913), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(new_n890), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n716), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(new_n866), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n460), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(new_n888), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n867), .A2(new_n460), .A3(new_n886), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n924), .A2(new_n803), .A3(new_n885), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n912), .B1(new_n925), .B2(G148gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n904), .B1(new_n911), .B2(new_n926), .ZN(G1345gat));
  NAND3_X1  g726(.A1(new_n903), .A2(new_n212), .A3(new_n716), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n910), .A2(new_n716), .ZN(new_n929));
  OAI211_X1 g728(.A(KEYINPUT125), .B(new_n928), .C1(new_n929), .C2(new_n212), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT125), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n212), .B1(new_n910), .B2(new_n716), .ZN(new_n932));
  INV_X1    g731(.A(new_n928), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n930), .A2(new_n934), .ZN(G1346gat));
  AOI21_X1  g734(.A(G162gat), .B1(new_n903), .B2(new_n673), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n707), .A2(new_n213), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n936), .B1(new_n910), .B2(new_n937), .ZN(G1347gat));
  NOR2_X1   g737(.A1(new_n773), .A2(new_n399), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n676), .A2(new_n461), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n867), .A2(new_n282), .A3(new_n522), .A4(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n942), .A2(KEYINPUT126), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n942), .A2(KEYINPUT126), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n939), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(G169gat), .B1(new_n941), .B2(new_n773), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1348gat));
  NOR3_X1   g746(.A1(new_n941), .A2(new_n361), .A3(new_n578), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n803), .B1(new_n943), .B2(new_n944), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n948), .B1(new_n949), .B2(new_n361), .ZN(G1349gat));
  OR3_X1    g749(.A1(new_n941), .A2(new_n653), .A3(new_n410), .ZN(new_n951));
  INV_X1    g750(.A(G183gat), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n952), .B1(new_n941), .B2(new_n653), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n951), .B(new_n953), .C1(KEYINPUT127), .C2(KEYINPUT60), .ZN(new_n954));
  NAND2_X1  g753(.A1(KEYINPUT127), .A2(KEYINPUT60), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n954), .B(new_n955), .ZN(G1350gat));
  OAI211_X1 g755(.A(new_n396), .B(new_n673), .C1(new_n943), .C2(new_n944), .ZN(new_n957));
  AOI211_X1 g756(.A(KEYINPUT61), .B(new_n396), .C1(new_n942), .C2(new_n673), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT61), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n942), .A2(new_n673), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n959), .B1(new_n960), .B2(G190gat), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n957), .B1(new_n958), .B2(new_n961), .ZN(G1351gat));
  NAND2_X1  g761(.A1(new_n695), .A2(new_n940), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n906), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n964), .A2(new_n231), .A3(new_n636), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n963), .B1(new_n922), .B2(new_n923), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n966), .A2(new_n636), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n965), .B1(new_n967), .B2(new_n231), .ZN(G1352gat));
  NAND3_X1  g767(.A1(new_n964), .A2(new_n232), .A3(new_n803), .ZN(new_n969));
  XOR2_X1   g768(.A(new_n969), .B(KEYINPUT62), .Z(new_n970));
  AOI211_X1 g769(.A(new_n578), .B(new_n963), .C1(new_n922), .C2(new_n923), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n970), .B1(new_n971), .B2(new_n232), .ZN(G1353gat));
  AOI21_X1  g771(.A(new_n653), .B1(new_n239), .B2(new_n241), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n964), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n966), .A2(new_n716), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n975), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n976));
  AOI21_X1  g775(.A(KEYINPUT63), .B1(new_n975), .B2(G211gat), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n974), .B1(new_n976), .B2(new_n977), .ZN(G1354gat));
  AOI21_X1  g777(.A(G218gat), .B1(new_n964), .B2(new_n673), .ZN(new_n979));
  AND2_X1   g778(.A1(new_n673), .A2(G218gat), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n979), .B1(new_n966), .B2(new_n980), .ZN(G1355gat));
endmodule


