

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790;

  XNOR2_X1 U374 ( .A(n373), .B(n526), .ZN(n773) );
  XNOR2_X1 U375 ( .A(n488), .B(n487), .ZN(n766) );
  AND2_X1 U376 ( .A1(n579), .A2(n565), .ZN(n566) );
  OR2_X1 U377 ( .A1(G902), .A2(n751), .ZN(n351) );
  AND2_X1 U378 ( .A1(n459), .A2(KEYINPUT70), .ZN(n352) );
  AND2_X1 U379 ( .A1(n476), .A2(n475), .ZN(n353) );
  NOR2_X2 U380 ( .A1(n787), .A2(n571), .ZN(n417) );
  XNOR2_X2 U381 ( .A(n418), .B(KEYINPUT35), .ZN(n787) );
  XNOR2_X2 U382 ( .A(n640), .B(KEYINPUT81), .ZN(n650) );
  XNOR2_X2 U383 ( .A(G143), .B(G128), .ZN(n510) );
  XNOR2_X2 U384 ( .A(n516), .B(n484), .ZN(n768) );
  XNOR2_X2 U385 ( .A(n427), .B(n483), .ZN(n516) );
  XNOR2_X2 U386 ( .A(G116), .B(G113), .ZN(n486) );
  NOR2_X1 U387 ( .A1(n755), .A2(G902), .ZN(n374) );
  AND2_X1 U388 ( .A1(n376), .A2(n789), .ZN(n628) );
  INV_X1 U389 ( .A(n446), .ZN(n693) );
  NAND2_X1 U390 ( .A1(n700), .A2(n696), .ZN(n710) );
  INV_X2 U391 ( .A(G953), .ZN(n782) );
  XNOR2_X1 U392 ( .A(n375), .B(KEYINPUT112), .ZN(n789) );
  AND2_X1 U393 ( .A1(n583), .A2(n582), .ZN(n692) );
  XNOR2_X1 U394 ( .A(n550), .B(n351), .ZN(n581) );
  INV_X1 U395 ( .A(KEYINPUT47), .ZN(n356) );
  AND2_X1 U396 ( .A1(n624), .A2(n377), .ZN(n376) );
  NAND2_X1 U397 ( .A1(n384), .A2(n383), .ZN(n388) );
  OR2_X1 U398 ( .A1(n710), .A2(KEYINPUT79), .ZN(n406) );
  INV_X1 U399 ( .A(n619), .ZN(n384) );
  INV_X1 U400 ( .A(n715), .ZN(n632) );
  XNOR2_X1 U401 ( .A(n611), .B(KEYINPUT1), .ZN(n715) );
  XNOR2_X1 U402 ( .A(n424), .B(n396), .ZN(n608) );
  XNOR2_X1 U403 ( .A(n561), .B(n560), .ZN(n583) );
  AND2_X1 U404 ( .A1(n401), .A2(n400), .ZN(n592) );
  XNOR2_X1 U405 ( .A(n403), .B(n402), .ZN(n401) );
  NOR2_X1 U406 ( .A1(n591), .A2(n782), .ZN(n403) );
  INV_X1 U407 ( .A(n513), .ZN(n379) );
  XNOR2_X1 U408 ( .A(n500), .B(KEYINPUT14), .ZN(n502) );
  XNOR2_X1 U409 ( .A(n382), .B(G140), .ZN(n526) );
  INV_X1 U410 ( .A(KEYINPUT89), .ZN(n359) );
  INV_X1 U411 ( .A(KEYINPUT32), .ZN(n415) );
  INV_X1 U412 ( .A(G137), .ZN(n382) );
  INV_X1 U413 ( .A(G900), .ZN(n400) );
  INV_X1 U414 ( .A(KEYINPUT105), .ZN(n402) );
  BUF_X1 U415 ( .A(G113), .Z(n437) );
  INV_X1 U416 ( .A(KEYINPUT101), .ZN(n407) );
  INV_X1 U417 ( .A(G101), .ZN(n380) );
  AND2_X1 U418 ( .A1(n386), .A2(n385), .ZN(n392) );
  XNOR2_X1 U419 ( .A(n416), .B(n414), .ZN(n785) );
  NAND2_X1 U420 ( .A1(n394), .A2(n397), .ZN(n387) );
  NOR2_X1 U421 ( .A1(n446), .A2(n356), .ZN(n355) );
  NAND2_X1 U422 ( .A1(n399), .A2(n398), .ZN(n394) );
  INV_X1 U423 ( .A(n618), .ZN(n398) );
  INV_X1 U424 ( .A(n388), .ZN(n393) );
  XNOR2_X1 U425 ( .A(n505), .B(KEYINPUT0), .ZN(n579) );
  NAND2_X1 U426 ( .A1(n372), .A2(KEYINPUT39), .ZN(n371) );
  INV_X2 U427 ( .A(n692), .ZN(n696) );
  NOR2_X1 U428 ( .A1(n621), .A2(n504), .ZN(n505) );
  AND2_X1 U429 ( .A1(n367), .A2(n365), .ZN(n364) );
  NOR2_X1 U430 ( .A1(n594), .A2(n361), .ZN(n597) );
  AND2_X1 U431 ( .A1(n369), .A2(n368), .ZN(n367) );
  XNOR2_X1 U432 ( .A(n395), .B(n595), .ZN(n596) );
  AND2_X2 U433 ( .A1(n718), .A2(n719), .ZN(n716) );
  NAND2_X1 U434 ( .A1(n608), .A2(n633), .ZN(n395) );
  INV_X1 U435 ( .A(n583), .ZN(n409) );
  XNOR2_X1 U436 ( .A(n520), .B(n519), .ZN(n611) );
  AND2_X1 U437 ( .A1(n459), .A2(n370), .ZN(n361) );
  NOR2_X1 U438 ( .A1(n606), .A2(KEYINPUT70), .ZN(n366) );
  XNOR2_X1 U439 ( .A(n449), .B(n448), .ZN(n755) );
  NOR2_X1 U440 ( .A1(n735), .A2(G953), .ZN(n501) );
  XNOR2_X1 U441 ( .A(n412), .B(n410), .ZN(n663) );
  XNOR2_X1 U442 ( .A(n360), .B(n359), .ZN(n735) );
  XNOR2_X1 U443 ( .A(n461), .B(n521), .ZN(n532) );
  XNOR2_X1 U444 ( .A(n774), .B(G146), .ZN(n518) );
  XNOR2_X1 U445 ( .A(n381), .B(n379), .ZN(n515) );
  XNOR2_X1 U446 ( .A(n556), .B(n413), .ZN(n412) );
  XNOR2_X1 U447 ( .A(n547), .B(n511), .ZN(n774) );
  XNOR2_X1 U448 ( .A(n526), .B(n514), .ZN(n381) );
  XNOR2_X1 U449 ( .A(n425), .B(KEYINPUT103), .ZN(n396) );
  XNOR2_X1 U450 ( .A(n553), .B(n551), .ZN(n411) );
  XNOR2_X1 U451 ( .A(n437), .B(G122), .ZN(n553) );
  XNOR2_X1 U452 ( .A(n510), .B(G134), .ZN(n547) );
  XNOR2_X1 U453 ( .A(n486), .B(n485), .ZN(n488) );
  XNOR2_X1 U454 ( .A(n552), .B(n554), .ZN(n413) );
  XNOR2_X1 U455 ( .A(n575), .B(n415), .ZN(n414) );
  AND2_X1 U456 ( .A1(n356), .A2(n405), .ZN(n404) );
  XOR2_X1 U457 ( .A(KEYINPUT17), .B(KEYINPUT87), .Z(n490) );
  XOR2_X1 U458 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n554) );
  XNOR2_X1 U459 ( .A(KEYINPUT86), .B(G110), .ZN(n483) );
  NAND2_X1 U460 ( .A1(G234), .A2(G237), .ZN(n500) );
  INV_X1 U461 ( .A(KEYINPUT3), .ZN(n485) );
  XOR2_X1 U462 ( .A(G140), .B(G104), .Z(n552) );
  XNOR2_X1 U463 ( .A(KEYINPUT5), .B(G137), .ZN(n507) );
  XNOR2_X1 U464 ( .A(n513), .B(n510), .ZN(n422) );
  NOR2_X2 U465 ( .A1(n706), .A2(n707), .ZN(n711) );
  NAND2_X1 U466 ( .A1(n357), .A2(n354), .ZN(n623) );
  NAND2_X1 U467 ( .A1(n355), .A2(n406), .ZN(n354) );
  NAND2_X1 U468 ( .A1(n358), .A2(n404), .ZN(n357) );
  NAND2_X1 U469 ( .A1(n693), .A2(n710), .ZN(n358) );
  NAND2_X1 U470 ( .A1(n502), .A2(G952), .ZN(n360) );
  NAND2_X1 U471 ( .A1(n364), .A2(n362), .ZN(n607) );
  NAND2_X1 U472 ( .A1(n366), .A2(n363), .ZN(n362) );
  INV_X1 U473 ( .A(n459), .ZN(n363) );
  NAND2_X1 U474 ( .A1(n366), .A2(n593), .ZN(n365) );
  NAND2_X1 U475 ( .A1(n606), .A2(KEYINPUT70), .ZN(n368) );
  NAND2_X1 U476 ( .A1(n352), .A2(n370), .ZN(n369) );
  INV_X1 U477 ( .A(n593), .ZN(n370) );
  INV_X1 U478 ( .A(n372), .ZN(n443) );
  NAND2_X1 U479 ( .A1(n597), .A2(n596), .ZN(n372) );
  NAND2_X1 U480 ( .A1(n466), .A2(n465), .ZN(n641) );
  NAND2_X1 U481 ( .A1(n443), .A2(n467), .ZN(n465) );
  AND2_X2 U482 ( .A1(n371), .A2(n469), .ZN(n466) );
  XNOR2_X1 U483 ( .A(n411), .B(n373), .ZN(n410) );
  XNOR2_X2 U484 ( .A(n525), .B(n524), .ZN(n373) );
  XNOR2_X2 U485 ( .A(n374), .B(n537), .ZN(n718) );
  NAND2_X1 U486 ( .A1(n620), .A2(n715), .ZN(n375) );
  INV_X1 U487 ( .A(n690), .ZN(n377) );
  XNOR2_X2 U488 ( .A(n378), .B(n539), .ZN(n738) );
  NAND2_X1 U489 ( .A1(n453), .A2(n715), .ZN(n378) );
  XNOR2_X2 U490 ( .A(n380), .B(KEYINPUT69), .ZN(n513) );
  NAND2_X1 U491 ( .A1(n696), .A2(n457), .ZN(n383) );
  NAND2_X1 U492 ( .A1(n387), .A2(n456), .ZN(n385) );
  NAND2_X1 U493 ( .A1(n388), .A2(n456), .ZN(n386) );
  NAND2_X1 U494 ( .A1(n392), .A2(n389), .ZN(n620) );
  NAND2_X1 U495 ( .A1(n390), .A2(n393), .ZN(n389) );
  AND2_X1 U496 ( .A1(n391), .A2(n394), .ZN(n390) );
  AND2_X1 U497 ( .A1(n397), .A2(KEYINPUT36), .ZN(n391) );
  NAND2_X1 U498 ( .A1(n618), .A2(n457), .ZN(n397) );
  NOR2_X1 U499 ( .A1(n696), .A2(n457), .ZN(n399) );
  NAND2_X1 U500 ( .A1(n502), .A2(G902), .ZN(n591) );
  INV_X1 U501 ( .A(KEYINPUT79), .ZN(n405) );
  XNOR2_X2 U502 ( .A(n408), .B(n407), .ZN(n700) );
  NAND2_X1 U503 ( .A1(n581), .A2(n409), .ZN(n408) );
  NAND2_X1 U504 ( .A1(n417), .A2(n785), .ZN(n452) );
  AND2_X1 U505 ( .A1(n585), .A2(n574), .ZN(n416) );
  NAND2_X1 U506 ( .A1(n563), .A2(n626), .ZN(n418) );
  NOR2_X1 U507 ( .A1(n668), .A2(n643), .ZN(n496) );
  XNOR2_X1 U508 ( .A(n420), .B(n419), .ZN(n668) );
  XNOR2_X1 U509 ( .A(n766), .B(n494), .ZN(n419) );
  XNOR2_X1 U510 ( .A(n768), .B(n421), .ZN(n420) );
  XNOR2_X1 U511 ( .A(n493), .B(n422), .ZN(n421) );
  XNOR2_X1 U512 ( .A(n424), .B(n425), .ZN(n423) );
  NOR2_X2 U513 ( .A1(n655), .A2(G902), .ZN(n424) );
  XOR2_X1 U514 ( .A(n512), .B(G472), .Z(n425) );
  XNOR2_X1 U515 ( .A(n463), .B(n462), .ZN(n642) );
  INV_X1 U516 ( .A(KEYINPUT85), .ZN(n462) );
  XNOR2_X1 U517 ( .A(G902), .B(KEYINPUT15), .ZN(n463) );
  XNOR2_X1 U518 ( .A(n522), .B(n458), .ZN(n606) );
  XNOR2_X1 U519 ( .A(KEYINPUT96), .B(KEYINPUT21), .ZN(n458) );
  AND2_X1 U520 ( .A1(n572), .A2(n716), .ZN(n453) );
  NAND2_X1 U521 ( .A1(n642), .A2(G234), .ZN(n461) );
  XNOR2_X1 U522 ( .A(G128), .B(G119), .ZN(n527) );
  INV_X1 U523 ( .A(KEYINPUT10), .ZN(n524) );
  XNOR2_X1 U524 ( .A(n498), .B(KEYINPUT88), .ZN(n633) );
  XNOR2_X1 U525 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U526 ( .A(KEYINPUT4), .B(G131), .ZN(n511) );
  XNOR2_X1 U527 ( .A(n491), .B(KEYINPUT18), .ZN(n492) );
  OR2_X1 U528 ( .A1(G237), .A2(G902), .ZN(n497) );
  INV_X1 U529 ( .A(G902), .ZN(n557) );
  XNOR2_X1 U530 ( .A(n534), .B(n533), .ZN(n536) );
  INV_X1 U531 ( .A(KEYINPUT95), .ZN(n533) );
  XOR2_X1 U532 ( .A(KEYINPUT9), .B(G122), .Z(n545) );
  XNOR2_X1 U533 ( .A(G116), .B(G107), .ZN(n544) );
  XNOR2_X1 U534 ( .A(G143), .B(G131), .ZN(n551) );
  NOR2_X1 U535 ( .A1(G237), .A2(G953), .ZN(n506) );
  NAND2_X1 U536 ( .A1(n478), .A2(n477), .ZN(n476) );
  NOR2_X1 U537 ( .A1(n645), .A2(n654), .ZN(n477) );
  NAND2_X1 U538 ( .A1(n474), .A2(n654), .ZN(n473) );
  NAND2_X1 U539 ( .A1(n471), .A2(n480), .ZN(n470) );
  NAND2_X1 U540 ( .A1(n706), .A2(KEYINPUT39), .ZN(n469) );
  AND2_X1 U541 ( .A1(n600), .A2(n468), .ZN(n467) );
  INV_X1 U542 ( .A(KEYINPUT39), .ZN(n468) );
  INV_X1 U543 ( .A(KEYINPUT19), .ZN(n499) );
  XNOR2_X1 U544 ( .A(KEYINPUT16), .B(G122), .ZN(n484) );
  XNOR2_X1 U545 ( .A(n531), .B(KEYINPUT23), .ZN(n448) );
  XNOR2_X1 U546 ( .A(n530), .B(n773), .ZN(n449) );
  AND2_X1 U547 ( .A1(n658), .A2(G953), .ZN(n758) );
  INV_X1 U548 ( .A(KEYINPUT36), .ZN(n456) );
  INV_X1 U549 ( .A(n636), .ZN(n454) );
  INV_X1 U550 ( .A(KEYINPUT120), .ZN(n444) );
  AND2_X1 U551 ( .A1(n650), .A2(n662), .ZN(n426) );
  XOR2_X1 U552 ( .A(G104), .B(G107), .Z(n427) );
  AND2_X1 U553 ( .A1(n612), .A2(n611), .ZN(n428) );
  AND2_X1 U554 ( .A1(n447), .A2(n611), .ZN(n429) );
  AND2_X1 U555 ( .A1(n762), .A2(KEYINPUT65), .ZN(n430) );
  XNOR2_X1 U556 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n431) );
  BUF_X1 U557 ( .A(n655), .Z(n432) );
  NAND2_X1 U558 ( .A1(n490), .A2(n489), .ZN(n435) );
  NAND2_X1 U559 ( .A1(n433), .A2(n434), .ZN(n436) );
  NAND2_X1 U560 ( .A1(n435), .A2(n436), .ZN(n494) );
  INV_X1 U561 ( .A(n490), .ZN(n433) );
  INV_X1 U562 ( .A(n489), .ZN(n434) );
  NAND2_X1 U563 ( .A1(n704), .A2(n643), .ZN(n478) );
  AND2_X1 U564 ( .A1(n579), .A2(n738), .ZN(n540) );
  BUF_X1 U565 ( .A(n766), .Z(n438) );
  XNOR2_X1 U566 ( .A(n439), .B(n440), .ZN(n786) );
  NAND2_X1 U567 ( .A1(n739), .A2(n428), .ZN(n439) );
  XOR2_X1 U568 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n440) );
  XNOR2_X1 U569 ( .A(n423), .B(KEYINPUT6), .ZN(n616) );
  BUF_X1 U570 ( .A(n616), .Z(n572) );
  NOR2_X1 U571 ( .A1(n618), .A2(n696), .ZN(n441) );
  NAND2_X1 U572 ( .A1(n466), .A2(n465), .ZN(n442) );
  XNOR2_X1 U573 ( .A(n766), .B(n513), .ZN(n455) );
  XNOR2_X1 U574 ( .A(n455), .B(n509), .ZN(n464) );
  XNOR2_X1 U575 ( .A(n464), .B(n518), .ZN(n655) );
  NOR2_X1 U576 ( .A1(n703), .A2(n705), .ZN(n737) );
  AND2_X2 U577 ( .A1(n481), .A2(n762), .ZN(n703) );
  XNOR2_X1 U578 ( .A(n445), .B(n444), .ZN(n742) );
  AND2_X1 U579 ( .A1(n741), .A2(n740), .ZN(n445) );
  NAND2_X1 U580 ( .A1(n750), .A2(G210), .ZN(n672) );
  NAND2_X2 U581 ( .A1(n479), .A2(n353), .ZN(n750) );
  NAND2_X1 U582 ( .A1(n612), .A2(n429), .ZN(n446) );
  INV_X1 U583 ( .A(n621), .ZN(n447) );
  AND2_X2 U584 ( .A1(n426), .A2(n762), .ZN(n704) );
  NAND2_X1 U585 ( .A1(n450), .A2(n589), .ZN(n590) );
  XNOR2_X1 U586 ( .A(n452), .B(n451), .ZN(n450) );
  INV_X1 U587 ( .A(KEYINPUT44), .ZN(n451) );
  NAND2_X1 U588 ( .A1(n715), .A2(n716), .ZN(n578) );
  NAND2_X1 U589 ( .A1(n443), .A2(n454), .ZN(n625) );
  INV_X1 U590 ( .A(KEYINPUT111), .ZN(n457) );
  XNOR2_X1 U591 ( .A(n592), .B(n460), .ZN(n459) );
  INV_X1 U592 ( .A(KEYINPUT106), .ZN(n460) );
  NOR2_X2 U593 ( .A1(n666), .A2(n758), .ZN(n667) );
  NOR2_X2 U594 ( .A1(n659), .A2(n758), .ZN(n661) );
  NOR2_X2 U595 ( .A1(n673), .A2(n758), .ZN(n675) );
  NAND2_X1 U596 ( .A1(n472), .A2(n470), .ZN(n479) );
  NOR2_X1 U597 ( .A1(n703), .A2(n473), .ZN(n472) );
  NAND2_X1 U598 ( .A1(n641), .A2(n692), .ZN(n603) );
  INV_X1 U599 ( .A(n704), .ZN(n471) );
  NAND2_X1 U600 ( .A1(n480), .A2(n642), .ZN(n474) );
  NAND2_X1 U601 ( .A1(n481), .A2(n430), .ZN(n475) );
  XNOR2_X1 U602 ( .A(n653), .B(KEYINPUT80), .ZN(n481) );
  INV_X1 U603 ( .A(n645), .ZN(n480) );
  BUF_X1 U604 ( .A(n423), .Z(n721) );
  BUF_X1 U605 ( .A(n750), .Z(n754) );
  XNOR2_X2 U606 ( .A(G146), .B(G125), .ZN(n525) );
  XNOR2_X1 U607 ( .A(KEYINPUT22), .B(KEYINPUT67), .ZN(n482) );
  INV_X1 U608 ( .A(KEYINPUT4), .ZN(n491) );
  INV_X1 U609 ( .A(n685), .ZN(n571) );
  XNOR2_X1 U610 ( .A(n525), .B(n492), .ZN(n493) );
  XNOR2_X1 U611 ( .A(n538), .B(KEYINPUT73), .ZN(n539) );
  XNOR2_X1 U612 ( .A(KEYINPUT75), .B(KEYINPUT38), .ZN(n599) );
  XNOR2_X1 U613 ( .A(KEYINPUT71), .B(G469), .ZN(n519) );
  XNOR2_X1 U614 ( .A(n619), .B(n499), .ZN(n621) );
  INV_X1 U615 ( .A(n642), .ZN(n643) );
  XOR2_X1 U616 ( .A(KEYINPUT72), .B(G119), .Z(n487) );
  NAND2_X1 U617 ( .A1(G224), .A2(n782), .ZN(n489) );
  NAND2_X1 U618 ( .A1(G210), .A2(n497), .ZN(n495) );
  XNOR2_X1 U619 ( .A(n496), .B(n495), .ZN(n598) );
  NAND2_X1 U620 ( .A1(n497), .A2(G214), .ZN(n498) );
  NAND2_X1 U621 ( .A1(n598), .A2(n633), .ZN(n619) );
  XNOR2_X1 U622 ( .A(n501), .B(KEYINPUT90), .ZN(n593) );
  XNOR2_X1 U623 ( .A(G898), .B(KEYINPUT91), .ZN(n761) );
  NAND2_X1 U624 ( .A1(G953), .A2(n761), .ZN(n769) );
  NOR2_X1 U625 ( .A1(n769), .A2(n591), .ZN(n503) );
  NOR2_X1 U626 ( .A1(n593), .A2(n503), .ZN(n504) );
  XNOR2_X1 U627 ( .A(n506), .B(KEYINPUT76), .ZN(n555) );
  NAND2_X1 U628 ( .A1(n555), .A2(G210), .ZN(n508) );
  XNOR2_X1 U629 ( .A(n508), .B(n507), .ZN(n509) );
  INV_X1 U630 ( .A(KEYINPUT74), .ZN(n512) );
  NAND2_X1 U631 ( .A1(G227), .A2(n782), .ZN(n514) );
  XNOR2_X1 U632 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U633 ( .A(n518), .B(n517), .ZN(n744) );
  NOR2_X1 U634 ( .A1(n744), .A2(G902), .ZN(n520) );
  XOR2_X1 U635 ( .A(KEYINPUT20), .B(KEYINPUT93), .Z(n521) );
  NAND2_X1 U636 ( .A1(G221), .A2(n532), .ZN(n522) );
  INV_X1 U637 ( .A(n606), .ZN(n719) );
  NAND2_X1 U638 ( .A1(G234), .A2(n782), .ZN(n523) );
  XOR2_X1 U639 ( .A(KEYINPUT8), .B(n523), .Z(n541) );
  NAND2_X1 U640 ( .A1(n541), .A2(G221), .ZN(n531) );
  XOR2_X1 U641 ( .A(KEYINPUT24), .B(G110), .Z(n528) );
  XNOR2_X1 U642 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U643 ( .A(n529), .B(KEYINPUT92), .Z(n530) );
  NAND2_X1 U644 ( .A1(G217), .A2(n532), .ZN(n534) );
  XNOR2_X1 U645 ( .A(KEYINPUT94), .B(KEYINPUT25), .ZN(n535) );
  INV_X1 U646 ( .A(KEYINPUT33), .ZN(n538) );
  XNOR2_X1 U647 ( .A(n540), .B(KEYINPUT34), .ZN(n563) );
  XNOR2_X1 U648 ( .A(KEYINPUT100), .B(G478), .ZN(n550) );
  XOR2_X1 U649 ( .A(KEYINPUT99), .B(KEYINPUT7), .Z(n543) );
  NAND2_X1 U650 ( .A1(G217), .A2(n541), .ZN(n542) );
  XOR2_X1 U651 ( .A(n543), .B(n542), .Z(n549) );
  XNOR2_X1 U652 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U653 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U654 ( .A(n549), .B(n548), .ZN(n751) );
  AND2_X1 U655 ( .A1(n555), .A2(G214), .ZN(n556) );
  NAND2_X1 U656 ( .A1(n663), .A2(n557), .ZN(n561) );
  XOR2_X1 U657 ( .A(KEYINPUT13), .B(KEYINPUT97), .Z(n559) );
  XNOR2_X1 U658 ( .A(KEYINPUT98), .B(G475), .ZN(n558) );
  XOR2_X1 U659 ( .A(n559), .B(n558), .Z(n560) );
  NAND2_X1 U660 ( .A1(n581), .A2(n583), .ZN(n562) );
  XOR2_X1 U661 ( .A(n562), .B(KEYINPUT104), .Z(n626) );
  INV_X1 U662 ( .A(n718), .ZN(n568) );
  NOR2_X1 U663 ( .A1(n583), .A2(n581), .ZN(n708) );
  NAND2_X1 U664 ( .A1(n719), .A2(n708), .ZN(n564) );
  XOR2_X1 U665 ( .A(KEYINPUT102), .B(n564), .Z(n565) );
  XNOR2_X1 U666 ( .A(n566), .B(n482), .ZN(n573) );
  NOR2_X1 U667 ( .A1(n573), .A2(n715), .ZN(n567) );
  AND2_X1 U668 ( .A1(n568), .A2(n567), .ZN(n570) );
  INV_X1 U669 ( .A(n608), .ZN(n569) );
  NAND2_X1 U670 ( .A1(n570), .A2(n569), .ZN(n685) );
  NOR2_X1 U671 ( .A1(n573), .A2(n572), .ZN(n585) );
  NOR2_X1 U672 ( .A1(n718), .A2(n632), .ZN(n574) );
  XOR2_X1 U673 ( .A(KEYINPUT66), .B(KEYINPUT77), .Z(n575) );
  NAND2_X1 U674 ( .A1(n716), .A2(n611), .ZN(n594) );
  INV_X1 U675 ( .A(n721), .ZN(n576) );
  NOR2_X1 U676 ( .A1(n594), .A2(n576), .ZN(n577) );
  NAND2_X1 U677 ( .A1(n579), .A2(n577), .ZN(n680) );
  NOR2_X1 U678 ( .A1(n721), .A2(n578), .ZN(n726) );
  NAND2_X1 U679 ( .A1(n726), .A2(n579), .ZN(n580) );
  XOR2_X1 U680 ( .A(KEYINPUT31), .B(n580), .Z(n699) );
  NAND2_X1 U681 ( .A1(n680), .A2(n699), .ZN(n584) );
  INV_X1 U682 ( .A(n581), .ZN(n582) );
  NAND2_X1 U683 ( .A1(n584), .A2(n710), .ZN(n588) );
  NAND2_X1 U684 ( .A1(n632), .A2(n585), .ZN(n586) );
  XNOR2_X1 U685 ( .A(KEYINPUT83), .B(n586), .ZN(n587) );
  NAND2_X1 U686 ( .A1(n587), .A2(n718), .ZN(n678) );
  AND2_X1 U687 ( .A1(n588), .A2(n678), .ZN(n589) );
  XNOR2_X2 U688 ( .A(n590), .B(n431), .ZN(n762) );
  INV_X1 U689 ( .A(KEYINPUT30), .ZN(n595) );
  INV_X1 U690 ( .A(n598), .ZN(n636) );
  XNOR2_X2 U691 ( .A(n636), .B(n599), .ZN(n706) );
  INV_X1 U692 ( .A(n706), .ZN(n600) );
  INV_X1 U693 ( .A(KEYINPUT108), .ZN(n601) );
  XNOR2_X1 U694 ( .A(n601), .B(KEYINPUT40), .ZN(n602) );
  XNOR2_X2 U695 ( .A(n603), .B(n602), .ZN(n677) );
  INV_X1 U696 ( .A(n633), .ZN(n707) );
  NAND2_X1 U697 ( .A1(n711), .A2(n708), .ZN(n605) );
  XOR2_X1 U698 ( .A(KEYINPUT109), .B(KEYINPUT41), .Z(n604) );
  XNOR2_X2 U699 ( .A(n605), .B(n604), .ZN(n739) );
  NOR2_X1 U700 ( .A1(n718), .A2(n607), .ZN(n617) );
  NAND2_X1 U701 ( .A1(n617), .A2(n608), .ZN(n610) );
  INV_X1 U702 ( .A(KEYINPUT28), .ZN(n609) );
  XNOR2_X1 U703 ( .A(n610), .B(n609), .ZN(n612) );
  NOR2_X2 U704 ( .A1(n677), .A2(n786), .ZN(n615) );
  INV_X1 U705 ( .A(KEYINPUT82), .ZN(n613) );
  XOR2_X1 U706 ( .A(n613), .B(KEYINPUT46), .Z(n614) );
  XNOR2_X1 U707 ( .A(n615), .B(n614), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U709 ( .A1(n710), .A2(KEYINPUT79), .ZN(n622) );
  AND2_X1 U710 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U711 ( .A(n625), .B(KEYINPUT107), .ZN(n627) );
  AND2_X1 U712 ( .A1(n627), .A2(n626), .ZN(n690) );
  NAND2_X1 U713 ( .A1(n629), .A2(n628), .ZN(n631) );
  INV_X1 U714 ( .A(KEYINPUT48), .ZN(n630) );
  XNOR2_X1 U715 ( .A(n631), .B(n630), .ZN(n639) );
  AND2_X1 U716 ( .A1(n441), .A2(n632), .ZN(n634) );
  NAND2_X1 U717 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U718 ( .A(n635), .B(KEYINPUT43), .ZN(n637) );
  AND2_X1 U719 ( .A1(n637), .A2(n636), .ZN(n702) );
  INV_X1 U720 ( .A(n702), .ZN(n638) );
  NAND2_X1 U721 ( .A1(n639), .A2(n638), .ZN(n640) );
  INV_X1 U722 ( .A(n700), .ZN(n686) );
  NAND2_X1 U723 ( .A1(n442), .A2(n686), .ZN(n662) );
  NAND2_X1 U724 ( .A1(KEYINPUT2), .A2(n643), .ZN(n644) );
  XOR2_X1 U725 ( .A(n644), .B(KEYINPUT68), .Z(n645) );
  AND2_X1 U726 ( .A1(KEYINPUT2), .A2(KEYINPUT78), .ZN(n646) );
  AND2_X1 U727 ( .A1(n662), .A2(n646), .ZN(n647) );
  NAND2_X1 U728 ( .A1(n650), .A2(n647), .ZN(n652) );
  AND2_X1 U729 ( .A1(n662), .A2(KEYINPUT2), .ZN(n648) );
  NOR2_X1 U730 ( .A1(n648), .A2(KEYINPUT78), .ZN(n649) );
  NAND2_X1 U731 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U732 ( .A1(n652), .A2(n651), .ZN(n653) );
  INV_X1 U733 ( .A(KEYINPUT65), .ZN(n654) );
  NAND2_X1 U734 ( .A1(n750), .A2(G472), .ZN(n657) );
  XNOR2_X1 U735 ( .A(n432), .B(KEYINPUT62), .ZN(n656) );
  XNOR2_X1 U736 ( .A(n657), .B(n656), .ZN(n659) );
  INV_X1 U737 ( .A(G952), .ZN(n658) );
  INV_X1 U738 ( .A(KEYINPUT63), .ZN(n660) );
  XNOR2_X1 U739 ( .A(n661), .B(n660), .ZN(G57) );
  XNOR2_X1 U740 ( .A(n662), .B(G134), .ZN(G36) );
  NAND2_X1 U741 ( .A1(n750), .A2(G475), .ZN(n665) );
  XNOR2_X1 U742 ( .A(n663), .B(KEYINPUT59), .ZN(n664) );
  XNOR2_X1 U743 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U744 ( .A(n667), .B(KEYINPUT60), .ZN(G60) );
  XOR2_X1 U745 ( .A(KEYINPUT84), .B(KEYINPUT54), .Z(n669) );
  XNOR2_X1 U746 ( .A(n669), .B(KEYINPUT55), .ZN(n670) );
  XNOR2_X1 U747 ( .A(n668), .B(n670), .ZN(n671) );
  XNOR2_X1 U748 ( .A(n672), .B(n671), .ZN(n673) );
  XOR2_X1 U749 ( .A(KEYINPUT121), .B(KEYINPUT56), .Z(n674) );
  XNOR2_X1 U750 ( .A(n675), .B(n674), .ZN(G51) );
  XNOR2_X1 U751 ( .A(G131), .B(KEYINPUT127), .ZN(n676) );
  XNOR2_X1 U752 ( .A(n677), .B(n676), .ZN(G33) );
  XNOR2_X1 U753 ( .A(G101), .B(n678), .ZN(G3) );
  NOR2_X1 U754 ( .A1(n680), .A2(n696), .ZN(n679) );
  XOR2_X1 U755 ( .A(G104), .B(n679), .Z(G6) );
  NOR2_X1 U756 ( .A1(n680), .A2(n700), .ZN(n684) );
  XOR2_X1 U757 ( .A(KEYINPUT27), .B(KEYINPUT113), .Z(n682) );
  XNOR2_X1 U758 ( .A(G107), .B(KEYINPUT26), .ZN(n681) );
  XNOR2_X1 U759 ( .A(n682), .B(n681), .ZN(n683) );
  XNOR2_X1 U760 ( .A(n684), .B(n683), .ZN(G9) );
  XNOR2_X1 U761 ( .A(G110), .B(n685), .ZN(G12) );
  XOR2_X1 U762 ( .A(KEYINPUT114), .B(KEYINPUT29), .Z(n688) );
  NAND2_X1 U763 ( .A1(n693), .A2(n686), .ZN(n687) );
  XNOR2_X1 U764 ( .A(n688), .B(n687), .ZN(n689) );
  XNOR2_X1 U765 ( .A(G128), .B(n689), .ZN(G30) );
  XNOR2_X1 U766 ( .A(G143), .B(n690), .ZN(n691) );
  XNOR2_X1 U767 ( .A(n691), .B(KEYINPUT115), .ZN(G45) );
  NAND2_X1 U768 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U769 ( .A(n694), .B(KEYINPUT116), .ZN(n695) );
  XNOR2_X1 U770 ( .A(G146), .B(n695), .ZN(G48) );
  NOR2_X1 U771 ( .A1(n696), .A2(n699), .ZN(n698) );
  XNOR2_X1 U772 ( .A(n437), .B(KEYINPUT117), .ZN(n697) );
  XNOR2_X1 U773 ( .A(n698), .B(n697), .ZN(G15) );
  NOR2_X1 U774 ( .A1(n700), .A2(n699), .ZN(n701) );
  XOR2_X1 U775 ( .A(G116), .B(n701), .Z(G18) );
  XOR2_X1 U776 ( .A(G140), .B(n702), .Z(G42) );
  NOR2_X1 U777 ( .A1(n704), .A2(KEYINPUT2), .ZN(n705) );
  NAND2_X1 U778 ( .A1(n707), .A2(n706), .ZN(n709) );
  NAND2_X1 U779 ( .A1(n709), .A2(n708), .ZN(n713) );
  NAND2_X1 U780 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U781 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U782 ( .A1(n714), .A2(n738), .ZN(n731) );
  NOR2_X1 U783 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U784 ( .A(n717), .B(KEYINPUT50), .ZN(n724) );
  NOR2_X1 U785 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U786 ( .A(n720), .B(KEYINPUT49), .ZN(n722) );
  NAND2_X1 U787 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U788 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U789 ( .A(n725), .B(KEYINPUT118), .ZN(n727) );
  NOR2_X1 U790 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U791 ( .A(KEYINPUT51), .B(n728), .ZN(n729) );
  NAND2_X1 U792 ( .A1(n729), .A2(n739), .ZN(n730) );
  NAND2_X1 U793 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U794 ( .A(n732), .B(KEYINPUT52), .ZN(n733) );
  XNOR2_X1 U795 ( .A(n733), .B(KEYINPUT119), .ZN(n734) );
  NOR2_X1 U796 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U797 ( .A1(n737), .A2(n736), .ZN(n741) );
  NAND2_X1 U798 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U799 ( .A1(n742), .A2(G953), .ZN(n743) );
  XNOR2_X1 U800 ( .A(n743), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U801 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n746) );
  XNOR2_X1 U802 ( .A(n744), .B(KEYINPUT57), .ZN(n745) );
  XNOR2_X1 U803 ( .A(n746), .B(n745), .ZN(n748) );
  NAND2_X1 U804 ( .A1(n750), .A2(G469), .ZN(n747) );
  XOR2_X1 U805 ( .A(n748), .B(n747), .Z(n749) );
  NOR2_X1 U806 ( .A1(n758), .A2(n749), .ZN(G54) );
  NAND2_X1 U807 ( .A1(n754), .A2(G478), .ZN(n752) );
  XNOR2_X1 U808 ( .A(n752), .B(n751), .ZN(n753) );
  NOR2_X1 U809 ( .A1(n758), .A2(n753), .ZN(G63) );
  NAND2_X1 U810 ( .A1(n754), .A2(G217), .ZN(n756) );
  XNOR2_X1 U811 ( .A(n756), .B(n755), .ZN(n757) );
  NOR2_X1 U812 ( .A1(n758), .A2(n757), .ZN(G66) );
  NAND2_X1 U813 ( .A1(G953), .A2(G224), .ZN(n759) );
  XOR2_X1 U814 ( .A(KEYINPUT61), .B(n759), .Z(n760) );
  NOR2_X1 U815 ( .A1(n761), .A2(n760), .ZN(n765) );
  INV_X1 U816 ( .A(n762), .ZN(n763) );
  NOR2_X1 U817 ( .A1(G953), .A2(n763), .ZN(n764) );
  NOR2_X1 U818 ( .A1(n765), .A2(n764), .ZN(n772) );
  XNOR2_X1 U819 ( .A(n438), .B(G101), .ZN(n767) );
  XNOR2_X1 U820 ( .A(n768), .B(n767), .ZN(n770) );
  NAND2_X1 U821 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U822 ( .A(n772), .B(n771), .ZN(G69) );
  XNOR2_X1 U823 ( .A(n773), .B(KEYINPUT123), .ZN(n775) );
  XNOR2_X1 U824 ( .A(n775), .B(n774), .ZN(n779) );
  XNOR2_X1 U825 ( .A(G227), .B(n779), .ZN(n776) );
  NAND2_X1 U826 ( .A1(n776), .A2(G900), .ZN(n777) );
  NAND2_X1 U827 ( .A1(n777), .A2(G953), .ZN(n778) );
  XOR2_X1 U828 ( .A(KEYINPUT125), .B(n778), .Z(n784) );
  XOR2_X1 U829 ( .A(KEYINPUT124), .B(n779), .Z(n780) );
  XNOR2_X1 U830 ( .A(n426), .B(n780), .ZN(n781) );
  NAND2_X1 U831 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U832 ( .A1(n784), .A2(n783), .ZN(G72) );
  XNOR2_X1 U833 ( .A(G119), .B(n785), .ZN(G21) );
  XOR2_X1 U834 ( .A(n786), .B(G137), .Z(G39) );
  XOR2_X1 U835 ( .A(G122), .B(n787), .Z(n788) );
  XNOR2_X1 U836 ( .A(KEYINPUT126), .B(n788), .ZN(G24) );
  XOR2_X1 U837 ( .A(n789), .B(G125), .Z(n790) );
  XNOR2_X1 U838 ( .A(KEYINPUT37), .B(n790), .ZN(G27) );
endmodule

