//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 1 0 0 1 1 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 1 0 0 0 0 1 0 0 0 0 1 1 0 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n815,
    new_n816, new_n817, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1012, new_n1013, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1020, new_n1021, new_n1022, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1049, new_n1050;
  AND2_X1   g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(KEYINPUT41), .ZN(new_n203));
  XNOR2_X1  g002(.A(G190gat), .B(G218gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT15), .ZN(new_n206));
  INV_X1    g005(.A(G43gat), .ZN(new_n207));
  INV_X1    g006(.A(G50gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G43gat), .A2(G50gat), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n206), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT90), .B(G36gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G29gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT91), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT91), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n212), .A2(new_n215), .A3(G29gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT14), .ZN(new_n217));
  INV_X1    g016(.A(G29gat), .ZN(new_n218));
  INV_X1    g017(.A(G36gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n222), .A2(KEYINPUT89), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT89), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n224), .B1(new_n220), .B2(new_n221), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n214), .B(new_n216), .C1(new_n223), .C2(new_n225), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n214), .A2(new_n216), .ZN(new_n227));
  INV_X1    g026(.A(new_n211), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n209), .A2(new_n206), .A3(new_n210), .ZN(new_n229));
  AND3_X1   g028(.A1(new_n228), .A2(new_n222), .A3(new_n229), .ZN(new_n230));
  AOI22_X1  g029(.A1(new_n211), .A2(new_n226), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT17), .ZN(new_n232));
  NAND2_X1  g031(.A1(G99gat), .A2(G106gat), .ZN(new_n233));
  INV_X1    g032(.A(G85gat), .ZN(new_n234));
  INV_X1    g033(.A(G92gat), .ZN(new_n235));
  AOI22_X1  g034(.A1(KEYINPUT8), .A2(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT7), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n237), .B1(new_n234), .B2(new_n235), .ZN(new_n238));
  NAND3_X1  g037(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n236), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  XOR2_X1   g039(.A(G99gat), .B(G106gat), .Z(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n211), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n230), .A2(new_n216), .A3(new_n214), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT17), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT92), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT92), .ZN(new_n248));
  AOI211_X1 g047(.A(new_n248), .B(KEYINPUT17), .C1(new_n243), .C2(new_n244), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n232), .B(new_n242), .C1(new_n247), .C2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT99), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n245), .A2(new_n246), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n248), .B1(new_n231), .B2(KEYINPUT17), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n245), .A2(KEYINPUT92), .A3(new_n246), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n256), .A2(KEYINPUT99), .A3(new_n242), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n202), .A2(KEYINPUT41), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n259), .B1(new_n231), .B2(new_n242), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n205), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  AOI211_X1 g061(.A(new_n260), .B(new_n204), .C1(new_n252), .C2(new_n257), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n203), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n250), .A2(new_n251), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT99), .B1(new_n256), .B2(new_n242), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n261), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(new_n204), .ZN(new_n268));
  INV_X1    g067(.A(new_n203), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n258), .A2(new_n261), .A3(new_n205), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(G134gat), .B(G162gat), .Z(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  AND3_X1   g072(.A1(new_n264), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n273), .B1(new_n264), .B2(new_n271), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  XOR2_X1   g075(.A(G183gat), .B(G211gat), .Z(new_n277));
  XNOR2_X1  g076(.A(G127gat), .B(G155gat), .ZN(new_n278));
  XOR2_X1   g077(.A(new_n278), .B(KEYINPUT20), .Z(new_n279));
  XNOR2_X1  g078(.A(G57gat), .B(G64gat), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT94), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT9), .ZN(new_n282));
  INV_X1    g081(.A(G71gat), .ZN(new_n283));
  INV_X1    g082(.A(G78gat), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n280), .B1(new_n281), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G71gat), .B(G78gat), .ZN(new_n287));
  OAI211_X1 g086(.A(KEYINPUT94), .B(new_n282), .C1(new_n283), .C2(new_n284), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n286), .A2(KEYINPUT95), .A3(new_n287), .A4(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n285), .A2(new_n281), .ZN(new_n290));
  XOR2_X1   g089(.A(G57gat), .B(G64gat), .Z(new_n291));
  NAND4_X1  g090(.A1(new_n290), .A2(new_n291), .A3(new_n287), .A4(new_n288), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT95), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n286), .A2(new_n288), .ZN(new_n296));
  INV_X1    g095(.A(new_n287), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT96), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT21), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  AOI22_X1  g101(.A1(new_n289), .A2(new_n294), .B1(new_n297), .B2(new_n296), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT96), .B1(new_n303), .B2(KEYINPUT21), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n302), .A2(new_n304), .A3(G231gat), .A4(G233gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  AOI22_X1  g105(.A1(new_n302), .A2(new_n304), .B1(G231gat), .B2(G233gat), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n279), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n307), .ZN(new_n309));
  INV_X1    g108(.A(new_n279), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n309), .A2(new_n305), .A3(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n312), .B(KEYINPUT98), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n308), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n313), .B1(new_n308), .B2(new_n311), .ZN(new_n316));
  XNOR2_X1  g115(.A(G15gat), .B(G22gat), .ZN(new_n317));
  INV_X1    g116(.A(G1gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n317), .A2(KEYINPUT16), .A3(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n319), .B1(new_n318), .B2(new_n317), .ZN(new_n320));
  INV_X1    g119(.A(G8gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n320), .B(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n322), .B1(KEYINPUT21), .B2(new_n303), .ZN(new_n323));
  NOR3_X1   g122(.A1(new_n315), .A2(new_n316), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n323), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n311), .ZN(new_n326));
  INV_X1    g125(.A(new_n313), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n325), .B1(new_n328), .B2(new_n314), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n277), .B1(new_n324), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n323), .B1(new_n315), .B2(new_n316), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n328), .A2(new_n325), .A3(new_n314), .ZN(new_n332));
  INV_X1    g131(.A(new_n277), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  AND2_X1   g133(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n276), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT100), .ZN(new_n337));
  INV_X1    g136(.A(new_n242), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n299), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n295), .A2(new_n298), .A3(KEYINPUT100), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(new_n242), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n303), .A2(KEYINPUT100), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n339), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n299), .A2(new_n337), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n344), .A2(new_n242), .A3(new_n340), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT10), .B1(new_n345), .B2(new_n339), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n303), .A2(KEYINPUT10), .A3(new_n338), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT101), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n347), .B(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(G230gat), .A2(G233gat), .ZN(new_n351));
  MUX2_X1   g150(.A(new_n343), .B(new_n350), .S(new_n351), .Z(new_n352));
  XOR2_X1   g151(.A(G120gat), .B(G148gat), .Z(new_n353));
  XNOR2_X1  g152(.A(new_n353), .B(KEYINPUT103), .ZN(new_n354));
  XOR2_X1   g153(.A(G176gat), .B(G204gat), .Z(new_n355));
  XNOR2_X1  g154(.A(new_n354), .B(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n351), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT102), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n359), .B1(new_n346), .B2(new_n349), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT10), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n343), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n347), .B(KEYINPUT101), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n362), .A2(KEYINPUT102), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n358), .B1(new_n360), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n357), .B1(new_n343), .B2(new_n351), .ZN(new_n366));
  OAI22_X1  g165(.A1(new_n352), .A2(new_n357), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OR3_X1    g166(.A1(new_n336), .A2(KEYINPUT104), .A3(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT104), .B1(new_n336), .B2(new_n367), .ZN(new_n369));
  AND2_X1   g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT3), .ZN(new_n371));
  XNOR2_X1  g170(.A(G155gat), .B(G162gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(G155gat), .A2(G162gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT77), .ZN(new_n374));
  XNOR2_X1  g173(.A(G141gat), .B(G148gat), .ZN(new_n375));
  AND2_X1   g174(.A1(new_n373), .A2(KEYINPUT2), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n372), .B(new_n374), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n373), .A2(KEYINPUT2), .ZN(new_n379));
  INV_X1    g178(.A(G141gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n380), .A2(G148gat), .ZN(new_n381));
  INV_X1    g180(.A(G148gat), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n382), .A2(G141gat), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n379), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n372), .B1(new_n384), .B2(new_n374), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n371), .B1(new_n378), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT1), .ZN(new_n387));
  INV_X1    g186(.A(G113gat), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n388), .A2(G120gat), .ZN(new_n389));
  INV_X1    g188(.A(G120gat), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n390), .A2(G113gat), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n387), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(G134gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(G127gat), .ZN(new_n394));
  INV_X1    g193(.A(G127gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(G134gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n392), .A2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(KEYINPUT70), .B(G113gat), .ZN(new_n399));
  OAI21_X1  g198(.A(KEYINPUT69), .B1(new_n388), .B2(G120gat), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT69), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n401), .A2(new_n390), .A3(G113gat), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n399), .A2(G120gat), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n394), .A2(new_n396), .A3(new_n387), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n398), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  XOR2_X1   g204(.A(G155gat), .B(G162gat), .Z(new_n406));
  NAND2_X1  g205(.A1(new_n382), .A2(G141gat), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n380), .A2(G148gat), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n407), .A2(new_n408), .B1(KEYINPUT2), .B2(new_n373), .ZN(new_n409));
  INV_X1    g208(.A(new_n374), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n406), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n411), .A2(KEYINPUT3), .A3(new_n377), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n386), .A2(new_n405), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n377), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n400), .A2(new_n402), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n388), .A2(KEYINPUT70), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT70), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(G113gat), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(new_n418), .A3(G120gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n404), .ZN(new_n421));
  AOI22_X1  g220(.A1(new_n420), .A2(new_n421), .B1(new_n392), .B2(new_n397), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n414), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT4), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT78), .B(KEYINPUT4), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n414), .A2(new_n422), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(G225gat), .A2(G233gat), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n430), .A2(KEYINPUT5), .ZN(new_n431));
  AND4_X1   g230(.A1(new_n413), .A2(new_n425), .A3(new_n428), .A4(new_n431), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n412), .A2(new_n405), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n430), .B1(new_n433), .B2(new_n386), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n426), .B1(new_n414), .B2(new_n422), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT79), .ZN(new_n436));
  OAI22_X1  g235(.A1(new_n435), .A2(new_n436), .B1(new_n423), .B2(KEYINPUT4), .ZN(new_n437));
  AOI211_X1 g236(.A(KEYINPUT79), .B(new_n426), .C1(new_n414), .C2(new_n422), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n434), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT5), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n414), .B(new_n422), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n440), .B1(new_n441), .B2(new_n430), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n432), .B1(new_n439), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(G1gat), .B(G29gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n445), .B(KEYINPUT0), .ZN(new_n446));
  XNOR2_X1  g245(.A(G57gat), .B(G85gat), .ZN(new_n447));
  XOR2_X1   g246(.A(new_n446), .B(new_n447), .Z(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n444), .A2(KEYINPUT6), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT85), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n444), .A2(new_n452), .A3(new_n449), .ZN(new_n453));
  OAI21_X1  g252(.A(KEYINPUT85), .B1(new_n443), .B2(new_n448), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n442), .ZN(new_n456));
  INV_X1    g255(.A(new_n432), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n448), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT80), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n443), .A2(KEYINPUT80), .A3(new_n448), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT6), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n451), .B1(new_n455), .B2(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(G8gat), .B(G36gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(G64gat), .B(G92gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n464), .B(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  AND2_X1   g266(.A1(G211gat), .A2(G218gat), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n468), .A2(KEYINPUT22), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(G204gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(G197gat), .ZN(new_n472));
  INV_X1    g271(.A(G197gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(G204gat), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT72), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n472), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n475), .B1(new_n472), .B2(new_n474), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n470), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g277(.A1(G211gat), .A2(G218gat), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n468), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n473), .A2(G204gat), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n471), .A2(G197gat), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT72), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n472), .A2(new_n474), .A3(new_n475), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n480), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n486), .A2(new_n487), .A3(new_n470), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n481), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT23), .ZN(new_n490));
  NOR3_X1   g289(.A1(new_n490), .A2(G169gat), .A3(G176gat), .ZN(new_n491));
  AOI22_X1  g290(.A1(new_n491), .A2(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n492));
  INV_X1    g291(.A(G169gat), .ZN(new_n493));
  INV_X1    g292(.A(G176gat), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(new_n494), .A3(KEYINPUT23), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT23), .B1(new_n493), .B2(new_n494), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT65), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AND3_X1   g297(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(G183gat), .A2(G190gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n492), .A2(new_n498), .A3(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT25), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n490), .B1(G169gat), .B2(G176gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(G169gat), .A2(G176gat), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n495), .A2(new_n508), .A3(KEYINPUT25), .A4(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n499), .B1(new_n502), .B2(new_n501), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n507), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT28), .ZN(new_n515));
  INV_X1    g314(.A(G190gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n516), .B1(new_n517), .B2(KEYINPUT27), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT27), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n519), .B1(KEYINPUT66), .B2(G183gat), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n515), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(KEYINPUT27), .B(G183gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n522), .A2(KEYINPUT28), .A3(new_n516), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(new_n509), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT67), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n525), .A2(KEYINPUT67), .A3(new_n509), .ZN(new_n529));
  NOR2_X1   g328(.A1(G169gat), .A2(G176gat), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT26), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT68), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n530), .A2(KEYINPUT68), .A3(new_n531), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n528), .A2(new_n529), .A3(new_n534), .A4(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n524), .A2(new_n536), .A3(new_n502), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n514), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(G226gat), .A2(G233gat), .ZN(new_n539));
  XOR2_X1   g338(.A(new_n539), .B(KEYINPUT73), .Z(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  AND3_X1   g340(.A1(new_n524), .A2(new_n536), .A3(new_n502), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n512), .B1(new_n505), .B2(new_n506), .ZN(new_n543));
  OAI21_X1  g342(.A(KEYINPUT74), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT74), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n509), .B1(new_n495), .B2(new_n497), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n511), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT25), .B1(new_n547), .B2(new_n498), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n545), .B(new_n537), .C1(new_n548), .C2(new_n512), .ZN(new_n549));
  AOI21_X1  g348(.A(KEYINPUT29), .B1(new_n544), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n539), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n489), .B(new_n541), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n489), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n539), .B1(new_n544), .B2(new_n549), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT29), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n540), .B1(new_n538), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n553), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n467), .B1(new_n552), .B2(new_n557), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n552), .A2(new_n557), .A3(new_n467), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n558), .B1(new_n559), .B2(KEYINPUT30), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n552), .A2(new_n557), .A3(new_n467), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT30), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n561), .A2(KEYINPUT76), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT76), .B1(new_n561), .B2(new_n562), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n560), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n487), .B1(new_n486), .B2(new_n470), .ZN(new_n566));
  AOI211_X1 g365(.A(new_n480), .B(new_n469), .C1(new_n484), .C2(new_n485), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n555), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n414), .B1(new_n568), .B2(new_n371), .ZN(new_n569));
  INV_X1    g368(.A(G228gat), .ZN(new_n570));
  INV_X1    g369(.A(G233gat), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT29), .B1(new_n414), .B2(new_n371), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n574), .A2(new_n489), .ZN(new_n575));
  NOR3_X1   g374(.A1(new_n569), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n414), .ZN(new_n577));
  AOI21_X1  g376(.A(KEYINPUT29), .B1(new_n481), .B2(new_n488), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n577), .B1(new_n578), .B2(KEYINPUT3), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n386), .A2(new_n555), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(new_n553), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n572), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(G22gat), .B1(new_n576), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n573), .B1(new_n569), .B2(new_n575), .ZN(new_n584));
  INV_X1    g383(.A(G22gat), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n579), .A2(new_n581), .A3(new_n572), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G78gat), .B(G106gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(KEYINPUT31), .B(G50gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n591), .A2(KEYINPUT81), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n583), .A2(new_n587), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n592), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n584), .A2(new_n585), .A3(new_n586), .A4(new_n594), .ZN(new_n595));
  OAI211_X1 g394(.A(G22gat), .B(new_n591), .C1(new_n576), .C2(new_n582), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n593), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT35), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n422), .B1(new_n542), .B2(new_n543), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n514), .A2(new_n405), .A3(new_n537), .ZN(new_n600));
  NAND2_X1  g399(.A1(G227gat), .A2(G233gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT64), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT33), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(KEYINPUT32), .ZN(new_n606));
  XOR2_X1   g405(.A(G15gat), .B(G43gat), .Z(new_n607));
  XNOR2_X1  g406(.A(G71gat), .B(G99gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n605), .A2(new_n606), .A3(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n609), .ZN(new_n611));
  OAI211_X1 g410(.A(new_n603), .B(KEYINPUT32), .C1(new_n604), .C2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n599), .A2(new_n600), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT71), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n602), .A2(KEYINPUT34), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n615), .B1(new_n614), .B2(new_n616), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT34), .ZN(new_n619));
  AOI22_X1  g418(.A1(new_n599), .A2(new_n600), .B1(G227gat), .B2(G233gat), .ZN(new_n620));
  OAI22_X1  g419(.A1(new_n617), .A2(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n613), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n614), .A2(new_n616), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT71), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n620), .A2(new_n619), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n626), .A2(new_n627), .A3(new_n610), .A4(new_n612), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n597), .A2(new_n598), .A3(new_n622), .A4(new_n628), .ZN(new_n629));
  NOR3_X1   g428(.A1(new_n463), .A2(new_n565), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT6), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n444), .A2(new_n449), .ZN(new_n632));
  AND4_X1   g431(.A1(KEYINPUT80), .A2(new_n456), .A3(new_n448), .A4(new_n457), .ZN(new_n633));
  AOI21_X1  g432(.A(KEYINPUT80), .B1(new_n443), .B2(new_n448), .ZN(new_n634));
  OAI211_X1 g433(.A(new_n631), .B(new_n632), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT76), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n636), .B1(new_n559), .B2(KEYINPUT30), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n561), .A2(KEYINPUT76), .A3(new_n562), .ZN(new_n638));
  AOI22_X1  g437(.A1(new_n635), .A2(new_n450), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AND4_X1   g438(.A1(KEYINPUT30), .A2(new_n552), .A3(new_n557), .A4(new_n467), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT75), .ZN(new_n641));
  NOR3_X1   g440(.A1(new_n640), .A2(new_n641), .A3(new_n558), .ZN(new_n642));
  INV_X1    g441(.A(new_n558), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n552), .A2(new_n557), .A3(KEYINPUT30), .A4(new_n467), .ZN(new_n644));
  AOI21_X1  g443(.A(KEYINPUT75), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT86), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n622), .A2(new_n628), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n647), .B1(new_n648), .B2(new_n597), .ZN(new_n649));
  AND4_X1   g448(.A1(new_n647), .A2(new_n597), .A3(new_n622), .A4(new_n628), .ZN(new_n650));
  OAI211_X1 g449(.A(new_n639), .B(new_n646), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n630), .B1(new_n651), .B2(KEYINPUT35), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT39), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n413), .A2(new_n425), .A3(new_n428), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT83), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n654), .A2(new_n655), .A3(new_n430), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n655), .B1(new_n654), .B2(new_n430), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n653), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n654), .A2(new_n430), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(KEYINPUT83), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n441), .A2(new_n430), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n662), .A2(new_n653), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n661), .A2(new_n656), .A3(new_n663), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n659), .A2(new_n664), .A3(KEYINPUT40), .A4(new_n448), .ZN(new_n665));
  AND3_X1   g464(.A1(new_n665), .A2(new_n454), .A3(new_n453), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n659), .A2(new_n664), .A3(new_n448), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT40), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT84), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n667), .A2(KEYINPUT84), .A3(new_n668), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n565), .A2(new_n666), .A3(new_n671), .A4(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n460), .A2(new_n461), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n674), .A2(new_n631), .A3(new_n454), .A4(new_n453), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT37), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n552), .A2(new_n676), .A3(new_n557), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n677), .A2(new_n466), .ZN(new_n678));
  INV_X1    g477(.A(new_n549), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n545), .B1(new_n514), .B2(new_n537), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n551), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n538), .A2(new_n555), .ZN(new_n682));
  INV_X1    g481(.A(new_n540), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n676), .B1(new_n685), .B2(new_n489), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n553), .B(new_n541), .C1(new_n550), .C2(new_n551), .ZN(new_n687));
  AOI21_X1  g486(.A(KEYINPUT38), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n559), .B1(new_n678), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n677), .A2(new_n466), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n676), .B1(new_n552), .B2(new_n557), .ZN(new_n691));
  OAI21_X1  g490(.A(KEYINPUT38), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n675), .A2(new_n689), .A3(new_n450), .A4(new_n692), .ZN(new_n693));
  AND3_X1   g492(.A1(new_n673), .A2(new_n693), .A3(new_n597), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n622), .A2(new_n628), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT36), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n451), .B1(new_n462), .B2(new_n632), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n641), .B1(new_n640), .B2(new_n558), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n643), .A2(KEYINPUT75), .A3(new_n644), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n563), .A2(new_n564), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n698), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n697), .B1(new_n703), .B2(new_n597), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n694), .B1(new_n704), .B2(KEYINPUT82), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT82), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n697), .B(new_n706), .C1(new_n703), .C2(new_n597), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n652), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n322), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n709), .B(new_n232), .C1(new_n247), .C2(new_n249), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT93), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n711), .B1(new_n245), .B2(new_n322), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n245), .A2(new_n711), .A3(new_n322), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(G229gat), .A2(G233gat), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n710), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT18), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n710), .A2(new_n715), .A3(KEYINPUT18), .A4(new_n716), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n716), .B(KEYINPUT13), .Z(new_n721));
  INV_X1    g520(.A(new_n714), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n722), .A2(new_n712), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n245), .A2(new_n322), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n721), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n719), .A2(new_n720), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(G113gat), .B(G141gat), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT11), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(new_n493), .ZN(new_n729));
  XNOR2_X1  g528(.A(KEYINPUT87), .B(G197gat), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(new_n731));
  XOR2_X1   g530(.A(KEYINPUT88), .B(KEYINPUT12), .Z(new_n732));
  XOR2_X1   g531(.A(new_n731), .B(new_n732), .Z(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n726), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n719), .A2(new_n733), .A3(new_n720), .A4(new_n725), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n708), .A2(new_n738), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n370), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n698), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT106), .ZN(new_n742));
  XOR2_X1   g541(.A(KEYINPUT105), .B(G1gat), .Z(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n742), .B(new_n744), .ZN(G1324gat));
  INV_X1    g544(.A(new_n740), .ZN(new_n746));
  INV_X1    g545(.A(new_n565), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(KEYINPUT42), .B1(new_n748), .B2(new_n321), .ZN(new_n749));
  XOR2_X1   g548(.A(KEYINPUT16), .B(G8gat), .Z(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  MUX2_X1   g550(.A(KEYINPUT42), .B(new_n749), .S(new_n751), .Z(G1325gat));
  OAI21_X1  g551(.A(G15gat), .B1(new_n746), .B2(new_n697), .ZN(new_n753));
  OR2_X1    g552(.A1(new_n695), .A2(G15gat), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n753), .B1(new_n746), .B2(new_n754), .ZN(G1326gat));
  INV_X1    g554(.A(new_n597), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g556(.A(KEYINPUT43), .B(G22gat), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(G1327gat));
  NAND2_X1  g558(.A1(new_n330), .A2(new_n334), .ZN(new_n760));
  INV_X1    g559(.A(new_n367), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR4_X1   g561(.A1(new_n708), .A2(new_n738), .A3(new_n276), .A4(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n763), .A2(new_n218), .A3(new_n698), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT45), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT111), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n673), .A2(new_n693), .A3(new_n597), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n639), .A2(new_n646), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n756), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n767), .A2(new_n769), .A3(new_n697), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT109), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n770), .B1(new_n652), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(KEYINPUT86), .B1(new_n756), .B2(new_n695), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n648), .A2(new_n647), .A3(new_n597), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n598), .B1(new_n703), .B2(new_n775), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n776), .A2(KEYINPUT109), .A3(new_n630), .ZN(new_n777));
  OAI21_X1  g576(.A(KEYINPUT110), .B1(new_n772), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n652), .A2(new_n771), .ZN(new_n779));
  OAI21_X1  g578(.A(KEYINPUT109), .B1(new_n776), .B2(new_n630), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT110), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n779), .A2(new_n780), .A3(new_n781), .A4(new_n770), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n778), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n276), .A2(KEYINPUT44), .ZN(new_n784));
  OAI211_X1 g583(.A(KEYINPUT108), .B(KEYINPUT44), .C1(new_n708), .C2(new_n276), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT108), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n597), .B1(new_n639), .B2(new_n646), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT82), .B1(new_n787), .B2(new_n696), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n707), .A2(new_n788), .A3(new_n767), .ZN(new_n789));
  INV_X1    g588(.A(new_n652), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n276), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT44), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n786), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AOI22_X1  g592(.A1(new_n783), .A2(new_n784), .B1(new_n785), .B2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT107), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n720), .A2(new_n725), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n733), .B1(new_n796), .B2(new_n719), .ZN(new_n797));
  INV_X1    g596(.A(new_n736), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n795), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n735), .A2(KEYINPUT107), .A3(new_n736), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n762), .A2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n766), .B1(new_n794), .B2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n785), .A2(new_n793), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n778), .A2(new_n782), .A3(new_n784), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n809), .A2(KEYINPUT111), .A3(new_n803), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n698), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n806), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n765), .B1(new_n813), .B2(new_n218), .ZN(G1328gat));
  INV_X1    g613(.A(new_n212), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n763), .A2(new_n815), .A3(new_n565), .ZN(new_n816));
  XOR2_X1   g615(.A(new_n816), .B(KEYINPUT46), .Z(new_n817));
  NOR3_X1   g616(.A1(new_n806), .A2(new_n811), .A3(new_n747), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n817), .B1(new_n818), .B2(new_n815), .ZN(G1329gat));
  INV_X1    g618(.A(KEYINPUT112), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n804), .B1(new_n807), .B2(new_n808), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n207), .B1(new_n821), .B2(new_n696), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n695), .A2(G43gat), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n763), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT47), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n820), .B1(new_n822), .B2(new_n826), .ZN(new_n827));
  OR3_X1    g626(.A1(new_n822), .A2(new_n826), .A3(new_n820), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n805), .A2(new_n696), .A3(new_n810), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n824), .B1(new_n829), .B2(G43gat), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n827), .B(new_n828), .C1(new_n830), .C2(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g630(.A1(new_n805), .A2(new_n756), .A3(new_n810), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n756), .A2(new_n208), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT113), .ZN(new_n834));
  AOI22_X1  g633(.A1(new_n832), .A2(G50gat), .B1(new_n763), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n208), .B1(new_n821), .B2(new_n756), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n763), .A2(new_n834), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT48), .ZN(new_n838));
  OAI22_X1  g637(.A1(new_n835), .A2(KEYINPUT48), .B1(new_n836), .B2(new_n838), .ZN(G1331gat));
  NOR3_X1   g638(.A1(new_n336), .A2(new_n761), .A3(new_n801), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n783), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n698), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g642(.A(new_n747), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n846));
  XOR2_X1   g645(.A(new_n845), .B(new_n846), .Z(G1333gat));
  NAND3_X1  g646(.A1(new_n841), .A2(G71gat), .A3(new_n696), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n841), .A2(new_n648), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n848), .B1(new_n849), .B2(G71gat), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g650(.A1(new_n841), .A2(new_n756), .ZN(new_n852));
  XOR2_X1   g651(.A(KEYINPUT114), .B(G78gat), .Z(new_n853));
  XNOR2_X1  g652(.A(new_n852), .B(new_n853), .ZN(G1335gat));
  NAND3_X1  g653(.A1(new_n779), .A2(new_n780), .A3(new_n770), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n802), .A2(new_n760), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(new_n276), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n855), .A2(KEYINPUT51), .A3(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(KEYINPUT51), .B1(new_n855), .B2(new_n857), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n367), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(G85gat), .B1(new_n862), .B2(new_n698), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n794), .A2(new_n761), .A3(new_n856), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n812), .A2(new_n234), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(G1336gat));
  AOI21_X1  g665(.A(G92gat), .B1(new_n862), .B2(new_n565), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n809), .A2(new_n760), .A3(new_n367), .A4(new_n802), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n565), .A2(G92gat), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n868), .B(KEYINPUT52), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT52), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n869), .A2(new_n870), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n872), .B1(new_n873), .B2(new_n867), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n871), .A2(new_n874), .ZN(G1337gat));
  AOI21_X1  g674(.A(G99gat), .B1(new_n862), .B2(new_n648), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n696), .A2(G99gat), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n876), .B1(new_n864), .B2(new_n877), .ZN(G1338gat));
  INV_X1    g677(.A(G106gat), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n879), .B1(new_n864), .B2(new_n756), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n597), .A2(G106gat), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n367), .B(new_n881), .C1(new_n859), .C2(new_n860), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(KEYINPUT115), .ZN(new_n883));
  OAI21_X1  g682(.A(KEYINPUT53), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(G106gat), .B1(new_n869), .B2(new_n597), .ZN(new_n885));
  XNOR2_X1  g684(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n885), .A2(new_n882), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n884), .A2(new_n887), .ZN(G1339gat));
  NOR3_X1   g687(.A1(new_n262), .A2(new_n263), .A3(new_n203), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n269), .B1(new_n268), .B2(new_n270), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n272), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n264), .A2(new_n271), .A3(new_n273), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n723), .A2(new_n724), .A3(new_n721), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n716), .B1(new_n710), .B2(new_n715), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n731), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n736), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n367), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n365), .A2(new_n366), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT54), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n900), .B(new_n351), .C1(new_n346), .C2(new_n349), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n356), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n346), .A2(new_n349), .A3(new_n359), .ZN(new_n903));
  AOI21_X1  g702(.A(KEYINPUT102), .B1(new_n362), .B2(new_n363), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n351), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n900), .B1(new_n350), .B2(new_n358), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n902), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n899), .B1(new_n907), .B2(KEYINPUT55), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n350), .A2(new_n358), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT54), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n356), .B(new_n901), .C1(new_n910), .C2(new_n365), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT55), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n908), .A2(new_n799), .A3(new_n800), .A4(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n893), .B1(new_n898), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n736), .A2(new_n896), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n916), .B1(new_n911), .B2(new_n912), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n908), .B(new_n917), .C1(new_n274), .C2(new_n275), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n760), .B1(new_n915), .B2(new_n919), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n802), .A2(new_n335), .A3(new_n276), .A4(new_n761), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n812), .A2(new_n565), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n756), .A2(new_n695), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT117), .ZN(new_n927));
  OAI21_X1  g726(.A(G113gat), .B1(new_n927), .B2(new_n738), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n924), .A2(new_n775), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n930), .A2(new_n399), .A3(new_n801), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n928), .A2(new_n931), .ZN(G1340gat));
  NOR3_X1   g731(.A1(new_n927), .A2(new_n390), .A3(new_n761), .ZN(new_n933));
  AOI21_X1  g732(.A(G120gat), .B1(new_n930), .B2(new_n367), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n933), .A2(new_n934), .ZN(G1341gat));
  OAI21_X1  g734(.A(G127gat), .B1(new_n927), .B2(new_n760), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n930), .A2(new_n395), .A3(new_n335), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1342gat));
  OAI21_X1  g737(.A(G134gat), .B1(new_n927), .B2(new_n276), .ZN(new_n939));
  NOR4_X1   g738(.A1(new_n893), .A2(new_n801), .A3(new_n760), .A4(new_n367), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n914), .A2(new_n898), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(new_n276), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(new_n918), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n940), .B1(new_n943), .B2(new_n760), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n944), .A2(new_n812), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n893), .A2(new_n747), .ZN(new_n946));
  AOI211_X1 g745(.A(G134gat), .B(new_n946), .C1(new_n773), .C2(new_n774), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  XOR2_X1   g747(.A(new_n948), .B(KEYINPUT56), .Z(new_n949));
  NAND2_X1  g748(.A1(new_n939), .A2(new_n949), .ZN(G1343gat));
  AOI21_X1  g749(.A(new_n597), .B1(new_n920), .B2(new_n921), .ZN(new_n951));
  XOR2_X1   g750(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  OAI21_X1  g752(.A(KEYINPUT119), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT119), .ZN(new_n955));
  OAI211_X1 g754(.A(new_n955), .B(new_n952), .C1(new_n944), .C2(new_n597), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT121), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n913), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(KEYINPUT121), .B1(new_n911), .B2(new_n912), .ZN(new_n959));
  OAI211_X1 g758(.A(new_n737), .B(new_n908), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n898), .B(KEYINPUT120), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n893), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n760), .B1(new_n962), .B2(new_n919), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(new_n921), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n756), .A2(KEYINPUT57), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n954), .A2(new_n956), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n923), .A2(new_n697), .ZN(new_n968));
  INV_X1    g767(.A(new_n968), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n967), .A2(new_n737), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(KEYINPUT122), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT122), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n967), .A2(new_n972), .A3(new_n737), .A4(new_n969), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n971), .A2(G141gat), .A3(new_n973), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n696), .A2(new_n597), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n924), .A2(new_n975), .ZN(new_n976));
  AND3_X1   g775(.A1(new_n976), .A2(new_n380), .A3(new_n737), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n977), .A2(KEYINPUT58), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n974), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n953), .B1(new_n922), .B2(new_n756), .ZN(new_n980));
  AOI22_X1  g779(.A1(new_n980), .A2(new_n955), .B1(new_n964), .B2(new_n965), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n968), .B1(new_n981), .B2(new_n954), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n380), .B1(new_n982), .B2(new_n801), .ZN(new_n983));
  OAI21_X1  g782(.A(KEYINPUT58), .B1(new_n983), .B2(new_n977), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n979), .A2(new_n984), .ZN(G1344gat));
  AOI211_X1 g784(.A(KEYINPUT59), .B(new_n382), .C1(new_n982), .C2(new_n367), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT59), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n368), .A2(new_n738), .A3(new_n369), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n988), .A2(new_n963), .ZN(new_n989));
  AOI21_X1  g788(.A(KEYINPUT57), .B1(new_n989), .B2(new_n756), .ZN(new_n990));
  NOR3_X1   g789(.A1(new_n944), .A2(new_n597), .A3(new_n952), .ZN(new_n991));
  OAI211_X1 g790(.A(new_n367), .B(new_n969), .C1(new_n990), .C2(new_n991), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n987), .B1(new_n992), .B2(G148gat), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n945), .A2(new_n975), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n747), .A2(new_n382), .A3(new_n367), .ZN(new_n995));
  OAI22_X1  g794(.A1(new_n986), .A2(new_n993), .B1(new_n994), .B2(new_n995), .ZN(G1345gat));
  INV_X1    g795(.A(new_n982), .ZN(new_n997));
  OAI21_X1  g796(.A(G155gat), .B1(new_n997), .B2(new_n760), .ZN(new_n998));
  INV_X1    g797(.A(G155gat), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n976), .A2(new_n999), .A3(new_n335), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n998), .A2(new_n1000), .ZN(G1346gat));
  OAI21_X1  g800(.A(G162gat), .B1(new_n997), .B2(new_n276), .ZN(new_n1002));
  OR2_X1    g801(.A1(new_n946), .A2(G162gat), .ZN(new_n1003));
  OAI21_X1  g802(.A(new_n1002), .B1(new_n994), .B2(new_n1003), .ZN(G1347gat));
  AOI211_X1 g803(.A(new_n698), .B(new_n747), .C1(new_n920), .C2(new_n921), .ZN(new_n1005));
  AND2_X1   g804(.A1(new_n1005), .A2(new_n775), .ZN(new_n1006));
  NAND3_X1  g805(.A1(new_n1006), .A2(new_n493), .A3(new_n801), .ZN(new_n1007));
  XNOR2_X1  g806(.A(new_n1007), .B(KEYINPUT123), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1005), .A2(new_n925), .ZN(new_n1009));
  OAI21_X1  g808(.A(G169gat), .B1(new_n1009), .B2(new_n738), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1008), .A2(new_n1010), .ZN(G1348gat));
  NAND3_X1  g810(.A1(new_n1006), .A2(new_n494), .A3(new_n367), .ZN(new_n1012));
  OAI21_X1  g811(.A(G176gat), .B1(new_n1009), .B2(new_n761), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n1012), .A2(new_n1013), .ZN(G1349gat));
  NAND3_X1  g813(.A1(new_n1006), .A2(new_n522), .A3(new_n335), .ZN(new_n1015));
  OAI21_X1  g814(.A(G183gat), .B1(new_n1009), .B2(new_n760), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g816(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n1018));
  XNOR2_X1  g817(.A(new_n1017), .B(new_n1018), .ZN(G1350gat));
  OAI21_X1  g818(.A(G190gat), .B1(new_n1009), .B2(new_n276), .ZN(new_n1020));
  XNOR2_X1  g819(.A(new_n1020), .B(KEYINPUT61), .ZN(new_n1021));
  NAND3_X1  g820(.A1(new_n1006), .A2(new_n516), .A3(new_n893), .ZN(new_n1022));
  NAND2_X1  g821(.A1(new_n1021), .A2(new_n1022), .ZN(G1351gat));
  NAND2_X1  g822(.A1(new_n1005), .A2(new_n975), .ZN(new_n1024));
  NOR3_X1   g823(.A1(new_n1024), .A2(G197gat), .A3(new_n802), .ZN(new_n1025));
  XNOR2_X1  g824(.A(new_n1025), .B(KEYINPUT125), .ZN(new_n1026));
  NOR3_X1   g825(.A1(new_n696), .A2(new_n747), .A3(new_n698), .ZN(new_n1027));
  OAI21_X1  g826(.A(new_n1027), .B1(new_n990), .B2(new_n991), .ZN(new_n1028));
  OAI21_X1  g827(.A(G197gat), .B1(new_n1028), .B2(new_n738), .ZN(new_n1029));
  NAND2_X1  g828(.A1(new_n1026), .A2(new_n1029), .ZN(G1352gat));
  OAI211_X1 g829(.A(new_n367), .B(new_n1027), .C1(new_n990), .C2(new_n991), .ZN(new_n1031));
  NAND2_X1  g830(.A1(new_n1031), .A2(G204gat), .ZN(new_n1032));
  NOR2_X1   g831(.A1(new_n761), .A2(G204gat), .ZN(new_n1033));
  NAND3_X1  g832(.A1(new_n1005), .A2(new_n975), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g833(.A1(new_n1034), .A2(KEYINPUT126), .ZN(new_n1035));
  INV_X1    g834(.A(KEYINPUT126), .ZN(new_n1036));
  NAND4_X1  g835(.A1(new_n1005), .A2(new_n1036), .A3(new_n975), .A4(new_n1033), .ZN(new_n1037));
  NAND2_X1  g836(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g837(.A(KEYINPUT127), .ZN(new_n1039));
  AOI21_X1  g838(.A(new_n1039), .B1(new_n1038), .B2(KEYINPUT62), .ZN(new_n1040));
  INV_X1    g839(.A(KEYINPUT62), .ZN(new_n1041));
  AOI211_X1 g840(.A(KEYINPUT127), .B(new_n1041), .C1(new_n1035), .C2(new_n1037), .ZN(new_n1042));
  OAI221_X1 g841(.A(new_n1032), .B1(KEYINPUT62), .B2(new_n1038), .C1(new_n1040), .C2(new_n1042), .ZN(G1353gat));
  OR3_X1    g842(.A1(new_n1024), .A2(G211gat), .A3(new_n760), .ZN(new_n1044));
  OAI211_X1 g843(.A(new_n335), .B(new_n1027), .C1(new_n990), .C2(new_n991), .ZN(new_n1045));
  AND3_X1   g844(.A1(new_n1045), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1046));
  AOI21_X1  g845(.A(KEYINPUT63), .B1(new_n1045), .B2(G211gat), .ZN(new_n1047));
  OAI21_X1  g846(.A(new_n1044), .B1(new_n1046), .B2(new_n1047), .ZN(G1354gat));
  OAI21_X1  g847(.A(G218gat), .B1(new_n1028), .B2(new_n276), .ZN(new_n1049));
  OR2_X1    g848(.A1(new_n276), .A2(G218gat), .ZN(new_n1050));
  OAI21_X1  g849(.A(new_n1049), .B1(new_n1024), .B2(new_n1050), .ZN(G1355gat));
endmodule


