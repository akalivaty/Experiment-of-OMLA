//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 1 0 1 0 0 1 0 0 1 0 1 1 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n762, new_n763, new_n764,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  INV_X1    g002(.A(G140), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G125), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G140), .ZN(new_n192));
  AND3_X1   g006(.A1(new_n190), .A2(new_n192), .A3(KEYINPUT19), .ZN(new_n193));
  AOI21_X1  g007(.A(KEYINPUT19), .B1(new_n190), .B2(new_n192), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n188), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n190), .A2(new_n192), .A3(KEYINPUT16), .ZN(new_n196));
  OR3_X1    g010(.A1(new_n191), .A2(KEYINPUT16), .A3(G140), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n197), .A3(G146), .ZN(new_n198));
  INV_X1    g012(.A(G237), .ZN(new_n199));
  INV_X1    g013(.A(G953), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(G214), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G131), .ZN(new_n204));
  NOR2_X1   g018(.A1(G237), .A2(G953), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(G143), .A3(G214), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n203), .A2(new_n204), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n204), .B1(new_n203), .B2(new_n206), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n195), .B(new_n198), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  XNOR2_X1  g024(.A(G125), .B(G140), .ZN(new_n211));
  XNOR2_X1  g025(.A(new_n211), .B(new_n188), .ZN(new_n212));
  INV_X1    g026(.A(new_n206), .ZN(new_n213));
  AOI21_X1  g027(.A(G143), .B1(new_n205), .B2(G214), .ZN(new_n214));
  OAI211_X1 g028(.A(KEYINPUT18), .B(G131), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(KEYINPUT18), .A2(G131), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n203), .A2(new_n206), .A3(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n212), .A2(new_n215), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n210), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT88), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(G113), .B(G122), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n222), .B(G104), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n210), .A2(KEYINPUT88), .A3(new_n218), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n221), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(G131), .B1(new_n213), .B2(new_n214), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT17), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n226), .A2(new_n227), .A3(new_n207), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n209), .A2(KEYINPUT17), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n196), .A2(new_n197), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(new_n188), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(KEYINPUT69), .A3(new_n198), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n231), .A2(new_n234), .A3(new_n188), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n230), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n223), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n237), .A2(new_n238), .A3(new_n218), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n225), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(G475), .A2(G902), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT20), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT20), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n240), .A2(new_n244), .A3(new_n241), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G478), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n247), .A2(KEYINPUT15), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n202), .A2(G128), .ZN(new_n250));
  INV_X1    g064(.A(G128), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G143), .ZN(new_n252));
  INV_X1    g066(.A(G134), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n250), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G116), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G122), .ZN(new_n256));
  INV_X1    g070(.A(G122), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G116), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n259), .A2(G107), .ZN(new_n260));
  XNOR2_X1  g074(.A(G116), .B(G122), .ZN(new_n261));
  INV_X1    g075(.A(G107), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n254), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT13), .B1(new_n202), .B2(G128), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n265), .B1(new_n251), .B2(G143), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n202), .A2(KEYINPUT13), .A3(G128), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n253), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n250), .A2(new_n252), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G134), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT14), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n261), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n257), .A2(G116), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n262), .B1(new_n275), .B2(KEYINPUT14), .ZN(new_n276));
  AOI22_X1  g090(.A1(new_n254), .A2(new_n272), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT89), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n278), .B1(new_n259), .B2(G107), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n261), .A2(KEYINPUT89), .A3(new_n262), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT90), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n277), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n282), .B1(new_n277), .B2(new_n281), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n270), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(KEYINPUT9), .B(G234), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(G217), .A3(new_n200), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n277), .A2(new_n281), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT90), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n283), .ZN(new_n293));
  INV_X1    g107(.A(new_n289), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n293), .A2(new_n270), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n290), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G902), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n249), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  AOI211_X1 g112(.A(G902), .B(new_n248), .C1(new_n290), .C2(new_n295), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G952), .ZN(new_n301));
  AOI211_X1 g115(.A(G953), .B(new_n301), .C1(G234), .C2(G237), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  XNOR2_X1  g117(.A(KEYINPUT21), .B(G898), .ZN(new_n304));
  XOR2_X1   g118(.A(new_n304), .B(KEYINPUT91), .Z(new_n305));
  AOI211_X1 g119(.A(new_n297), .B(new_n200), .C1(G234), .C2(G237), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n303), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n238), .B1(new_n237), .B2(new_n218), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n212), .A2(new_n215), .A3(new_n217), .ZN(new_n310));
  AOI211_X1 g124(.A(new_n223), .B(new_n310), .C1(new_n230), .C2(new_n236), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n297), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G475), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n246), .A2(new_n300), .A3(new_n308), .A4(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT92), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n244), .B1(new_n240), .B2(new_n241), .ZN(new_n317));
  INV_X1    g131(.A(new_n241), .ZN(new_n318));
  AOI211_X1 g132(.A(KEYINPUT20), .B(new_n318), .C1(new_n225), .C2(new_n239), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n313), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n321), .A2(KEYINPUT92), .A3(new_n308), .A4(new_n300), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT2), .ZN(new_n324));
  INV_X1    g138(.A(G113), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(new_n325), .A3(KEYINPUT65), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT65), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n327), .B1(KEYINPUT2), .B2(G113), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(KEYINPUT2), .A2(G113), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(G116), .B(G119), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n329), .A2(new_n330), .A3(new_n332), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n262), .A2(KEYINPUT75), .A3(KEYINPUT3), .A4(G104), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n262), .A2(KEYINPUT75), .A3(G104), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT3), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n339), .B1(new_n262), .B2(G104), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n337), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G101), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G104), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT3), .B1(new_n344), .B2(G107), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n262), .A2(KEYINPUT75), .A3(G104), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(G101), .A3(new_n337), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n343), .A2(KEYINPUT4), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT4), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n347), .A2(new_n350), .A3(G101), .A4(new_n337), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n351), .A2(KEYINPUT76), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n351), .A2(KEYINPUT76), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n336), .B(new_n349), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(G110), .B(G122), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n262), .A2(G104), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n344), .A2(G107), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n342), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n358), .B1(new_n341), .B2(new_n342), .ZN(new_n359));
  INV_X1    g173(.A(G119), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G116), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n255), .A2(G119), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n362), .A3(KEYINPUT5), .ZN(new_n363));
  OR3_X1    g177(.A1(new_n255), .A2(KEYINPUT5), .A3(G119), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(new_n364), .A3(G113), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT79), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT79), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n363), .A2(new_n364), .A3(new_n367), .A4(G113), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n359), .A2(new_n366), .A3(new_n335), .A4(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n354), .A2(new_n355), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n188), .A2(G143), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n202), .A2(G146), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT0), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n374), .A2(new_n251), .ZN(new_n375));
  NOR2_X1   g189(.A1(KEYINPUT0), .A2(G128), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n373), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n371), .B(new_n372), .C1(new_n374), .C2(new_n251), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(G125), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT1), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n381), .B1(G143), .B2(new_n188), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n373), .B1(new_n382), .B2(new_n251), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT80), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n251), .A2(KEYINPUT1), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(new_n371), .A3(new_n372), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n383), .A2(new_n384), .A3(new_n191), .A4(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n251), .B1(new_n371), .B2(KEYINPUT1), .ZN(new_n388));
  XNOR2_X1  g202(.A(G143), .B(G146), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n191), .B(new_n386), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(KEYINPUT80), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n380), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT81), .ZN(new_n393));
  INV_X1    g207(.A(G224), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n393), .B1(new_n394), .B2(G953), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n200), .A2(KEYINPUT81), .A3(G224), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OR2_X1    g211(.A1(new_n397), .A2(KEYINPUT85), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(KEYINPUT85), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n392), .A2(KEYINPUT7), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT84), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n391), .A2(new_n401), .A3(new_n387), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n401), .B1(new_n391), .B2(new_n387), .ZN(new_n403));
  NOR3_X1   g217(.A1(new_n402), .A2(new_n403), .A3(new_n380), .ZN(new_n404));
  INV_X1    g218(.A(new_n397), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n405), .A2(KEYINPUT7), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n370), .B(new_n400), .C1(new_n404), .C2(new_n406), .ZN(new_n407));
  XOR2_X1   g221(.A(new_n355), .B(KEYINPUT8), .Z(new_n408));
  NAND3_X1  g222(.A1(new_n366), .A2(new_n335), .A3(new_n368), .ZN(new_n409));
  INV_X1    g223(.A(new_n358), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n343), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  OR2_X1    g226(.A1(new_n412), .A2(KEYINPUT83), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n359), .A2(new_n335), .A3(new_n365), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n414), .B1(new_n412), .B2(KEYINPUT83), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n408), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n297), .B1(new_n407), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT86), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OAI211_X1 g233(.A(KEYINPUT86), .B(new_n297), .C1(new_n407), .C2(new_n416), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n354), .A2(new_n369), .ZN(new_n422));
  INV_X1    g236(.A(new_n355), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(KEYINPUT6), .A3(new_n370), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT6), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n422), .A2(new_n426), .A3(new_n423), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n392), .B(new_n405), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n425), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT82), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT82), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n425), .A2(new_n431), .A3(new_n427), .A4(new_n428), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n421), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(G210), .B1(G237), .B2(G902), .ZN(new_n435));
  XOR2_X1   g249(.A(new_n435), .B(KEYINPUT87), .Z(new_n436));
  NAND2_X1  g250(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n421), .A2(new_n433), .A3(new_n435), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G221), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n440), .B1(new_n288), .B2(new_n297), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n377), .A2(new_n378), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n442), .B(new_n349), .C1(new_n352), .C2(new_n353), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT11), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n444), .B1(new_n253), .B2(G137), .ZN(new_n445));
  INV_X1    g259(.A(G137), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(KEYINPUT11), .A3(G134), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n253), .A2(G137), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n445), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G131), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n445), .A2(new_n447), .A3(new_n204), .A4(new_n448), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT10), .ZN(new_n454));
  AND3_X1   g268(.A1(new_n385), .A2(new_n371), .A3(new_n372), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT1), .B1(new_n202), .B2(G146), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT77), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT77), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n371), .A2(new_n458), .A3(KEYINPUT1), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n457), .A2(G128), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n455), .B1(new_n460), .B2(new_n373), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n454), .B1(new_n411), .B2(new_n461), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n456), .A2(G128), .B1(new_n371), .B2(new_n372), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n463), .A2(new_n455), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(new_n454), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n359), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n443), .A2(new_n453), .A3(new_n462), .A4(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(KEYINPUT78), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n251), .B1(new_n382), .B2(new_n458), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n389), .B1(new_n469), .B2(new_n457), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n359), .B1(new_n470), .B2(new_n455), .ZN(new_n471));
  AOI22_X1  g285(.A1(new_n471), .A2(new_n454), .B1(new_n465), .B2(new_n359), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT78), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n472), .A2(new_n473), .A3(new_n453), .A4(new_n443), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n468), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT12), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n386), .B1(new_n388), .B2(new_n389), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n477), .B1(new_n343), .B2(new_n410), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n460), .A2(new_n373), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n386), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n478), .B1(new_n359), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n476), .B1(new_n481), .B2(new_n453), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n411), .A2(new_n461), .ZN(new_n483));
  OAI211_X1 g297(.A(KEYINPUT12), .B(new_n452), .C1(new_n483), .C2(new_n478), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n475), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n200), .A2(G227), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(KEYINPUT74), .ZN(new_n488));
  XNOR2_X1  g302(.A(G110), .B(G140), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n488), .B(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n491), .B1(new_n468), .B2(new_n474), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n472), .A2(new_n443), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n452), .ZN(new_n494));
  AOI22_X1  g308(.A1(new_n486), .A2(new_n491), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(G469), .B1(new_n495), .B2(G902), .ZN(new_n496));
  INV_X1    g310(.A(G469), .ZN(new_n497));
  AOI221_X4 g311(.A(new_n491), .B1(new_n482), .B2(new_n484), .C1(new_n468), .C2(new_n474), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n490), .B1(new_n475), .B2(new_n494), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n497), .B(new_n297), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n441), .B1(new_n496), .B2(new_n500), .ZN(new_n501));
  AND4_X1   g315(.A1(new_n187), .A2(new_n323), .A3(new_n439), .A4(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT72), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n360), .A2(G128), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT68), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT68), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(new_n360), .A3(G128), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n251), .A2(G119), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n505), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(KEYINPUT24), .B(G110), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT23), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n512), .B1(new_n360), .B2(G128), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n251), .A2(KEYINPUT23), .A3(G119), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n504), .A3(new_n514), .ZN(new_n515));
  AOI22_X1  g329(.A1(new_n509), .A2(new_n511), .B1(G110), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n233), .A2(new_n235), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT70), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT70), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n233), .A2(new_n516), .A3(new_n519), .A4(new_n235), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n211), .A2(new_n188), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n198), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n515), .A2(G110), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n505), .A2(new_n507), .A3(new_n508), .ZN(new_n525));
  AOI22_X1  g339(.A1(new_n524), .A2(KEYINPUT71), .B1(new_n510), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT71), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n527), .B1(new_n515), .B2(G110), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n523), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n503), .B1(new_n521), .B2(new_n530), .ZN(new_n531));
  AOI211_X1 g345(.A(KEYINPUT72), .B(new_n529), .C1(new_n518), .C2(new_n520), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT22), .B(G137), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n200), .A2(G221), .A3(G234), .ZN(new_n534));
  XOR2_X1   g348(.A(new_n533), .B(new_n534), .Z(new_n535));
  NOR3_X1   g349(.A1(new_n531), .A2(new_n532), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n521), .A2(new_n530), .A3(new_n535), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n297), .ZN(new_n538));
  OAI21_X1  g352(.A(KEYINPUT25), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n521), .A2(new_n530), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(KEYINPUT72), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n521), .A2(new_n503), .A3(new_n530), .ZN(new_n542));
  INV_X1    g356(.A(new_n535), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT25), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n544), .A2(new_n545), .A3(new_n297), .A4(new_n537), .ZN(new_n546));
  INV_X1    g360(.A(G217), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n547), .B1(G234), .B2(new_n297), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n539), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT73), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT73), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n539), .A2(new_n546), .A3(new_n551), .A4(new_n548), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n544), .A2(new_n537), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n548), .A2(G902), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n550), .A2(new_n552), .A3(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(G472), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n253), .A2(G137), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n446), .A2(G134), .ZN(new_n559));
  OAI21_X1  g373(.A(G131), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n451), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n464), .A2(new_n561), .ZN(new_n562));
  AOI22_X1  g376(.A1(new_n450), .A2(new_n451), .B1(new_n377), .B2(new_n378), .ZN(new_n563));
  NOR3_X1   g377(.A1(new_n562), .A2(new_n563), .A3(new_n336), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT30), .ZN(new_n565));
  OR2_X1    g379(.A1(new_n565), .A2(KEYINPUT64), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(KEYINPUT64), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n566), .B(new_n567), .C1(new_n562), .C2(new_n563), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n452), .A2(new_n442), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n477), .A2(new_n451), .A3(new_n560), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n569), .A2(KEYINPUT64), .A3(new_n565), .A4(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n564), .B1(new_n572), .B2(new_n336), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n205), .A2(G210), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(KEYINPUT27), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT26), .B(G101), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT29), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n329), .A2(new_n330), .A3(new_n332), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n332), .B1(new_n329), .B2(new_n330), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n584), .B1(new_n569), .B2(new_n570), .ZN(new_n585));
  OAI21_X1  g399(.A(KEYINPUT28), .B1(new_n564), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(KEYINPUT67), .B1(new_n564), .B2(KEYINPUT28), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n569), .A2(new_n584), .A3(new_n570), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT67), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT28), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n586), .A2(new_n587), .A3(new_n591), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n580), .B(new_n581), .C1(new_n579), .C2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n592), .A2(new_n579), .ZN(new_n594));
  AOI21_X1  g408(.A(G902), .B1(new_n594), .B2(KEYINPUT29), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n557), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(G472), .A2(G902), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT66), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n598), .B1(new_n573), .B2(new_n578), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n584), .B1(new_n568), .B2(new_n571), .ZN(new_n600));
  NOR4_X1   g414(.A1(new_n600), .A2(KEYINPUT66), .A3(new_n564), .A4(new_n579), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT31), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n592), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n572), .A2(new_n336), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n605), .A2(new_n588), .A3(new_n578), .ZN(new_n606));
  OAI22_X1  g420(.A1(new_n604), .A2(new_n578), .B1(new_n606), .B2(KEYINPUT31), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n597), .B1(new_n603), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT32), .ZN(new_n609));
  INV_X1    g423(.A(new_n597), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n606), .A2(KEYINPUT66), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n573), .A2(new_n598), .A3(new_n578), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n611), .A2(KEYINPUT31), .A3(new_n612), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n600), .A2(new_n564), .A3(new_n579), .ZN(new_n614));
  AOI22_X1  g428(.A1(new_n614), .A2(new_n602), .B1(new_n592), .B2(new_n579), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n610), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT32), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n596), .B1(new_n609), .B2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n556), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n502), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G101), .ZN(G3));
  OAI21_X1  g436(.A(new_n297), .B1(new_n603), .B2(new_n607), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n616), .B1(new_n623), .B2(G472), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n501), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n625), .A2(new_n556), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n421), .A2(new_n435), .A3(new_n433), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n435), .B1(new_n421), .B2(new_n433), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n187), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(KEYINPUT93), .A2(KEYINPUT33), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n294), .B1(new_n293), .B2(new_n270), .ZN(new_n631));
  AOI211_X1 g445(.A(new_n269), .B(new_n289), .C1(new_n292), .C2(new_n283), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT93), .B(KEYINPUT33), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n290), .A2(new_n295), .A3(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n247), .A2(G902), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n633), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n297), .B1(new_n631), .B2(new_n632), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n247), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n320), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n308), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n629), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n626), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT94), .ZN(new_n645));
  XNOR2_X1  g459(.A(KEYINPUT34), .B(G104), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G6));
  NOR2_X1   g461(.A1(new_n320), .A2(new_n300), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n308), .B(KEYINPUT95), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n629), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n626), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT35), .B(G107), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G9));
  NOR2_X1   g468(.A1(new_n531), .A2(new_n532), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n543), .A2(KEYINPUT36), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n554), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n550), .A2(new_n552), .A3(new_n658), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n659), .A2(new_n624), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n502), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT37), .B(G110), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G12));
  INV_X1    g477(.A(new_n596), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n613), .A2(new_n615), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n617), .B1(new_n665), .B2(new_n597), .ZN(new_n666));
  AOI211_X1 g480(.A(KEYINPUT32), .B(new_n610), .C1(new_n613), .C2(new_n615), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n664), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n435), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n434), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n438), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n668), .A2(new_n671), .A3(new_n187), .A4(new_n501), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT96), .B(G900), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n302), .B1(new_n306), .B2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n648), .A2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n659), .A2(new_n677), .ZN(new_n678));
  OR2_X1    g492(.A1(new_n672), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G128), .ZN(G30));
  XOR2_X1   g494(.A(new_n674), .B(KEYINPUT39), .Z(new_n681));
  NAND2_X1  g495(.A1(new_n501), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT40), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n682), .A2(new_n683), .ZN(new_n686));
  OAI21_X1  g500(.A(KEYINPUT99), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n686), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT99), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n688), .A2(new_n689), .A3(new_n684), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n336), .B1(new_n562), .B2(new_n563), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n578), .B1(new_n691), .B2(new_n588), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT97), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n557), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n579), .B1(new_n564), .B2(new_n585), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(KEYINPUT97), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n599), .A2(new_n697), .A3(new_n601), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n557), .A2(new_n297), .ZN(new_n699));
  OAI21_X1  g513(.A(KEYINPUT98), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT98), .ZN(new_n701));
  INV_X1    g515(.A(new_n699), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n611), .A2(new_n612), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n701), .B(new_n702), .C1(new_n703), .C2(new_n697), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n705), .B1(new_n609), .B2(new_n618), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n706), .A2(new_n659), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n321), .A2(new_n300), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n187), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n439), .A2(KEYINPUT38), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n439), .A2(KEYINPUT38), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n687), .A2(new_n690), .A3(new_n707), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G143), .ZN(G45));
  NAND3_X1  g528(.A1(new_n320), .A2(new_n640), .A3(new_n675), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT100), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n320), .A2(new_n640), .A3(KEYINPUT100), .A4(new_n675), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n659), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n672), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(new_n188), .ZN(G48));
  INV_X1    g536(.A(new_n441), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n500), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n475), .A2(new_n494), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n491), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n475), .A2(new_n490), .A3(new_n485), .ZN(new_n727));
  AOI21_X1  g541(.A(G902), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g542(.A(KEYINPUT101), .B1(new_n728), .B2(new_n497), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n297), .B1(new_n498), .B2(new_n499), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT101), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n730), .A2(new_n731), .A3(G469), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n724), .B1(new_n729), .B2(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n620), .A2(new_n643), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(KEYINPUT102), .ZN(new_n735));
  XOR2_X1   g549(.A(KEYINPUT41), .B(G113), .Z(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G15));
  NAND3_X1  g551(.A1(new_n620), .A2(new_n651), .A3(new_n733), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G116), .ZN(G18));
  AND3_X1   g553(.A1(new_n659), .A2(new_n668), .A3(new_n323), .ZN(new_n740));
  INV_X1    g554(.A(new_n187), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n741), .B1(new_n670), .B2(new_n438), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n742), .A2(new_n733), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G119), .ZN(G21));
  OAI211_X1 g559(.A(new_n187), .B(new_n708), .C1(new_n627), .C2(new_n628), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n441), .B1(new_n728), .B2(new_n497), .ZN(new_n747));
  AOI22_X1  g561(.A1(new_n468), .A2(new_n474), .B1(new_n452), .B2(new_n493), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n727), .B1(new_n748), .B2(new_n490), .ZN(new_n749));
  AOI211_X1 g563(.A(KEYINPUT101), .B(new_n497), .C1(new_n749), .C2(new_n297), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n731), .B1(new_n730), .B2(G469), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n649), .B(new_n747), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n746), .A2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT103), .ZN(new_n754));
  AOI21_X1  g568(.A(G902), .B1(new_n613), .B2(new_n615), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n754), .B1(new_n755), .B2(new_n557), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n623), .A2(KEYINPUT103), .A3(G472), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n757), .A3(new_n608), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n758), .A2(new_n556), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n753), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G122), .ZN(G24));
  INV_X1    g575(.A(new_n720), .ZN(new_n762));
  INV_X1    g576(.A(new_n758), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(new_n743), .A3(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G125), .ZN(G27));
  INV_X1    g579(.A(KEYINPUT42), .ZN(new_n766));
  INV_X1    g580(.A(new_n436), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n767), .B1(new_n421), .B2(new_n433), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n627), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n719), .A2(new_n187), .A3(new_n769), .A4(new_n501), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n668), .A2(new_n552), .A3(new_n550), .A4(new_n555), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n766), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AOI22_X1  g586(.A1(new_n419), .A2(new_n420), .B1(new_n430), .B2(new_n432), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n438), .B(new_n187), .C1(new_n767), .C2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n717), .A2(new_n718), .ZN(new_n775));
  INV_X1    g589(.A(new_n500), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n486), .A2(new_n491), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n492), .A2(new_n494), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(G469), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(G469), .A2(G902), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n723), .B1(new_n776), .B2(new_n781), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n774), .A2(new_n775), .A3(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(KEYINPUT42), .A3(new_n620), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n772), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G131), .ZN(G33));
  NAND4_X1  g600(.A1(new_n769), .A2(new_n187), .A3(new_n501), .A4(new_n677), .ZN(new_n787));
  OAI21_X1  g601(.A(KEYINPUT104), .B1(new_n771), .B2(new_n787), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n774), .A2(new_n782), .A3(new_n676), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT104), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(new_n620), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G134), .ZN(G36));
  NAND2_X1  g607(.A1(new_n495), .A2(KEYINPUT45), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT45), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n475), .A2(new_n494), .A3(new_n490), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n490), .B1(new_n475), .B2(new_n485), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n794), .A2(G469), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n780), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT46), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n776), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT105), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n799), .A2(new_n803), .A3(KEYINPUT46), .A4(new_n780), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n799), .A2(KEYINPUT46), .A3(new_n780), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(KEYINPUT105), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n802), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n723), .ZN(new_n808));
  INV_X1    g622(.A(new_n681), .ZN(new_n809));
  OAI21_X1  g623(.A(KEYINPUT106), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT106), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n807), .A2(new_n811), .A3(new_n723), .A4(new_n681), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n321), .A2(new_n640), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(KEYINPUT43), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(new_n624), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n816), .A2(KEYINPUT44), .A3(new_n659), .ZN(new_n817));
  AOI21_X1  g631(.A(KEYINPUT44), .B1(new_n816), .B2(new_n659), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n818), .A2(new_n774), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n813), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G137), .ZN(G39));
  INV_X1    g635(.A(new_n774), .ZN(new_n822));
  AND4_X1   g636(.A1(new_n556), .A2(new_n822), .A3(new_n619), .A4(new_n719), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT47), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n808), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT47), .B1(new_n807), .B2(new_n723), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n823), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(G140), .ZN(G42));
  AND2_X1   g642(.A1(new_n710), .A2(new_n711), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n706), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT49), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n729), .A2(new_n732), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(new_n500), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n830), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  NOR4_X1   g649(.A1(new_n556), .A2(new_n741), .A3(new_n441), .A4(new_n814), .ZN(new_n836));
  XOR2_X1   g650(.A(new_n836), .B(KEYINPUT107), .Z(new_n837));
  OAI211_X1 g651(.A(new_n835), .B(new_n837), .C1(new_n831), .C2(new_n834), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n815), .A2(new_n303), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n839), .A2(new_n759), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n840), .A2(new_n741), .A3(new_n829), .A4(new_n733), .ZN(new_n841));
  XOR2_X1   g655(.A(new_n841), .B(KEYINPUT50), .Z(new_n842));
  AND2_X1   g656(.A1(new_n840), .A2(new_n822), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n808), .B(new_n824), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n833), .A2(new_n723), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n700), .B(new_n704), .C1(new_n666), .C2(new_n667), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n847), .A2(new_n556), .A3(new_n303), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n822), .A2(new_n733), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT112), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n320), .A2(new_n640), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n550), .A2(new_n552), .A3(new_n658), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n854), .A2(new_n758), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n849), .A2(new_n839), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n853), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n851), .B1(new_n850), .B2(new_n852), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n842), .B(new_n846), .C1(new_n860), .C2(KEYINPUT113), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(KEYINPUT51), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT111), .ZN(new_n863));
  OAI22_X1  g677(.A1(new_n844), .A2(new_n863), .B1(new_n723), .B2(new_n833), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n825), .A2(new_n826), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n865), .A2(KEYINPUT111), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n843), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n841), .B(KEYINPUT50), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(KEYINPUT51), .ZN(new_n869));
  AOI22_X1  g683(.A1(new_n867), .A2(new_n869), .B1(KEYINPUT113), .B2(KEYINPUT51), .ZN(new_n870));
  INV_X1    g684(.A(new_n860), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n862), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n857), .A2(new_n771), .ZN(new_n873));
  XOR2_X1   g687(.A(new_n873), .B(KEYINPUT48), .Z(new_n874));
  NAND2_X1  g688(.A1(new_n850), .A2(new_n641), .ZN(new_n875));
  AOI211_X1 g689(.A(new_n301), .B(G953), .C1(new_n840), .C2(new_n743), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n877), .B(KEYINPUT114), .Z(new_n878));
  NAND2_X1  g692(.A1(new_n872), .A2(new_n878), .ZN(new_n879));
  NOR4_X1   g693(.A1(new_n320), .A2(new_n298), .A3(new_n299), .A4(new_n674), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n437), .A2(new_n880), .A3(new_n187), .A4(new_n438), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n854), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n619), .A2(new_n782), .ZN(new_n883));
  AOI22_X1  g697(.A1(new_n783), .A2(new_n855), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n785), .A2(new_n792), .A3(new_n884), .ZN(new_n885));
  AOI22_X1  g699(.A1(new_n743), .A2(new_n740), .B1(new_n753), .B2(new_n759), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n769), .A2(new_n741), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n641), .A2(new_n648), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n626), .A2(new_n887), .A3(new_n649), .A4(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n502), .B1(new_n620), .B2(new_n660), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n620), .B(new_n733), .C1(new_n643), .C2(new_n651), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n886), .A2(new_n890), .A3(new_n891), .A4(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n885), .A2(new_n893), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n629), .A2(new_n619), .A3(new_n782), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n501), .A2(new_n675), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n746), .A2(new_n896), .ZN(new_n897));
  AOI22_X1  g711(.A1(new_n762), .A2(new_n895), .B1(new_n897), .B2(new_n707), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n898), .A2(KEYINPUT108), .A3(new_n679), .A4(new_n764), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT108), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n742), .A2(new_n719), .A3(new_n659), .A4(new_n733), .ZN(new_n901));
  OAI22_X1  g715(.A1(new_n901), .A2(new_n758), .B1(new_n672), .B2(new_n678), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n854), .A2(new_n847), .ZN(new_n903));
  AOI211_X1 g717(.A(new_n441), .B(new_n674), .C1(new_n496), .C2(new_n500), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n742), .A2(new_n708), .A3(new_n904), .ZN(new_n905));
  OAI22_X1  g719(.A1(new_n903), .A2(new_n905), .B1(new_n672), .B2(new_n720), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n900), .B1(new_n902), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n899), .A2(new_n907), .A3(KEYINPUT52), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n894), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT52), .B1(new_n899), .B2(new_n907), .ZN(new_n910));
  OAI21_X1  g724(.A(KEYINPUT53), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n899), .A2(new_n907), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT52), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT53), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT52), .B1(new_n902), .B2(new_n906), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n914), .A2(new_n915), .A3(new_n894), .A4(new_n916), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n911), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT109), .B1(new_n918), .B2(KEYINPUT54), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n915), .B1(new_n909), .B2(new_n910), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT54), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n891), .A2(KEYINPUT53), .A3(new_n890), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n885), .A2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT110), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n886), .A2(new_n924), .A3(new_n892), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n924), .B1(new_n886), .B2(new_n892), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n914), .A2(new_n916), .A3(new_n923), .A4(new_n927), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n920), .A2(new_n921), .A3(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n919), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n918), .A2(KEYINPUT109), .A3(KEYINPUT54), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n879), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(G952), .A2(G953), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT115), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n838), .B1(new_n933), .B2(new_n935), .ZN(G75));
  XNOR2_X1  g750(.A(new_n428), .B(KEYINPUT117), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT55), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n425), .A2(new_n427), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT116), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n938), .B(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n920), .A2(new_n928), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(G902), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(G210), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT56), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n941), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n200), .A2(G952), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT118), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n943), .A2(new_n767), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n941), .A2(new_n946), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n947), .A2(new_n952), .ZN(G51));
  XNOR2_X1  g767(.A(new_n799), .B(KEYINPUT120), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n943), .A2(new_n954), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n780), .B(KEYINPUT57), .Z(new_n956));
  AOI21_X1  g770(.A(new_n921), .B1(new_n920), .B2(new_n928), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n956), .B1(new_n929), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n749), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT119), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n955), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n958), .A2(KEYINPUT119), .A3(new_n749), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n948), .B1(new_n961), .B2(new_n962), .ZN(G54));
  AND2_X1   g777(.A1(KEYINPUT58), .A2(G475), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n944), .A2(new_n240), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n240), .B1(new_n944), .B2(new_n964), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n965), .A2(new_n966), .A3(new_n948), .ZN(G60));
  NOR2_X1   g781(.A1(new_n929), .A2(new_n957), .ZN(new_n968));
  NAND2_X1  g782(.A1(G478), .A2(G902), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT59), .Z(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n633), .A2(new_n635), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n949), .B1(new_n968), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n931), .A2(new_n932), .A3(new_n971), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n633), .A2(new_n635), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n973), .B1(new_n974), .B2(new_n975), .ZN(G63));
  XNOR2_X1  g790(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n977));
  NAND2_X1  g791(.A1(G217), .A2(G902), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n977), .B(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n979), .B1(new_n920), .B2(new_n928), .ZN(new_n980));
  OR2_X1    g794(.A1(new_n980), .A2(new_n553), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n657), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n981), .A2(new_n949), .A3(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT61), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n983), .B(new_n984), .ZN(G66));
  INV_X1    g799(.A(new_n305), .ZN(new_n986));
  OAI21_X1  g800(.A(G953), .B1(new_n986), .B2(new_n394), .ZN(new_n987));
  INV_X1    g801(.A(new_n893), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n987), .B1(new_n988), .B2(G953), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n940), .B1(G898), .B2(new_n200), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n989), .B(new_n990), .ZN(G69));
  INV_X1    g805(.A(KEYINPUT124), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n193), .A2(new_n194), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n572), .B(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT122), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n995), .B1(new_n902), .B2(new_n721), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n762), .A2(new_n895), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n764), .A2(new_n679), .A3(new_n997), .A4(KEYINPUT122), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT62), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n713), .A2(new_n996), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  OR4_X1    g814(.A1(new_n771), .A2(new_n682), .A3(new_n774), .A4(new_n888), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n820), .A2(new_n1000), .A3(new_n827), .A4(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT123), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n713), .A2(new_n996), .A3(new_n998), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1003), .B1(new_n1004), .B2(KEYINPUT62), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1005), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n1004), .A2(new_n1003), .A3(KEYINPUT62), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1002), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  OAI211_X1 g822(.A(new_n992), .B(new_n994), .C1(new_n1008), .C2(G953), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n200), .B1(G227), .B2(G900), .ZN(new_n1010));
  AND2_X1   g824(.A1(new_n820), .A2(new_n827), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n813), .A2(new_n620), .A3(new_n742), .A4(new_n708), .ZN(new_n1012));
  AND4_X1   g826(.A1(new_n785), .A2(new_n996), .A3(new_n998), .A4(new_n792), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n1011), .A2(new_n200), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n994), .B1(G900), .B2(G953), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1010), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1009), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1007), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1018), .A2(new_n1005), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n200), .B1(new_n1019), .B2(new_n1002), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n992), .B1(new_n1020), .B2(new_n994), .ZN(new_n1021));
  OAI21_X1  g835(.A(KEYINPUT125), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n994), .B1(new_n1008), .B2(G953), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1023), .A2(KEYINPUT124), .ZN(new_n1024));
  INV_X1    g838(.A(KEYINPUT125), .ZN(new_n1025));
  NAND4_X1  g839(.A1(new_n1024), .A2(new_n1025), .A3(new_n1009), .A4(new_n1016), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1022), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g841(.A(new_n1023), .ZN(new_n1028));
  AND2_X1   g842(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1010), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1027), .A2(new_n1030), .ZN(G72));
  NAND2_X1  g845(.A1(new_n1008), .A2(new_n988), .ZN(new_n1032));
  XOR2_X1   g846(.A(new_n699), .B(KEYINPUT63), .Z(new_n1033));
  INV_X1    g847(.A(new_n1033), .ZN(new_n1034));
  AOI211_X1 g848(.A(new_n573), .B(new_n579), .C1(new_n1032), .C2(new_n1034), .ZN(new_n1035));
  AND4_X1   g849(.A1(new_n988), .A2(new_n1011), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1036));
  OAI211_X1 g850(.A(new_n573), .B(new_n579), .C1(new_n1036), .C2(new_n1033), .ZN(new_n1037));
  XOR2_X1   g851(.A(new_n580), .B(KEYINPUT126), .Z(new_n1038));
  INV_X1    g852(.A(new_n703), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n1033), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n948), .B1(new_n918), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1037), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g856(.A(KEYINPUT127), .B1(new_n1035), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1044));
  NAND3_X1  g858(.A1(new_n1044), .A2(new_n574), .A3(new_n578), .ZN(new_n1045));
  INV_X1    g859(.A(KEYINPUT127), .ZN(new_n1046));
  NAND4_X1  g860(.A1(new_n1045), .A2(new_n1046), .A3(new_n1037), .A4(new_n1041), .ZN(new_n1047));
  NAND2_X1  g861(.A1(new_n1043), .A2(new_n1047), .ZN(G57));
endmodule


