//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n187));
  XNOR2_X1  g001(.A(G110), .B(G140), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT78), .ZN(new_n189));
  XOR2_X1   g003(.A(KEYINPUT70), .B(G953), .Z(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G227), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n189), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT12), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT3), .ZN(new_n194));
  INV_X1    g008(.A(G104), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n194), .B1(new_n195), .B2(G107), .ZN(new_n196));
  INV_X1    g010(.A(G107), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(KEYINPUT3), .A3(G104), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G101), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT79), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n201), .B1(new_n197), .B2(G104), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n195), .A2(KEYINPUT79), .A3(G107), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n199), .A2(new_n200), .A3(new_n202), .A4(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT83), .B1(new_n197), .B2(G104), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT83), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(new_n195), .A3(G107), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n197), .A2(G104), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G101), .ZN(new_n210));
  AND2_X1   g024(.A1(new_n204), .A2(new_n210), .ZN(new_n211));
  OR2_X1    g025(.A1(KEYINPUT64), .A2(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(KEYINPUT64), .A2(G143), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n212), .A2(KEYINPUT65), .A3(G146), .A4(new_n213), .ZN(new_n214));
  AND2_X1   g028(.A1(KEYINPUT64), .A2(G143), .ZN(new_n215));
  NOR2_X1   g029(.A1(KEYINPUT64), .A2(G143), .ZN(new_n216));
  INV_X1    g030(.A(G146), .ZN(new_n217));
  NOR3_X1   g031(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n219));
  INV_X1    g033(.A(G143), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n219), .B1(new_n220), .B2(G146), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n214), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G128), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n217), .B1(new_n215), .B2(new_n216), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n223), .B1(new_n224), .B2(KEYINPUT1), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  AND2_X1   g040(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n227));
  NOR2_X1   g041(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G128), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n212), .A2(G146), .A3(new_n213), .ZN(new_n231));
  INV_X1    g045(.A(new_n221), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n230), .B1(new_n233), .B2(new_n214), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n211), .B1(new_n226), .B2(new_n234), .ZN(new_n235));
  NOR3_X1   g049(.A1(new_n227), .A2(new_n228), .A3(new_n223), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n215), .A2(new_n216), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n221), .B1(new_n237), .B2(G146), .ZN(new_n238));
  NOR4_X1   g052(.A1(new_n215), .A2(new_n216), .A3(new_n219), .A4(new_n217), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n236), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n204), .A2(new_n210), .ZN(new_n241));
  OAI22_X1  g055(.A1(new_n227), .A2(new_n228), .B1(new_n220), .B2(G146), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G128), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n220), .A2(G146), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n224), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n240), .A2(new_n241), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n235), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G134), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G137), .ZN(new_n250));
  INV_X1    g064(.A(G137), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(KEYINPUT11), .A3(G134), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT11), .B1(new_n251), .B2(G134), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n250), .B(new_n252), .C1(new_n253), .C2(KEYINPUT66), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT11), .ZN(new_n255));
  OAI211_X1 g069(.A(KEYINPUT66), .B(new_n255), .C1(new_n249), .C2(G137), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(G131), .B1(new_n254), .B2(new_n257), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n252), .A2(new_n250), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT66), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n249), .A2(G137), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n260), .B1(new_n261), .B2(KEYINPUT11), .ZN(new_n262));
  INV_X1    g076(.A(G131), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n259), .A2(new_n262), .A3(new_n263), .A4(new_n256), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n258), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n193), .B1(new_n248), .B2(new_n265), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n258), .A2(new_n264), .ZN(new_n267));
  AOI211_X1 g081(.A(KEYINPUT12), .B(new_n267), .C1(new_n235), .C2(new_n247), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT84), .B(KEYINPUT10), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n240), .A2(new_n246), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n204), .A2(new_n210), .A3(KEYINPUT10), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n235), .A2(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AND3_X1   g088(.A1(new_n197), .A2(KEYINPUT3), .A3(G104), .ZN(new_n275));
  AOI21_X1  g089(.A(KEYINPUT3), .B1(new_n197), .B2(G104), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n202), .B(new_n203), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT80), .ZN(new_n278));
  AND3_X1   g092(.A1(new_n277), .A2(new_n278), .A3(G101), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n278), .B1(new_n277), .B2(G101), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n204), .A2(KEYINPUT4), .ZN(new_n281));
  NOR3_X1   g095(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(KEYINPUT0), .A2(G128), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n284), .B1(new_n238), .B2(new_n239), .ZN(new_n285));
  OR2_X1    g099(.A1(KEYINPUT0), .A2(G128), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n283), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n287), .B1(new_n224), .B2(new_n244), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(KEYINPUT81), .B(KEYINPUT4), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n277), .A2(G101), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n285), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  NOR3_X1   g106(.A1(new_n282), .A2(KEYINPUT82), .A3(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT82), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n277), .A2(G101), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT80), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n277), .A2(new_n278), .A3(G101), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n296), .A2(KEYINPUT4), .A3(new_n297), .A4(new_n204), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n285), .A2(new_n289), .A3(new_n291), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n294), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n267), .B(new_n274), .C1(new_n293), .C2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n192), .B1(new_n269), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n301), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT82), .B1(new_n282), .B2(new_n292), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n298), .A2(new_n299), .A3(new_n294), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n267), .B1(new_n306), .B2(new_n274), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n302), .B1(new_n308), .B2(new_n192), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n187), .B(G469), .C1(new_n309), .C2(G902), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n269), .A2(new_n301), .ZN(new_n311));
  INV_X1    g125(.A(new_n192), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n274), .B1(new_n293), .B2(new_n300), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n265), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(new_n301), .A3(new_n192), .ZN(new_n316));
  AOI21_X1  g130(.A(G902), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G469), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT85), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G902), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n192), .B1(new_n315), .B2(new_n301), .ZN(new_n321));
  AND3_X1   g135(.A1(new_n269), .A2(new_n301), .A3(new_n192), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n318), .B(new_n320), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n310), .A2(new_n319), .A3(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT9), .B(G234), .ZN(new_n325));
  OAI21_X1  g139(.A(G221), .B1(new_n325), .B2(G902), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(G214), .B1(G237), .B2(G902), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT2), .B(G113), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  OR2_X1    g145(.A1(KEYINPUT68), .A2(G119), .ZN(new_n332));
  NAND2_X1  g146(.A1(KEYINPUT68), .A2(G119), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(G116), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(G119), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n331), .B(new_n334), .C1(G116), .C2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n333), .ZN(new_n337));
  NOR2_X1   g151(.A1(KEYINPUT68), .A2(G119), .ZN(new_n338));
  INV_X1    g152(.A(G116), .ZN(new_n339));
  NOR3_X1   g153(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n335), .A2(G116), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n330), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n336), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n297), .A2(KEYINPUT4), .A3(new_n204), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n343), .B(new_n291), .C1(new_n344), .C2(new_n280), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT5), .ZN(new_n346));
  NOR3_X1   g160(.A1(new_n340), .A2(new_n346), .A3(new_n341), .ZN(new_n347));
  OAI21_X1  g161(.A(G113), .B1(new_n334), .B2(KEYINPUT5), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n211), .B(new_n336), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(G110), .B(G122), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n345), .A2(new_n351), .A3(new_n349), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(KEYINPUT6), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n283), .B1(new_n233), .B2(new_n214), .ZN(new_n356));
  OAI21_X1  g170(.A(G125), .B1(new_n356), .B2(new_n288), .ZN(new_n357));
  INV_X1    g171(.A(G125), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n240), .A2(new_n246), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G224), .ZN(new_n361));
  OR2_X1    g175(.A1(new_n361), .A2(G953), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n362), .B(KEYINPUT86), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n360), .B(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT6), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n350), .A2(new_n365), .A3(new_n352), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n355), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  XOR2_X1   g181(.A(new_n351), .B(KEYINPUT8), .Z(new_n368));
  OAI21_X1  g182(.A(new_n336), .B1(new_n347), .B2(new_n348), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n241), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n368), .B1(new_n349), .B2(new_n370), .ZN(new_n371));
  AND4_X1   g185(.A1(KEYINPUT7), .A2(new_n357), .A3(new_n359), .A4(new_n362), .ZN(new_n372));
  AOI22_X1  g186(.A1(new_n357), .A2(new_n359), .B1(KEYINPUT7), .B2(new_n362), .ZN(new_n373));
  NOR3_X1   g187(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(G902), .B1(new_n374), .B2(new_n354), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n367), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(G210), .B1(G237), .B2(G902), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n377), .B(KEYINPUT87), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n378), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n367), .A2(new_n375), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n329), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n327), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT20), .ZN(new_n385));
  INV_X1    g199(.A(G140), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G125), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n358), .A2(G140), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n388), .A3(KEYINPUT16), .ZN(new_n389));
  OR3_X1    g203(.A1(new_n358), .A2(KEYINPUT16), .A3(G140), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n390), .A3(G146), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(KEYINPUT75), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n389), .A2(new_n390), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n217), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT75), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n389), .A2(new_n390), .A3(new_n395), .A4(G146), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n392), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT89), .ZN(new_n398));
  INV_X1    g212(.A(G237), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n190), .A2(G143), .A3(G214), .A4(new_n399), .ZN(new_n400));
  OR2_X1    g214(.A1(KEYINPUT70), .A2(G953), .ZN(new_n401));
  NAND2_X1  g215(.A1(KEYINPUT70), .A2(G953), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n401), .A2(G214), .A3(new_n399), .A4(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n237), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n398), .B1(new_n405), .B2(new_n263), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n400), .A2(new_n404), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(KEYINPUT89), .A3(G131), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n397), .B1(new_n409), .B2(KEYINPUT17), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT17), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n405), .A2(new_n263), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n406), .A2(new_n411), .A3(new_n408), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(KEYINPUT91), .ZN(new_n414));
  AOI21_X1  g228(.A(KEYINPUT89), .B1(new_n407), .B2(G131), .ZN(new_n415));
  AOI211_X1 g229(.A(new_n398), .B(new_n263), .C1(new_n400), .C2(new_n404), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT91), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n417), .A2(new_n418), .A3(new_n411), .A4(new_n412), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n410), .A2(new_n414), .A3(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(G113), .B(G122), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n421), .B(new_n195), .ZN(new_n422));
  NAND2_X1  g236(.A1(KEYINPUT18), .A2(G131), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n405), .A2(KEYINPUT88), .A3(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT88), .ZN(new_n425));
  OAI211_X1 g239(.A(KEYINPUT18), .B(G131), .C1(new_n407), .C2(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(G125), .B(G140), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n427), .B(new_n217), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n424), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n420), .A2(new_n422), .A3(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n422), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT90), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n427), .A2(new_n432), .ZN(new_n433));
  XOR2_X1   g247(.A(new_n433), .B(KEYINPUT19), .Z(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n391), .B1(new_n435), .B2(G146), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n436), .B1(new_n417), .B2(new_n412), .ZN(new_n437));
  INV_X1    g251(.A(new_n429), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n431), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n430), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(G475), .A2(G902), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n385), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n441), .ZN(new_n443));
  AOI211_X1 g257(.A(KEYINPUT20), .B(new_n443), .C1(new_n430), .C2(new_n439), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n422), .B1(new_n420), .B2(new_n429), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(G902), .B1(new_n446), .B2(new_n430), .ZN(new_n447));
  INV_X1    g261(.A(G475), .ZN(new_n448));
  OAI22_X1  g262(.A1(new_n442), .A2(new_n444), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(G116), .B(G122), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n450), .B(new_n197), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n212), .A2(G128), .A3(new_n213), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n220), .A2(G128), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n452), .A2(new_n249), .A3(new_n454), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n452), .A2(KEYINPUT13), .A3(new_n454), .ZN(new_n456));
  OAI21_X1  g270(.A(G134), .B1(new_n452), .B2(KEYINPUT13), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n451), .B(new_n455), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  NOR3_X1   g272(.A1(new_n215), .A2(new_n216), .A3(new_n223), .ZN(new_n459));
  OAI21_X1  g273(.A(G134), .B1(new_n459), .B2(new_n453), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n455), .ZN(new_n461));
  INV_X1    g275(.A(G122), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(G116), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n197), .B1(new_n463), .B2(KEYINPUT14), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(new_n450), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(G217), .ZN(new_n467));
  NOR3_X1   g281(.A1(new_n325), .A2(new_n467), .A3(G953), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n458), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(KEYINPUT92), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT92), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n458), .A2(new_n466), .A3(new_n471), .A4(new_n468), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n458), .A2(new_n466), .ZN(new_n473));
  INV_X1    g287(.A(new_n468), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n470), .A2(new_n472), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(G478), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n477), .A2(KEYINPUT15), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n476), .A2(new_n320), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT94), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n476), .A2(KEYINPUT94), .A3(new_n320), .A4(new_n479), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n476), .A2(KEYINPUT93), .A3(new_n320), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(KEYINPUT93), .B1(new_n476), .B2(new_n320), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n484), .B1(new_n478), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(G952), .ZN(new_n490));
  AOI211_X1 g304(.A(G953), .B(new_n490), .C1(G234), .C2(G237), .ZN(new_n491));
  AOI211_X1 g305(.A(new_n320), .B(new_n190), .C1(G234), .C2(G237), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(KEYINPUT95), .ZN(new_n493));
  XNOR2_X1  g307(.A(KEYINPUT21), .B(G898), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n491), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n489), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n449), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n384), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(G472), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n288), .B1(new_n222), .B2(new_n284), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n265), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n250), .ZN(new_n503));
  OAI21_X1  g317(.A(G131), .B1(new_n503), .B2(new_n261), .ZN(new_n504));
  AOI22_X1  g318(.A1(G128), .A2(new_n242), .B1(new_n224), .B2(new_n244), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n504), .B(new_n264), .C1(new_n234), .C2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT30), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n502), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n507), .B1(new_n502), .B2(new_n506), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n343), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n343), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n502), .A2(new_n506), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT69), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n502), .A2(new_n506), .A3(KEYINPUT69), .A4(new_n511), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n190), .A2(G210), .A3(new_n399), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n516), .B(KEYINPUT27), .ZN(new_n517));
  XNOR2_X1  g331(.A(KEYINPUT26), .B(G101), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n517), .B(new_n518), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n510), .A2(new_n514), .A3(new_n515), .A4(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT31), .ZN(new_n521));
  AND2_X1   g335(.A1(new_n514), .A2(new_n515), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT31), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n522), .A2(new_n523), .A3(new_n519), .A4(new_n510), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT28), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n512), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n502), .A2(new_n506), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n343), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n514), .A2(new_n530), .A3(new_n515), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n528), .B1(new_n531), .B2(KEYINPUT28), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n532), .A2(new_n519), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n500), .B(new_n320), .C1(new_n525), .C2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT32), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n521), .B(new_n524), .C1(new_n532), .C2(new_n519), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT32), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n536), .A2(new_n537), .A3(new_n500), .A4(new_n320), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT72), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n519), .A2(KEYINPUT29), .ZN(new_n541));
  AOI211_X1 g355(.A(new_n528), .B(new_n541), .C1(new_n531), .C2(KEYINPUT28), .ZN(new_n542));
  OAI21_X1  g356(.A(KEYINPUT71), .B1(new_n542), .B2(G902), .ZN(new_n543));
  INV_X1    g357(.A(new_n519), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n522), .A2(new_n544), .A3(new_n510), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n545), .B1(new_n532), .B2(new_n544), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT29), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n544), .A2(new_n547), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n532), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT71), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n550), .A2(new_n551), .A3(new_n320), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n543), .A2(new_n548), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(G472), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n539), .A2(new_n540), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n540), .B1(new_n539), .B2(new_n554), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n467), .B1(G234), .B2(new_n320), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n427), .A2(new_n217), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n391), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n332), .A2(G128), .A3(new_n333), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n223), .A2(KEYINPUT23), .A3(G119), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(G110), .ZN(new_n565));
  AOI21_X1  g379(.A(G128), .B1(new_n332), .B2(new_n333), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n564), .B(new_n565), .C1(KEYINPUT23), .C2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT73), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n332), .A2(new_n568), .A3(G128), .A4(new_n333), .ZN(new_n569));
  NOR3_X1   g383(.A1(new_n337), .A2(new_n338), .A3(new_n223), .ZN(new_n570));
  OAI21_X1  g384(.A(KEYINPUT73), .B1(new_n335), .B2(G128), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n565), .A2(KEYINPUT24), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT24), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(G110), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT74), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n572), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n575), .B1(new_n572), .B2(new_n574), .ZN(new_n577));
  OAI221_X1 g391(.A(new_n569), .B1(new_n570), .B2(new_n571), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n561), .B1(new_n567), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n576), .A2(new_n577), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n332), .A2(new_n333), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT23), .B1(new_n584), .B2(new_n223), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n562), .A2(new_n563), .ZN(new_n586));
  OAI21_X1  g400(.A(G110), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AND4_X1   g401(.A1(KEYINPUT76), .A2(new_n397), .A3(new_n583), .A4(new_n587), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n562), .B(new_n563), .C1(new_n566), .C2(KEYINPUT23), .ZN(new_n589));
  AOI22_X1  g403(.A1(G110), .A2(new_n589), .B1(new_n581), .B2(new_n582), .ZN(new_n590));
  AOI21_X1  g404(.A(KEYINPUT76), .B1(new_n590), .B2(new_n397), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n580), .B1(new_n588), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n593));
  XNOR2_X1  g407(.A(KEYINPUT22), .B(G137), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT76), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n392), .A2(new_n394), .A3(new_n396), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n583), .A2(new_n587), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n590), .A2(KEYINPUT76), .A3(new_n397), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n603), .A2(new_n580), .A3(new_n595), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n597), .A2(new_n320), .A3(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT25), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n597), .A2(KEYINPUT25), .A3(new_n604), .A4(new_n320), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n559), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n595), .B1(new_n603), .B2(new_n580), .ZN(new_n610));
  AOI211_X1 g424(.A(new_n579), .B(new_n596), .C1(new_n601), .C2(new_n602), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n558), .A2(G902), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(KEYINPUT77), .B1(new_n557), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT77), .ZN(new_n617));
  INV_X1    g431(.A(new_n615), .ZN(new_n618));
  NOR4_X1   g432(.A1(new_n555), .A2(new_n556), .A3(new_n617), .A4(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n499), .B1(new_n616), .B2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(G101), .ZN(G3));
  NAND2_X1  g435(.A1(new_n536), .A2(new_n320), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(G472), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n623), .A2(new_n534), .ZN(new_n624));
  AND4_X1   g438(.A1(new_n615), .A2(new_n624), .A3(new_n326), .A4(new_n324), .ZN(new_n625));
  INV_X1    g439(.A(new_n487), .ZN(new_n626));
  AOI21_X1  g440(.A(G478), .B1(new_n626), .B2(new_n485), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n458), .A2(new_n466), .A3(KEYINPUT96), .A4(new_n468), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n475), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT96), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n469), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g445(.A(KEYINPUT33), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT33), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n470), .A2(new_n475), .A3(new_n633), .A4(new_n472), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n477), .B1(new_n635), .B2(new_n320), .ZN(new_n636));
  OAI21_X1  g450(.A(KEYINPUT97), .B1(new_n627), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n477), .B1(new_n486), .B2(new_n487), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT97), .ZN(new_n639));
  AOI21_X1  g453(.A(G902), .B1(new_n632), .B2(new_n634), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n638), .B(new_n639), .C1(new_n477), .C2(new_n640), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n449), .ZN(new_n643));
  INV_X1    g457(.A(new_n381), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n380), .B1(new_n367), .B2(new_n375), .ZN(new_n645));
  OAI211_X1 g459(.A(new_n496), .B(new_n328), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n625), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT98), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT34), .B(G104), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G6));
  NAND2_X1  g465(.A1(new_n440), .A2(new_n441), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(KEYINPUT20), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT99), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n440), .A2(new_n385), .A3(new_n441), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n444), .A2(KEYINPUT99), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n646), .ZN(new_n660));
  INV_X1    g474(.A(new_n430), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n320), .B1(new_n661), .B2(new_n445), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n489), .B1(G475), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n659), .A2(new_n660), .A3(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n625), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT35), .B(G107), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G9));
  AOI21_X1  g482(.A(KEYINPUT25), .B1(new_n612), .B2(new_n320), .ZN(new_n669));
  INV_X1    g483(.A(new_n608), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n558), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT100), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n596), .A2(KEYINPUT36), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n592), .B(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n613), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n671), .A2(new_n672), .A3(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n675), .ZN(new_n677));
  OAI21_X1  g491(.A(KEYINPUT100), .B1(new_n609), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n384), .A2(new_n498), .A3(new_n624), .A4(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT37), .B(G110), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G12));
  NAND2_X1  g497(.A1(new_n539), .A2(new_n554), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(KEYINPUT72), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n310), .A2(new_n319), .A3(new_n323), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n676), .A2(new_n678), .A3(new_n382), .ZN(new_n687));
  INV_X1    g501(.A(new_n326), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  AOI22_X1  g503(.A1(new_n535), .A2(new_n538), .B1(new_n553), .B2(G472), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n540), .ZN(new_n691));
  INV_X1    g505(.A(G900), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n491), .B1(new_n493), .B2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  AND4_X1   g508(.A1(new_n657), .A2(new_n663), .A3(new_n656), .A4(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n685), .A2(new_n689), .A3(new_n691), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G128), .ZN(G30));
  INV_X1    g511(.A(new_n327), .ZN(new_n698));
  XOR2_X1   g512(.A(new_n693), .B(KEYINPUT39), .Z(new_n699));
  NAND3_X1  g513(.A1(new_n698), .A2(KEYINPUT40), .A3(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(KEYINPUT40), .B1(new_n698), .B2(new_n699), .ZN(new_n702));
  OAI21_X1  g516(.A(KEYINPUT102), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n702), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT102), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n704), .A2(new_n705), .A3(new_n700), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n644), .A2(new_n645), .ZN(new_n707));
  XOR2_X1   g521(.A(new_n707), .B(KEYINPUT38), .Z(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n531), .A2(new_n544), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n520), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(G902), .B1(new_n711), .B2(KEYINPUT101), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n712), .B1(KEYINPUT101), .B2(new_n711), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(G472), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n539), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  AOI22_X1  g530(.A1(new_n653), .A2(new_n655), .B1(new_n662), .B2(G475), .ZN(new_n717));
  INV_X1    g531(.A(new_n489), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n609), .A2(new_n677), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n718), .A2(new_n719), .A3(new_n328), .ZN(new_n720));
  NOR4_X1   g534(.A1(new_n709), .A2(new_n716), .A3(new_n717), .A4(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n703), .A2(new_n706), .A3(new_n721), .ZN(new_n722));
  XOR2_X1   g536(.A(new_n722), .B(new_n237), .Z(G45));
  NOR2_X1   g537(.A1(new_n643), .A2(new_n693), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n685), .A2(new_n689), .A3(new_n691), .A4(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G146), .ZN(G48));
  OAI21_X1  g540(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(G469), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n326), .A3(new_n323), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n557), .A2(new_n615), .A3(new_n647), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(KEYINPUT41), .B(G113), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n731), .B(new_n732), .ZN(G15));
  NAND4_X1  g547(.A1(new_n557), .A2(new_n665), .A3(new_n615), .A4(new_n730), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G116), .ZN(G18));
  NOR4_X1   g549(.A1(new_n687), .A2(new_n449), .A3(new_n729), .A4(new_n497), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n736), .A2(new_n685), .A3(new_n691), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G119), .ZN(G21));
  NAND2_X1  g552(.A1(new_n382), .A2(new_n718), .ZN(new_n739));
  NOR4_X1   g553(.A1(new_n717), .A2(new_n739), .A3(new_n729), .A4(new_n495), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT103), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n532), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n544), .B1(new_n532), .B2(new_n741), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n500), .B(new_n320), .C1(new_n744), .C2(new_n525), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(new_n615), .A3(new_n623), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n746), .A2(KEYINPUT104), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(KEYINPUT104), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n740), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G122), .ZN(G24));
  NAND2_X1  g564(.A1(new_n745), .A2(new_n623), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n751), .A2(new_n719), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n383), .A2(new_n729), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n724), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G125), .ZN(G27));
  NAND2_X1  g569(.A1(new_n637), .A2(new_n641), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n653), .A2(new_n655), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n662), .A2(G475), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NOR4_X1   g573(.A1(new_n644), .A2(new_n645), .A3(new_n688), .A4(new_n329), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n302), .A2(KEYINPUT106), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n761), .A2(new_n316), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT107), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT106), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n313), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n762), .A2(new_n763), .A3(G469), .A4(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n765), .A2(G469), .A3(new_n316), .A4(new_n761), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(KEYINPUT107), .ZN(new_n768));
  NAND2_X1  g582(.A1(G469), .A2(G902), .ZN(new_n769));
  XOR2_X1   g583(.A(new_n769), .B(KEYINPUT105), .Z(new_n770));
  AND2_X1   g584(.A1(new_n323), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n766), .A2(new_n768), .A3(new_n771), .ZN(new_n772));
  AND4_X1   g586(.A1(new_n759), .A2(new_n694), .A3(new_n760), .A4(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT108), .B1(new_n684), .B2(new_n615), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT108), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n690), .A2(new_n618), .A3(new_n775), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n773), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(KEYINPUT42), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n772), .A2(new_n760), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n643), .A2(KEYINPUT42), .A3(new_n693), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n557), .A2(new_n615), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(new_n263), .ZN(G33));
  NAND4_X1  g597(.A1(new_n557), .A2(new_n615), .A3(new_n695), .A4(new_n779), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G134), .ZN(G36));
  NOR3_X1   g599(.A1(new_n644), .A2(new_n329), .A3(new_n645), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n449), .A2(new_n756), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(KEYINPUT43), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n624), .A2(new_n719), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT44), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n787), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n770), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n309), .A2(KEYINPUT45), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n795), .A2(new_n318), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n762), .A2(KEYINPUT45), .A3(new_n765), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n794), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(KEYINPUT46), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n323), .B1(new_n798), .B2(KEYINPUT46), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n326), .B(new_n699), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT109), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n798), .A2(KEYINPUT46), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n323), .A3(new_n799), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n806), .A2(KEYINPUT109), .A3(new_n326), .A4(new_n699), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n789), .A2(KEYINPUT44), .A3(new_n790), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n793), .A2(new_n804), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G137), .ZN(G39));
  INV_X1    g624(.A(KEYINPUT47), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n806), .B(new_n326), .C1(KEYINPUT110), .C2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n800), .A2(new_n801), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n811), .A2(KEYINPUT110), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n811), .A2(KEYINPUT110), .ZN(new_n815));
  OAI22_X1  g629(.A1(new_n813), .A2(new_n688), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n724), .A2(new_n618), .A3(new_n786), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n557), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n812), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  XOR2_X1   g633(.A(KEYINPUT111), .B(G140), .Z(new_n820));
  XNOR2_X1  g634(.A(new_n819), .B(new_n820), .ZN(G42));
  NAND2_X1  g635(.A1(new_n728), .A2(new_n323), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n708), .B1(KEYINPUT49), .B2(new_n822), .ZN(new_n823));
  OR2_X1    g637(.A1(new_n822), .A2(KEYINPUT49), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n615), .A2(new_n326), .A3(new_n328), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n825), .A2(new_n449), .A3(new_n756), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n823), .A2(new_n716), .A3(new_n824), .A4(new_n826), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n789), .B(new_n491), .C1(new_n748), .C2(new_n747), .ZN(new_n828));
  NOR4_X1   g642(.A1(new_n828), .A2(new_n328), .A3(new_n708), .A4(new_n729), .ZN(new_n829));
  NOR2_X1   g643(.A1(KEYINPUT118), .A2(KEYINPUT50), .ZN(new_n830));
  XOR2_X1   g644(.A(new_n829), .B(new_n830), .Z(new_n831));
  AND4_X1   g645(.A1(new_n491), .A2(new_n760), .A3(new_n323), .A4(new_n728), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n789), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n752), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n716), .A2(new_n615), .A3(new_n832), .ZN(new_n835));
  OR3_X1    g649(.A1(new_n835), .A2(new_n449), .A3(new_n642), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n831), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n828), .A2(new_n787), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n812), .A2(new_n816), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n822), .A2(new_n326), .ZN(new_n842));
  XOR2_X1   g656(.A(new_n842), .B(KEYINPUT117), .Z(new_n843));
  OAI21_X1  g657(.A(new_n839), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(KEYINPUT51), .B1(new_n838), .B2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n786), .A2(new_n758), .A3(new_n489), .A4(new_n694), .ZN(new_n846));
  NOR4_X1   g660(.A1(new_n327), .A2(new_n846), .A3(new_n658), .A4(new_n679), .ZN(new_n847));
  AOI22_X1  g661(.A1(new_n847), .A2(new_n557), .B1(new_n773), .B2(new_n752), .ZN(new_n848));
  AND4_X1   g662(.A1(new_n778), .A2(new_n848), .A3(new_n781), .A4(new_n784), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT113), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n660), .A2(new_n642), .A3(new_n449), .A4(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n717), .A2(new_n718), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n851), .B1(new_n646), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n850), .B1(new_n759), .B2(new_n660), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n625), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n681), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n557), .A2(KEYINPUT77), .A3(new_n615), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n685), .A2(new_n691), .A3(new_n615), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n617), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n856), .B1(new_n860), .B2(new_n499), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT112), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n685), .A2(new_n691), .A3(new_n615), .A4(new_n730), .ZN(new_n863));
  INV_X1    g677(.A(new_n647), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n737), .B(new_n749), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n863), .A2(new_n664), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n862), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n749), .A2(new_n737), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n868), .A2(KEYINPUT112), .A3(new_n731), .A4(new_n734), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n849), .A2(new_n861), .A3(new_n867), .A4(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n717), .A2(new_n739), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n693), .A2(KEYINPUT115), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n693), .A2(KEYINPUT115), .ZN(new_n873));
  AND4_X1   g687(.A1(new_n326), .A2(new_n719), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n715), .A2(new_n871), .A3(new_n772), .A4(new_n874), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n725), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n876), .A2(KEYINPUT52), .A3(new_n696), .A4(new_n754), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT52), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n725), .A2(new_n875), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n696), .A2(new_n754), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(KEYINPUT53), .B1(new_n870), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n880), .A2(KEYINPUT114), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n725), .A2(KEYINPUT52), .A3(new_n875), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT114), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n696), .A2(new_n886), .A3(new_n754), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n884), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT116), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n888), .A2(new_n889), .A3(new_n881), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n889), .B1(new_n888), .B2(new_n881), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n867), .A2(new_n869), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT53), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n893), .A2(new_n894), .A3(new_n861), .A4(new_n849), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n883), .B(KEYINPUT54), .C1(new_n892), .C2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n856), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n620), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n868), .A2(KEYINPUT53), .A3(new_n731), .A4(new_n734), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n778), .A2(new_n848), .A3(new_n781), .A4(new_n784), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n901), .B1(new_n890), .B2(new_n891), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n894), .B1(new_n870), .B2(new_n882), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT54), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n896), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n833), .B1(new_n774), .B2(new_n776), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n907), .B(KEYINPUT48), .Z(new_n908));
  NOR2_X1   g722(.A1(new_n490), .A2(G953), .ZN(new_n909));
  INV_X1    g723(.A(new_n753), .ZN(new_n910));
  OAI221_X1 g724(.A(new_n909), .B1(new_n643), .B2(new_n835), .C1(new_n828), .C2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n839), .B1(new_n841), .B2(new_n842), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(KEYINPUT51), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n912), .B1(new_n837), .B2(new_n914), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n845), .A2(new_n906), .A3(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(G952), .A2(G953), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n827), .B1(new_n916), .B2(new_n917), .ZN(G75));
  NOR2_X1   g732(.A1(new_n190), .A2(G952), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n320), .B1(new_n902), .B2(new_n903), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT56), .B1(new_n921), .B2(new_n378), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n355), .A2(new_n366), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT119), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n364), .B(KEYINPUT55), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n924), .B(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n920), .B1(new_n922), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n927), .B1(new_n922), .B2(new_n926), .ZN(G51));
  AND3_X1   g742(.A1(new_n921), .A2(new_n797), .A3(new_n796), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n321), .A2(new_n322), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n902), .A2(new_n903), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(KEYINPUT54), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n905), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n770), .B(KEYINPUT57), .Z(new_n934));
  AOI21_X1  g748(.A(new_n930), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n929), .B1(new_n935), .B2(KEYINPUT120), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT120), .ZN(new_n937));
  INV_X1    g751(.A(new_n934), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n938), .B1(new_n932), .B2(new_n905), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n937), .B1(new_n939), .B2(new_n930), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n919), .B1(new_n936), .B2(new_n940), .ZN(G54));
  AND2_X1   g755(.A1(KEYINPUT58), .A2(G475), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n921), .A2(new_n440), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n440), .B1(new_n921), .B2(new_n942), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n943), .A2(new_n944), .A3(new_n919), .ZN(G60));
  NAND2_X1  g759(.A1(G478), .A2(G902), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT59), .Z(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n906), .A2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT122), .ZN(new_n950));
  INV_X1    g764(.A(new_n635), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n947), .B1(new_n896), .B2(new_n905), .ZN(new_n953));
  OAI21_X1  g767(.A(KEYINPUT122), .B1(new_n953), .B2(new_n635), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n951), .A2(new_n947), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n904), .B1(new_n902), .B2(new_n903), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT121), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI211_X1 g775(.A(KEYINPUT121), .B(new_n956), .C1(new_n957), .C2(new_n958), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n919), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n955), .A2(new_n963), .ZN(G63));
  NAND2_X1  g778(.A1(G217), .A2(G902), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT60), .Z(new_n966));
  NAND3_X1  g780(.A1(new_n931), .A2(new_n674), .A3(new_n966), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n931), .A2(new_n966), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n920), .B(new_n967), .C1(new_n968), .C2(new_n612), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT61), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(G66));
  OAI21_X1  g785(.A(G953), .B1(new_n494), .B2(new_n361), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n893), .A2(new_n861), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n190), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n972), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n924), .B1(G898), .B2(new_n190), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT123), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n976), .B(new_n978), .ZN(G69));
  NAND3_X1  g793(.A1(new_n778), .A2(new_n781), .A3(new_n784), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n804), .A2(new_n807), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n774), .A2(new_n776), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n982), .A2(new_n717), .A3(new_n739), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n980), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  AND3_X1   g798(.A1(new_n884), .A2(new_n725), .A3(new_n887), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n984), .A2(new_n809), .A3(new_n819), .A4(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(new_n190), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n508), .A2(new_n509), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(new_n434), .ZN(new_n989));
  INV_X1    g803(.A(G227), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n989), .B1(new_n990), .B2(new_n975), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n987), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n692), .B1(new_n989), .B2(new_n990), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n722), .A2(new_n725), .A3(new_n884), .A4(new_n887), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT62), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n985), .A2(KEYINPUT62), .A3(new_n722), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n809), .A2(new_n819), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n852), .A2(new_n643), .ZN(new_n1000));
  AND4_X1   g814(.A1(new_n698), .A2(new_n1000), .A3(new_n699), .A4(new_n786), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n999), .B1(new_n860), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n998), .A2(new_n1002), .A3(KEYINPUT124), .ZN(new_n1003));
  INV_X1    g817(.A(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(KEYINPUT124), .B1(new_n998), .B2(new_n1002), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n989), .A2(new_n190), .ZN(new_n1007));
  OAI221_X1 g821(.A(new_n992), .B1(new_n190), .B2(new_n993), .C1(new_n1006), .C2(new_n1007), .ZN(G72));
  INV_X1    g822(.A(KEYINPUT127), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n522), .A2(new_n510), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(new_n519), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1005), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1012), .A2(new_n974), .A3(new_n1003), .ZN(new_n1013));
  XNOR2_X1  g827(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n500), .A2(new_n320), .ZN(new_n1015));
  XOR2_X1   g829(.A(new_n1014), .B(new_n1015), .Z(new_n1016));
  INV_X1    g830(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1011), .B1(new_n1013), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1017), .B1(new_n986), .B2(new_n973), .ZN(new_n1019));
  XOR2_X1   g833(.A(new_n545), .B(KEYINPUT126), .Z(new_n1020));
  AOI21_X1  g834(.A(new_n919), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  AND3_X1   g835(.A1(new_n1011), .A2(new_n545), .A3(new_n1017), .ZN(new_n1022));
  OAI211_X1 g836(.A(new_n883), .B(new_n1022), .C1(new_n892), .C2(new_n895), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1009), .B1(new_n1018), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(new_n1024), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1016), .B1(new_n1006), .B2(new_n974), .ZN(new_n1027));
  OAI211_X1 g841(.A(new_n1026), .B(KEYINPUT127), .C1(new_n1027), .C2(new_n1011), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1025), .A2(new_n1028), .ZN(G57));
endmodule


