//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 0 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 1 0 0 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:52 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0004(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n205));
  INV_X1    g0005(.A(G116), .ZN(new_n206));
  INV_X1    g0006(.A(G270), .ZN(new_n207));
  XNOR2_X1  g0007(.A(KEYINPUT65), .B(G77), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  XOR2_X1   g0009(.A(KEYINPUT66), .B(G244), .Z(new_n210));
  OAI221_X1 g0010(.A(new_n205), .B1(new_n206), .B2(new_n207), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT67), .ZN(new_n212));
  OR2_X1    g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G97), .A2(G257), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n211), .A2(new_n212), .ZN(new_n215));
  INV_X1    g0015(.A(G58), .ZN(new_n216));
  INV_X1    g0016(.A(G232), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  OAI22_X1  g0019(.A1(new_n216), .A2(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n220), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND4_X1  g0021(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G20), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT1), .Z(new_n225));
  OR2_X1    g0025(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n226), .A2(G50), .A3(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n223), .A2(G13), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  NOR2_X1   g0034(.A1(G257), .A2(G264), .ZN(new_n235));
  NOR3_X1   g0035(.A1(new_n234), .A2(new_n219), .A3(new_n235), .ZN(new_n236));
  AOI22_X1  g0036(.A1(new_n229), .A2(new_n232), .B1(new_n236), .B2(KEYINPUT0), .ZN(new_n237));
  OAI211_X1 g0037(.A(new_n225), .B(new_n237), .C1(KEYINPUT0), .C2(new_n236), .ZN(new_n238));
  INV_X1    g0038(.A(new_n238), .ZN(G361));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n217), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT2), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n242), .B(G226), .Z(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G264), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(new_n207), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G358));
  XNOR2_X1  g0047(.A(G50), .B(G68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G87), .B(G97), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(G107), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(new_n206), .ZN(new_n253));
  XOR2_X1   g0053(.A(new_n250), .B(new_n253), .Z(G351));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT3), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n256), .A2(new_n258), .A3(G223), .A4(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT76), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT3), .B(G33), .ZN(new_n263));
  NAND4_X1  g0063(.A1(new_n263), .A2(KEYINPUT76), .A3(G223), .A4(new_n259), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(G226), .A3(G1698), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G87), .ZN(new_n266));
  NAND4_X1  g0066(.A1(new_n262), .A2(new_n264), .A3(new_n265), .A4(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n230), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G1), .ZN(new_n273));
  INV_X1    g0073(.A(G41), .ZN(new_n274));
  INV_X1    g0074(.A(G45), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n273), .A2(new_n276), .B1(new_n268), .B2(new_n269), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G232), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n276), .A2(new_n273), .A3(G274), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n272), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G169), .ZN(new_n281));
  INV_X1    g0081(.A(G179), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n281), .B1(new_n282), .B2(new_n280), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT16), .ZN(new_n284));
  INV_X1    g0084(.A(G68), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT75), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n286), .B1(new_n255), .B2(KEYINPUT3), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n257), .A2(KEYINPUT75), .A3(G33), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n287), .A2(new_n256), .A3(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n289), .A2(KEYINPUT7), .A3(new_n231), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT7), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n291), .B1(new_n263), .B2(G20), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n285), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT74), .ZN(new_n294));
  NOR2_X1   g0094(.A1(G20), .A2(G33), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G159), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n294), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n295), .A2(KEYINPUT74), .A3(G159), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n216), .A2(new_n285), .ZN(new_n301));
  OAI21_X1  g0101(.A(G20), .B1(new_n301), .B2(new_n201), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n284), .B1(new_n293), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n256), .A2(new_n258), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n305), .A2(KEYINPUT7), .A3(new_n231), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n292), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G68), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n300), .A2(new_n302), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n308), .A2(new_n309), .A3(KEYINPUT16), .ZN(new_n310));
  NAND3_X1  g0110(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n230), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n304), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  XNOR2_X1  g0113(.A(KEYINPUT8), .B(G58), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT68), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT68), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n316), .A2(new_n216), .A3(KEYINPUT8), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n273), .A2(G13), .A3(G20), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n312), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(G1), .B2(new_n231), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n321), .B1(new_n318), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n313), .A2(new_n325), .ZN(new_n326));
  AND3_X1   g0126(.A1(new_n283), .A2(KEYINPUT18), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(KEYINPUT18), .B1(new_n283), .B2(new_n326), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n280), .A2(G200), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n272), .A2(G190), .A3(new_n278), .A4(new_n279), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n330), .A2(new_n313), .A3(new_n325), .A4(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT17), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n285), .B1(new_n292), .B2(new_n306), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n334), .A2(new_n303), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n322), .B1(new_n335), .B2(KEYINPUT16), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n324), .B1(new_n336), .B2(new_n304), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT17), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n337), .A2(new_n338), .A3(new_n330), .A4(new_n331), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n333), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT77), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n333), .A2(new_n339), .A3(KEYINPUT77), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n329), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n256), .A2(new_n258), .A3(G232), .A4(G1698), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT70), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT70), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n263), .A2(new_n347), .A3(G232), .A4(G1698), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G33), .A2(G97), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n263), .A2(G226), .A3(new_n259), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n346), .A2(new_n348), .A3(new_n349), .A4(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n271), .ZN(new_n352));
  OR2_X1    g0152(.A1(new_n277), .A2(KEYINPUT71), .ZN(new_n353));
  INV_X1    g0153(.A(G238), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n354), .B1(new_n277), .B2(KEYINPUT71), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n352), .A2(new_n279), .A3(new_n356), .ZN(new_n357));
  XOR2_X1   g0157(.A(KEYINPUT72), .B(KEYINPUT13), .Z(new_n358));
  NOR2_X1   g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n358), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n351), .A2(new_n271), .B1(new_n353), .B2(new_n355), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n360), .B1(new_n361), .B2(new_n279), .ZN(new_n362));
  OAI21_X1  g0162(.A(G169), .B1(new_n359), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT14), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n361), .A2(new_n279), .A3(new_n360), .ZN(new_n365));
  INV_X1    g0165(.A(new_n357), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT13), .ZN(new_n367));
  OAI211_X1 g0167(.A(G179), .B(new_n365), .C1(new_n366), .C2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n357), .A2(new_n358), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n365), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT14), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(new_n371), .A3(G169), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n364), .A2(new_n368), .A3(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n255), .A2(G20), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n374), .A2(G77), .B1(new_n295), .B2(G50), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(new_n231), .B2(G68), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n376), .A2(KEYINPUT11), .A3(new_n312), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n285), .B2(new_n323), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n319), .A2(G68), .ZN(new_n379));
  XNOR2_X1  g0179(.A(new_n379), .B(KEYINPUT12), .ZN(new_n380));
  AOI21_X1  g0180(.A(KEYINPUT11), .B1(new_n376), .B2(new_n312), .ZN(new_n381));
  NOR3_X1   g0181(.A1(new_n378), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n373), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n344), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n319), .A2(G50), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n315), .A2(new_n317), .A3(new_n374), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n295), .A2(G150), .ZN(new_n388));
  OAI21_X1  g0188(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n386), .B1(new_n390), .B2(new_n312), .ZN(new_n391));
  INV_X1    g0191(.A(G50), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n323), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n259), .A2(G222), .ZN(new_n396));
  NAND2_X1  g0196(.A1(G223), .A2(G1698), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n263), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n398), .B(new_n271), .C1(new_n208), .C2(new_n263), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n277), .A2(G226), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(new_n279), .A3(new_n400), .ZN(new_n401));
  OR2_X1    g0201(.A1(new_n401), .A2(G179), .ZN(new_n402));
  INV_X1    g0202(.A(G169), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  AND3_X1   g0204(.A1(new_n395), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G238), .A2(G1698), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n263), .B(new_n406), .C1(new_n217), .C2(G1698), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n407), .B(new_n271), .C1(G107), .C2(new_n263), .ZN(new_n408));
  INV_X1    g0208(.A(new_n277), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n408), .B(new_n279), .C1(new_n210), .C2(new_n409), .ZN(new_n410));
  OR2_X1    g0210(.A1(new_n410), .A2(G179), .ZN(new_n411));
  OAI22_X1  g0211(.A1(new_n209), .A2(new_n231), .B1(new_n314), .B2(new_n296), .ZN(new_n412));
  XNOR2_X1  g0212(.A(KEYINPUT15), .B(G87), .ZN(new_n413));
  NOR3_X1   g0213(.A1(new_n413), .A2(G20), .A3(new_n255), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n312), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(G77), .ZN(new_n416));
  OAI221_X1 g0216(.A(new_n415), .B1(new_n416), .B2(new_n323), .C1(new_n208), .C2(new_n319), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n410), .A2(new_n403), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n411), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT9), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n395), .A2(new_n420), .ZN(new_n421));
  AOI211_X1 g0221(.A(new_n386), .B(new_n393), .C1(new_n390), .C2(new_n312), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT9), .ZN(new_n423));
  INV_X1    g0223(.A(G190), .ZN(new_n424));
  OR2_X1    g0224(.A1(new_n401), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n401), .A2(G200), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n421), .A2(new_n423), .A3(new_n425), .A4(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT10), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n422), .A2(KEYINPUT9), .B1(G200), .B2(new_n401), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT10), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n429), .A2(new_n430), .A3(new_n425), .A4(new_n421), .ZN(new_n431));
  AOI211_X1 g0231(.A(new_n405), .B(new_n419), .C1(new_n428), .C2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n370), .A2(G200), .ZN(new_n433));
  OAI211_X1 g0233(.A(G190), .B(new_n365), .C1(new_n366), .C2(new_n367), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n433), .A2(new_n382), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT73), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT73), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n433), .A2(new_n437), .A3(new_n434), .A4(new_n382), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n417), .A2(KEYINPUT69), .B1(G200), .B2(new_n410), .ZN(new_n439));
  OAI221_X1 g0239(.A(new_n439), .B1(KEYINPUT69), .B2(new_n417), .C1(new_n424), .C2(new_n410), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n432), .A2(new_n436), .A3(new_n438), .A4(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n385), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(G97), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n320), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n273), .A2(G33), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n322), .A2(new_n319), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(G107), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n448), .B1(new_n290), .B2(new_n292), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n296), .A2(new_n416), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT6), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n444), .A2(new_n448), .ZN(new_n452));
  NOR2_X1   g0252(.A1(G97), .A2(G107), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n448), .A2(KEYINPUT6), .A3(G97), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n231), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n449), .A2(new_n450), .A3(new_n456), .ZN(new_n457));
  OAI221_X1 g0257(.A(new_n445), .B1(new_n444), .B2(new_n447), .C1(new_n457), .C2(new_n322), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n256), .A2(new_n258), .A3(G250), .A4(G1698), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT78), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n263), .A2(KEYINPUT78), .A3(G250), .A4(G1698), .ZN(new_n462));
  NAND2_X1  g0262(.A1(G33), .A2(G283), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n256), .A2(new_n258), .A3(G244), .A4(new_n259), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT4), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n263), .A2(KEYINPUT4), .A3(G244), .A4(new_n259), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n271), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n273), .A2(G45), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT5), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n274), .ZN(new_n473));
  NAND2_X1  g0273(.A1(KEYINPUT5), .A2(G41), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G274), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n473), .A2(new_n474), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n275), .A2(G1), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n478), .A2(new_n479), .B1(new_n268), .B2(new_n269), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n477), .B1(G257), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n470), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(new_n424), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n458), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT79), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n470), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g0286(.A(KEYINPUT79), .B(new_n271), .C1(new_n464), .C2(new_n469), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n486), .A2(new_n481), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G200), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT80), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n488), .A2(KEYINPUT80), .A3(G200), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n484), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n486), .A2(new_n282), .A3(new_n481), .A4(new_n487), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n482), .A2(new_n403), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n458), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n257), .A2(G33), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n499));
  OAI21_X1  g0299(.A(G303), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n256), .A2(new_n258), .A3(G257), .A4(new_n259), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n256), .A2(new_n258), .A3(G264), .A4(G1698), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  AND2_X1   g0303(.A1(new_n503), .A2(new_n271), .ZN(new_n504));
  INV_X1    g0304(.A(new_n474), .ZN(new_n505));
  NOR2_X1   g0305(.A1(KEYINPUT5), .A2(G41), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n479), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n270), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n476), .B1(new_n508), .B2(new_n207), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n504), .A2(new_n509), .A3(new_n282), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n320), .A2(new_n206), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n322), .A2(G116), .A3(new_n319), .A4(new_n446), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n311), .A2(new_n230), .B1(G20), .B2(new_n206), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n463), .B(new_n231), .C1(G33), .C2(new_n444), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n513), .A2(KEYINPUT20), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(KEYINPUT20), .B1(new_n513), .B2(new_n514), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n511), .B(new_n512), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n510), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(G169), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT82), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n520), .B1(new_n504), .B2(new_n509), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n480), .A2(G270), .B1(G274), .B2(new_n475), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n503), .A2(new_n271), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n522), .A2(new_n523), .A3(KEYINPUT82), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n519), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n518), .B1(new_n525), .B2(KEYINPUT21), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n513), .A2(new_n514), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT20), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n513), .A2(KEYINPUT20), .A3(new_n514), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n529), .A2(new_n530), .B1(new_n206), .B2(new_n320), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n403), .B1(new_n531), .B2(new_n512), .ZN(new_n532));
  AND3_X1   g0332(.A1(new_n522), .A2(new_n523), .A3(KEYINPUT82), .ZN(new_n533));
  AOI21_X1  g0333(.A(KEYINPUT82), .B1(new_n522), .B2(new_n523), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n532), .B(KEYINPUT21), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT83), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n521), .A2(new_n524), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n538), .A2(KEYINPUT83), .A3(KEYINPUT21), .A4(new_n532), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n526), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(G200), .B1(new_n533), .B2(new_n534), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n521), .A2(G190), .A3(new_n524), .ZN(new_n542));
  INV_X1    g0342(.A(new_n517), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT84), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n541), .A2(new_n542), .A3(KEYINPUT84), .A4(new_n543), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n320), .A2(new_n448), .ZN(new_n549));
  OAI22_X1  g0349(.A1(new_n447), .A2(new_n448), .B1(new_n549), .B2(KEYINPUT25), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n256), .A2(new_n258), .A3(new_n231), .A4(G87), .ZN(new_n551));
  NAND2_X1  g0351(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OR2_X1    g0353(.A1(KEYINPUT86), .A2(KEYINPUT23), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n448), .A2(G20), .ZN(new_n555));
  NAND2_X1  g0355(.A1(KEYINPUT86), .A2(KEYINPUT23), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n448), .A2(KEYINPUT86), .A3(KEYINPUT23), .A4(G20), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(KEYINPUT85), .A2(KEYINPUT22), .A3(G87), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n263), .A2(new_n561), .B1(G33), .B2(G116), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n553), .B(new_n559), .C1(new_n562), .C2(G20), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(KEYINPUT24), .ZN(new_n564));
  NAND2_X1  g0364(.A1(G33), .A2(G116), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n305), .B2(new_n560), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n231), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT24), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n567), .A2(new_n568), .A3(new_n553), .A4(new_n559), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n550), .B1(new_n570), .B2(new_n312), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n549), .A2(KEYINPUT25), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n256), .A2(new_n258), .A3(G257), .A4(G1698), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(KEYINPUT87), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT87), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n263), .A2(new_n576), .A3(G257), .A4(G1698), .ZN(new_n577));
  NAND2_X1  g0377(.A1(G33), .A2(G294), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n263), .A2(G250), .A3(new_n259), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n575), .A2(new_n577), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n580), .A2(new_n271), .B1(G264), .B2(new_n480), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n581), .A2(G190), .A3(new_n476), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n580), .A2(new_n271), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n480), .A2(G264), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n583), .A2(new_n476), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(G200), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n571), .A2(new_n573), .A3(new_n582), .A4(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT19), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n231), .B1(new_n349), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n453), .A2(new_n218), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n256), .A2(new_n258), .A3(new_n231), .A4(G68), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n588), .B1(new_n349), .B2(G20), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n312), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n413), .A2(new_n320), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n322), .A2(G87), .A3(new_n319), .A4(new_n446), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n256), .A2(new_n258), .A3(G244), .A4(G1698), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n256), .A2(new_n258), .A3(G238), .A4(new_n259), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n599), .A2(new_n600), .A3(new_n565), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n271), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n479), .A2(G274), .ZN(new_n603));
  INV_X1    g0403(.A(new_n269), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n471), .B(G250), .C1(new_n604), .C2(new_n230), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n602), .A2(G190), .A3(new_n603), .A4(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(G200), .ZN(new_n607));
  INV_X1    g0407(.A(new_n603), .ZN(new_n608));
  INV_X1    g0408(.A(new_n605), .ZN(new_n609));
  AOI211_X1 g0409(.A(new_n608), .B(new_n609), .C1(new_n601), .C2(new_n271), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n598), .B(new_n606), .C1(new_n607), .C2(new_n610), .ZN(new_n611));
  XNOR2_X1  g0411(.A(new_n413), .B(KEYINPUT81), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n595), .B(new_n596), .C1(new_n447), .C2(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n602), .A2(new_n282), .A3(new_n603), .A4(new_n605), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n613), .B(new_n614), .C1(new_n610), .C2(G169), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n587), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n570), .A2(new_n312), .ZN(new_n618));
  INV_X1    g0418(.A(new_n550), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n618), .A2(new_n573), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n585), .A2(new_n403), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n581), .A2(new_n282), .A3(new_n476), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n540), .A2(new_n548), .A3(new_n617), .A4(new_n623), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n443), .A2(new_n497), .A3(new_n624), .ZN(G372));
  OR2_X1    g0425(.A1(new_n327), .A2(new_n328), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n342), .A2(new_n343), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n373), .A2(new_n383), .B1(new_n419), .B2(new_n435), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT90), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n435), .A2(new_n419), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n384), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n626), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n428), .A2(new_n431), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n405), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n537), .A2(new_n539), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n538), .A2(new_n532), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT21), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n637), .A2(new_n638), .B1(new_n510), .B2(new_n517), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n636), .A2(new_n623), .A3(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT88), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n641), .B1(new_n610), .B2(new_n607), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n602), .A2(new_n603), .A3(new_n605), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n643), .A2(KEYINPUT88), .A3(G200), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n642), .A2(new_n606), .A3(new_n644), .A4(new_n598), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n587), .A2(new_n615), .A3(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n640), .A2(new_n646), .A3(new_n493), .A4(new_n496), .ZN(new_n647));
  XOR2_X1   g0447(.A(new_n615), .B(KEYINPUT89), .Z(new_n648));
  NAND2_X1  g0448(.A1(new_n611), .A2(new_n615), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT26), .B1(new_n496), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n645), .A2(new_n615), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n458), .A2(new_n495), .A3(new_n494), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT26), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n647), .A2(new_n648), .A3(new_n650), .A4(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n635), .B1(new_n657), .B2(new_n443), .ZN(G369));
  INV_X1    g0458(.A(G13), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(G20), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n273), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(G213), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(G343), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(new_n543), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n540), .A2(new_n548), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n670), .B1(new_n540), .B2(new_n669), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n671), .A2(G330), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n623), .A2(new_n666), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n620), .A2(new_n666), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n587), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n673), .B1(new_n675), .B2(new_n623), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n636), .A2(new_n639), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n667), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT91), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n679), .B(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n673), .B1(new_n681), .B2(new_n676), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n677), .A2(new_n682), .ZN(G399));
  NOR2_X1   g0483(.A1(new_n590), .A2(G116), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n234), .A2(G41), .ZN(new_n686));
  NOR3_X1   g0486(.A1(new_n685), .A2(new_n686), .A3(new_n273), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n687), .A2(KEYINPUT92), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n229), .A2(new_n686), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n687), .A2(KEYINPUT92), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n691), .B(KEYINPUT28), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT29), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n656), .A2(new_n693), .A3(new_n667), .ZN(new_n694));
  OAI21_X1  g0494(.A(KEYINPUT26), .B1(new_n651), .B2(new_n496), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n653), .A2(new_n654), .A3(new_n616), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n647), .A2(new_n648), .A3(new_n695), .A4(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n693), .B1(new_n697), .B2(new_n667), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(G330), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n610), .A2(G179), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n488), .A2(new_n538), .A3(new_n585), .A4(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n610), .A2(new_n470), .A3(new_n481), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n705), .A2(KEYINPUT30), .A3(new_n510), .A4(new_n581), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT30), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n510), .A2(new_n581), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n707), .B1(new_n708), .B2(new_n704), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n703), .A2(new_n706), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(KEYINPUT93), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT93), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n703), .A2(new_n706), .A3(new_n709), .A4(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n711), .A2(new_n666), .A3(new_n713), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n624), .A2(new_n497), .A3(new_n666), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT31), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n710), .A2(KEYINPUT31), .A3(new_n666), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n701), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n700), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n692), .B1(new_n720), .B2(G1), .ZN(G364));
  AOI21_X1  g0521(.A(new_n273), .B1(new_n660), .B2(G45), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n686), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT94), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n672), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(G330), .B2(new_n671), .ZN(new_n727));
  INV_X1    g0527(.A(new_n725), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n250), .A2(G45), .ZN(new_n729));
  AOI22_X1  g0529(.A1(new_n729), .A2(KEYINPUT95), .B1(new_n275), .B2(new_n229), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n234), .A2(new_n263), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n730), .B(new_n731), .C1(KEYINPUT95), .C2(new_n729), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n263), .A2(G355), .A3(new_n233), .ZN(new_n733));
  OAI211_X1 g0533(.A(new_n732), .B(new_n733), .C1(G116), .C2(new_n233), .ZN(new_n734));
  NOR2_X1   g0534(.A1(G13), .A2(G33), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G20), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n230), .B1(G20), .B2(new_n403), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n728), .B1(new_n734), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n737), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n231), .A2(new_n424), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n282), .A2(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR4_X1   g0545(.A1(new_n231), .A2(new_n282), .A3(new_n424), .A4(new_n607), .ZN(new_n746));
  AOI22_X1  g0546(.A1(new_n745), .A2(G322), .B1(new_n746), .B2(G326), .ZN(new_n747));
  INV_X1    g0547(.A(G294), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G179), .A2(G200), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n231), .B1(new_n749), .B2(G190), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n747), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n231), .A2(G190), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(new_n749), .ZN(new_n753));
  INV_X1    g0553(.A(G329), .ZN(new_n754));
  XOR2_X1   g0554(.A(KEYINPUT33), .B(G317), .Z(new_n755));
  NAND3_X1  g0555(.A1(new_n752), .A2(G179), .A3(G200), .ZN(new_n756));
  OAI221_X1 g0556(.A(new_n305), .B1(new_n753), .B2(new_n754), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n282), .A2(G200), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT97), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n742), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n757), .B1(new_n761), .B2(G303), .ZN(new_n762));
  INV_X1    g0562(.A(G283), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n759), .A2(new_n752), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n752), .A2(new_n743), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n751), .B(new_n765), .C1(G311), .C2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n750), .A2(new_n444), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n769), .B1(G50), .B2(new_n746), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n770), .B1(new_n216), .B2(new_n744), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n761), .A2(G87), .ZN(new_n772));
  INV_X1    g0572(.A(new_n756), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n305), .B1(new_n773), .B2(G68), .ZN(new_n774));
  OAI211_X1 g0574(.A(new_n772), .B(new_n774), .C1(new_n209), .C2(new_n766), .ZN(new_n775));
  INV_X1    g0575(.A(new_n764), .ZN(new_n776));
  AOI211_X1 g0576(.A(new_n771), .B(new_n775), .C1(G107), .C2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n753), .A2(new_n297), .ZN(new_n778));
  XOR2_X1   g0578(.A(KEYINPUT96), .B(KEYINPUT32), .Z(new_n779));
  XNOR2_X1  g0579(.A(new_n778), .B(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n768), .B1(new_n777), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT98), .ZN(new_n782));
  INV_X1    g0582(.A(new_n738), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n740), .B1(new_n671), .B2(new_n741), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n727), .A2(new_n784), .ZN(G396));
  NAND2_X1  g0585(.A1(new_n656), .A2(new_n667), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n417), .A2(new_n666), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n419), .B1(new_n440), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n788), .B1(new_n419), .B2(new_n667), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n786), .B(new_n789), .Z(new_n790));
  INV_X1    g0590(.A(new_n719), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n728), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT101), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n790), .A2(new_n791), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n218), .A2(new_n764), .B1(new_n760), .B2(new_n448), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n769), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n756), .A2(new_n763), .B1(new_n766), .B2(new_n206), .ZN(new_n798));
  XOR2_X1   g0598(.A(new_n798), .B(KEYINPUT99), .Z(new_n799));
  INV_X1    g0599(.A(new_n746), .ZN(new_n800));
  INV_X1    g0600(.A(G303), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n800), .A2(new_n801), .B1(new_n748), .B2(new_n744), .ZN(new_n802));
  INV_X1    g0602(.A(new_n753), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n802), .B1(G311), .B2(new_n803), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n797), .A2(new_n799), .A3(new_n305), .A4(new_n804), .ZN(new_n805));
  AOI22_X1  g0605(.A1(G150), .A2(new_n773), .B1(new_n746), .B2(G137), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT100), .ZN(new_n807));
  INV_X1    g0607(.A(G143), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n807), .B1(new_n808), .B2(new_n744), .C1(new_n297), .C2(new_n766), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT34), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n776), .A2(G68), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n810), .B(new_n811), .C1(new_n216), .C2(new_n750), .ZN(new_n812));
  INV_X1    g0612(.A(G132), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n263), .B1(new_n813), .B2(new_n753), .C1(new_n760), .C2(new_n392), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n805), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n728), .B1(new_n815), .B2(new_n738), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n783), .A2(new_n736), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n816), .B1(G77), .B2(new_n817), .C1(new_n736), .C2(new_n789), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n795), .A2(new_n818), .ZN(G384));
  NOR2_X1   g0619(.A1(new_n714), .A2(new_n716), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n717), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n789), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n382), .A2(new_n667), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n384), .A2(new_n435), .A3(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n373), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n828), .A2(new_n436), .A3(new_n438), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(new_n824), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(KEYINPUT104), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT104), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n829), .A2(new_n832), .A3(new_n824), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n827), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n823), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n336), .B1(KEYINPUT16), .B2(new_n335), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n325), .ZN(new_n837));
  INV_X1    g0637(.A(new_n664), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n837), .B1(new_n283), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n839), .A2(new_n332), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT37), .ZN(new_n841));
  XNOR2_X1  g0641(.A(KEYINPUT105), .B(KEYINPUT37), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n283), .A2(new_n326), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n326), .A2(new_n838), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n843), .A2(new_n332), .A3(new_n844), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n840), .A2(new_n841), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n837), .A2(new_n838), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n846), .B1(new_n344), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT38), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n846), .B(KEYINPUT38), .C1(new_n344), .C2(new_n847), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n853), .A2(KEYINPUT40), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n835), .A2(new_n854), .ZN(new_n855));
  AND3_X1   g0655(.A1(new_n829), .A2(new_n832), .A3(new_n824), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n832), .B1(new_n829), .B2(new_n824), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n826), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n844), .B1(new_n626), .B2(new_n340), .ZN(new_n859));
  INV_X1    g0659(.A(new_n842), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n845), .B(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n849), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n851), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n822), .A2(new_n858), .A3(new_n789), .A4(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(KEYINPUT40), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n855), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n822), .A2(new_n442), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n866), .B(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(G330), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n863), .A2(KEYINPUT39), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT39), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(new_n850), .B2(new_n851), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n384), .A2(new_n666), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n656), .A2(new_n789), .A3(new_n667), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n419), .A2(new_n667), .ZN(new_n878));
  XOR2_X1   g0678(.A(new_n878), .B(KEYINPUT103), .Z(new_n879));
  NAND2_X1  g0679(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n858), .A2(new_n880), .ZN(new_n881));
  OAI22_X1  g0681(.A1(new_n853), .A2(new_n881), .B1(new_n626), .B2(new_n838), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n876), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n869), .B(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n442), .B1(new_n694), .B2(new_n698), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n635), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n886), .B(KEYINPUT106), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n884), .B(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n273), .B2(new_n660), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n454), .A2(new_n455), .ZN(new_n890));
  OAI211_X1 g0690(.A(G116), .B(new_n232), .C1(new_n890), .C2(KEYINPUT35), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n891), .B(KEYINPUT102), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(KEYINPUT35), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(KEYINPUT36), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n208), .B1(new_n216), .B2(new_n285), .ZN(new_n896));
  OAI22_X1  g0696(.A1(new_n228), .A2(new_n896), .B1(G50), .B2(new_n285), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n897), .A2(G1), .A3(new_n659), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n889), .A2(new_n895), .A3(new_n898), .ZN(G367));
  NOR2_X1   g0699(.A1(new_n760), .A2(new_n206), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT46), .ZN(new_n901));
  OAI221_X1 g0701(.A(new_n305), .B1(new_n766), .B2(new_n763), .C1(new_n748), .C2(new_n756), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n902), .B1(new_n776), .B2(G97), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n745), .A2(G303), .B1(new_n746), .B2(G311), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n903), .B(new_n904), .C1(new_n448), .C2(new_n750), .ZN(new_n905));
  XNOR2_X1  g0705(.A(KEYINPUT109), .B(G317), .ZN(new_n906));
  AOI211_X1 g0706(.A(new_n901), .B(new_n905), .C1(new_n803), .C2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n750), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n745), .A2(G150), .B1(new_n908), .B2(G68), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n808), .B2(new_n800), .ZN(new_n910));
  INV_X1    g0710(.A(G137), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n263), .B1(new_n753), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(G50), .B2(new_n767), .ZN(new_n913));
  OAI221_X1 g0713(.A(new_n913), .B1(new_n216), .B2(new_n760), .C1(new_n209), .C2(new_n764), .ZN(new_n914));
  AOI211_X1 g0714(.A(new_n910), .B(new_n914), .C1(G159), .C2(new_n773), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n907), .A2(new_n915), .ZN(new_n916));
  XOR2_X1   g0716(.A(new_n916), .B(KEYINPUT47), .Z(new_n917));
  AOI21_X1  g0717(.A(new_n728), .B1(new_n917), .B2(new_n738), .ZN(new_n918));
  INV_X1    g0718(.A(new_n731), .ZN(new_n919));
  OAI221_X1 g0719(.A(new_n739), .B1(new_n233), .B2(new_n413), .C1(new_n246), .C2(new_n919), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n667), .A2(new_n598), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n652), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n648), .B2(new_n921), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n918), .B(new_n920), .C1(new_n741), .C2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT108), .ZN(new_n925));
  INV_X1    g0725(.A(new_n682), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n488), .A2(KEYINPUT80), .A3(G200), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT80), .B1(new_n488), .B2(G200), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n653), .B1(new_n929), .B2(new_n484), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n458), .A2(new_n666), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n653), .A2(new_n666), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT44), .B1(new_n926), .B2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT44), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n682), .A2(new_n937), .A3(new_n934), .ZN(new_n938));
  AND3_X1   g0738(.A1(new_n682), .A2(KEYINPUT45), .A3(new_n934), .ZN(new_n939));
  AOI21_X1  g0739(.A(KEYINPUT45), .B1(new_n682), .B2(new_n934), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n936), .A2(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n677), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n677), .B1(new_n939), .B2(new_n940), .C1(new_n936), .C2(new_n938), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n681), .A2(new_n676), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n679), .A2(new_n680), .ZN(new_n946));
  AOI21_X1  g0746(.A(KEYINPUT91), .B1(new_n678), .B2(new_n667), .ZN(new_n947));
  OR3_X1    g0747(.A1(new_n946), .A2(new_n676), .A3(new_n947), .ZN(new_n948));
  AND3_X1   g0748(.A1(new_n945), .A2(new_n948), .A3(new_n672), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n672), .B1(new_n945), .B2(new_n948), .ZN(new_n950));
  NOR4_X1   g0750(.A1(new_n700), .A2(new_n949), .A3(new_n719), .A4(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n943), .A2(new_n944), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n720), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n686), .B(KEYINPUT41), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n925), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n954), .ZN(new_n956));
  AOI211_X1 g0756(.A(KEYINPUT108), .B(new_n956), .C1(new_n952), .C2(new_n720), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n955), .A2(new_n957), .A3(new_n723), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n945), .A2(new_n935), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT42), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n923), .A2(KEYINPUT43), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n496), .B1(new_n932), .B2(new_n623), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n667), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n960), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT107), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n964), .B(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n961), .B1(new_n960), .B2(new_n963), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n923), .A2(KEYINPUT43), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n677), .A2(new_n935), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n966), .A2(new_n971), .A3(new_n969), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n924), .B1(new_n958), .B2(new_n975), .ZN(G387));
  NOR2_X1   g0776(.A1(new_n314), .A2(G50), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT50), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n684), .B1(new_n285), .B2(new_n416), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  AOI211_X1 g0779(.A(G45), .B(new_n979), .C1(new_n978), .C2(new_n977), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n731), .B1(new_n243), .B2(new_n275), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n685), .A2(new_n233), .A3(new_n263), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n983), .B1(new_n448), .B2(new_n234), .ZN(new_n984));
  NOR3_X1   g0784(.A1(new_n984), .A2(new_n738), .A3(new_n737), .ZN(new_n985));
  AOI22_X1  g0785(.A1(G311), .A2(new_n773), .B1(new_n746), .B2(G322), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n745), .A2(new_n906), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n986), .B(new_n987), .C1(new_n801), .C2(new_n766), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT48), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n989), .B1(new_n763), .B2(new_n750), .C1(new_n748), .C2(new_n760), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT49), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n803), .A2(G326), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n990), .A2(new_n991), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n263), .B1(new_n776), .B2(G116), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n992), .A2(new_n993), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n263), .B1(new_n766), .B2(new_n285), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n800), .A2(new_n297), .B1(new_n392), .B2(new_n744), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n997), .B(new_n998), .C1(G150), .C2(new_n803), .ZN(new_n999));
  INV_X1    g0799(.A(new_n318), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n776), .A2(G97), .B1(new_n1000), .B2(new_n773), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n761), .A2(new_n208), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n612), .A2(new_n750), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n999), .A2(new_n1001), .A3(new_n1002), .A4(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n783), .B1(new_n996), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n676), .A2(new_n741), .ZN(new_n1007));
  NOR4_X1   g0807(.A1(new_n985), .A2(new_n1006), .A3(new_n728), .A4(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n949), .A2(new_n950), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1008), .B1(new_n1009), .B2(new_n723), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n686), .B(KEYINPUT110), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n951), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n720), .A2(new_n1009), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1010), .B1(new_n1012), .B2(new_n1013), .ZN(G393));
  INV_X1    g0814(.A(new_n1011), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n943), .A2(new_n944), .A3(KEYINPUT111), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(KEYINPUT111), .B2(new_n943), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n952), .B(new_n1015), .C1(new_n1017), .C2(new_n951), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n935), .A2(new_n737), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n739), .B1(new_n444), .B2(new_n233), .C1(new_n253), .C2(new_n919), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n263), .B1(new_n803), .B2(G322), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n801), .B2(new_n756), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n448), .A2(new_n764), .B1(new_n760), .B2(new_n763), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1022), .B(new_n1023), .C1(G116), .C2(new_n908), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n745), .A2(G311), .B1(new_n746), .B2(G317), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT52), .Z(new_n1026));
  OAI211_X1 g0826(.A(new_n1024), .B(new_n1026), .C1(new_n748), .C2(new_n766), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT112), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n756), .A2(new_n392), .ZN(new_n1029));
  INV_X1    g0829(.A(G150), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n800), .A2(new_n1030), .B1(new_n297), .B2(new_n744), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT51), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(G68), .A2(new_n761), .B1(new_n776), .B2(G87), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n263), .B1(new_n753), .B2(new_n808), .C1(new_n314), .C2(new_n766), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n750), .A2(new_n416), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1032), .A2(new_n1033), .A3(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1028), .B1(new_n1029), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n728), .B1(new_n1038), .B2(new_n738), .ZN(new_n1039));
  AND3_X1   g0839(.A1(new_n1019), .A2(new_n1020), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n1017), .B2(new_n723), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1018), .A2(new_n1041), .ZN(G390));
  NAND2_X1  g0842(.A1(new_n881), .A2(new_n875), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n697), .A2(new_n789), .A3(new_n667), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n879), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n858), .A2(new_n1045), .ZN(new_n1046));
  AND2_X1   g0846(.A1(new_n851), .A2(new_n862), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1047), .A2(new_n874), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n873), .A2(new_n1043), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n822), .A2(new_n858), .A3(G330), .A4(new_n789), .ZN(new_n1050));
  OAI21_X1  g0850(.A(KEYINPUT113), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT114), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n719), .A2(new_n1052), .A3(new_n789), .A4(new_n858), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n714), .ZN(new_n1054));
  AOI221_X4 g0854(.A(new_n526), .B1(new_n537), .B2(new_n539), .C1(new_n546), .C2(new_n547), .ZN(new_n1055));
  AND3_X1   g0855(.A1(new_n623), .A2(new_n616), .A3(new_n587), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1055), .A2(new_n930), .A3(new_n1056), .A4(new_n667), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1054), .B1(new_n1057), .B2(KEYINPUT31), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n718), .ZN(new_n1059));
  OAI211_X1 g0859(.A(G330), .B(new_n789), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(KEYINPUT114), .B1(new_n1060), .B2(new_n834), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1053), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1049), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1048), .A2(new_n1046), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n852), .A2(KEYINPUT39), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1047), .A2(new_n871), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n874), .B1(new_n858), .B2(new_n880), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1064), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT113), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1050), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  AND3_X1   g0872(.A1(new_n1051), .A2(new_n1063), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n723), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n305), .B1(new_n753), .B2(new_n748), .C1(new_n444), .C2(new_n766), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(G107), .B2(new_n773), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n744), .A2(new_n206), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1035), .B(new_n1077), .C1(G283), .C2(new_n746), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1076), .A2(new_n1078), .A3(new_n772), .A4(new_n811), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n760), .A2(new_n1030), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT53), .ZN(new_n1081));
  INV_X1    g0881(.A(G128), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n800), .A2(new_n1082), .B1(new_n750), .B2(new_n297), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(G132), .B2(new_n745), .ZN(new_n1084));
  INV_X1    g0884(.A(G125), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n263), .B1(new_n753), .B2(new_n1085), .C1(new_n911), .C2(new_n756), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n776), .B2(G50), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1081), .A2(new_n1084), .A3(new_n1087), .ZN(new_n1088));
  XOR2_X1   g0888(.A(KEYINPUT54), .B(G143), .Z(new_n1089));
  AND2_X1   g0889(.A1(new_n767), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1079), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n728), .B1(new_n1091), .B2(new_n738), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1092), .B1(new_n1000), .B2(new_n817), .C1(new_n1067), .C2(new_n736), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1074), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n822), .A2(G330), .A3(new_n789), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1045), .B1(new_n1095), .B2(new_n834), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1062), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1060), .A2(new_n834), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1050), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n880), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n442), .B(G330), .C1(new_n1058), .C2(new_n820), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n885), .A2(new_n1102), .A3(new_n635), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT115), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n885), .A2(new_n1102), .A3(new_n635), .A4(KEYINPUT115), .ZN(new_n1106));
  AND2_X1   g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1101), .A2(KEYINPUT116), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT116), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1062), .A2(new_n1096), .B1(new_n1099), .B2(new_n880), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1109), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1108), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n1073), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT117), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1113), .A2(new_n1073), .A3(KEYINPUT117), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1113), .A2(new_n1073), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1119), .A2(new_n1011), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1094), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(G378));
  OAI22_X1  g0922(.A1(new_n766), .A2(new_n911), .B1(new_n750), .B2(new_n1030), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n800), .A2(new_n1085), .B1(new_n1082), .B2(new_n744), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n1123), .B(new_n1124), .C1(new_n761), .C2(new_n1089), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n813), .B2(new_n756), .ZN(new_n1126));
  XOR2_X1   g0926(.A(new_n1126), .B(KEYINPUT59), .Z(new_n1127));
  AOI21_X1  g0927(.A(G33), .B1(new_n803), .B2(G124), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  AOI211_X1 g0929(.A(G41), .B(new_n1129), .C1(G159), .C2(new_n776), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(KEYINPUT3), .A2(G33), .ZN(new_n1131));
  AOI21_X1  g0931(.A(G50), .B1(new_n1131), .B2(new_n274), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n764), .A2(new_n216), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT118), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n745), .A2(G107), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n746), .A2(G116), .B1(new_n908), .B2(G68), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1002), .A2(new_n305), .A3(new_n1135), .A4(new_n1136), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n612), .A2(new_n766), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n274), .B1(new_n753), .B2(new_n763), .C1(new_n444), .C2(new_n756), .ZN(new_n1139));
  NOR4_X1   g0939(.A1(new_n1134), .A2(new_n1137), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1140), .B(new_n1141), .ZN(new_n1142));
  NOR3_X1   g0942(.A1(new_n1130), .A2(new_n1132), .A3(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n725), .B1(new_n1143), .B2(new_n783), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n405), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n634), .A2(new_n1145), .ZN(new_n1146));
  XOR2_X1   g0946(.A(new_n1146), .B(KEYINPUT120), .Z(new_n1147));
  NOR2_X1   g0947(.A1(new_n422), .A2(new_n664), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1148), .B(new_n1149), .ZN(new_n1150));
  OR2_X1    g0950(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1144), .B1(new_n1153), .B2(new_n735), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n783), .A2(new_n392), .A3(new_n736), .ZN(new_n1155));
  AND2_X1   g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1153), .B1(new_n866), .B2(G330), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n835), .A2(new_n854), .B1(KEYINPUT40), .B2(new_n864), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1153), .ZN(new_n1159));
  NOR3_X1   g0959(.A1(new_n1158), .A2(new_n701), .A3(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n883), .B1(new_n1157), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1159), .B1(new_n1158), .B2(new_n701), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n866), .A2(G330), .A3(new_n1153), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1162), .B(new_n1163), .C1(new_n876), .C2(new_n882), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1161), .A2(new_n1164), .A3(KEYINPUT121), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT121), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1166), .B(new_n883), .C1(new_n1160), .C2(new_n1157), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1156), .B1(new_n1168), .B2(new_n723), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1111), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1161), .A2(new_n1164), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(KEYINPUT57), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1015), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n1113), .A2(KEYINPUT117), .A3(new_n1073), .ZN(new_n1174));
  AOI21_X1  g0974(.A(KEYINPUT117), .B1(new_n1113), .B2(new_n1073), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1107), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(KEYINPUT57), .B1(new_n1176), .B2(new_n1168), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1169), .B1(new_n1173), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT122), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  OAI211_X1 g0980(.A(KEYINPUT122), .B(new_n1169), .C1(new_n1173), .C2(new_n1177), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(G375));
  NOR2_X1   g0983(.A1(new_n760), .A2(new_n297), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n263), .B1(new_n753), .B2(new_n1082), .C1(new_n1030), .C2(new_n766), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n746), .A2(G132), .B1(new_n908), .B2(G50), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(new_n911), .C2(new_n744), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1134), .B(new_n1188), .C1(new_n773), .C2(new_n1089), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n305), .B1(new_n756), .B2(new_n206), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(G303), .B2(new_n803), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n745), .A2(G283), .B1(new_n746), .B2(G294), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1191), .B(new_n1192), .C1(new_n448), .C2(new_n766), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1004), .B1(new_n444), .B2(new_n760), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1193), .B(new_n1194), .C1(G77), .C2(new_n776), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1189), .A2(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1196), .A2(new_n783), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n725), .B1(G68), .B2(new_n817), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1198), .B(KEYINPUT124), .Z(new_n1199));
  AOI211_X1 g0999(.A(new_n1197), .B(new_n1199), .C1(new_n834), .C2(new_n735), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n1101), .B2(new_n723), .ZN(new_n1201));
  AND3_X1   g1001(.A1(new_n1110), .A2(KEYINPUT123), .A3(new_n1111), .ZN(new_n1202));
  AOI21_X1  g1002(.A(KEYINPUT123), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1112), .B(new_n1108), .C1(new_n1202), .C2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1201), .B1(new_n1204), .B2(new_n956), .ZN(G381));
  NAND3_X1  g1005(.A1(new_n1180), .A2(new_n1121), .A3(new_n1181), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(G393), .A2(G396), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  OR3_X1    g1008(.A1(G387), .A2(G384), .A3(G390), .ZN(new_n1209));
  OR4_X1    g1009(.A1(G381), .A2(new_n1206), .A3(new_n1208), .A4(new_n1209), .ZN(G407));
  INV_X1    g1010(.A(G213), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1211), .A2(G343), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1182), .A2(KEYINPUT125), .A3(new_n1121), .A4(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT125), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1212), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1214), .B1(new_n1206), .B2(new_n1215), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(G407), .A2(new_n1213), .A3(G213), .A4(new_n1216), .ZN(G409));
  NAND3_X1  g1017(.A1(new_n1176), .A2(new_n954), .A3(new_n1168), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1156), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1171), .A2(new_n723), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1218), .A2(new_n1121), .A3(new_n1219), .A4(new_n1220), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n1221), .A2(new_n1215), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1178), .A2(G378), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1110), .A2(KEYINPUT60), .A3(new_n1111), .ZN(new_n1224));
  XOR2_X1   g1024(.A(new_n1224), .B(KEYINPUT126), .Z(new_n1225));
  INV_X1    g1025(.A(KEYINPUT60), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n1113), .A2(new_n1226), .B1(new_n1203), .B2(new_n1202), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1225), .A2(new_n1227), .A3(new_n1015), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1228), .A2(G384), .A3(new_n1201), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(G384), .B1(new_n1228), .B2(new_n1201), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1222), .A2(new_n1223), .A3(new_n1232), .ZN(new_n1233));
  OAI211_X1 g1033(.A(G2897), .B(new_n1212), .C1(new_n1230), .C2(new_n1231), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1231), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1212), .A2(G2897), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1235), .A2(new_n1229), .A3(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1234), .A2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(new_n1223), .B2(new_n1222), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT63), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1233), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT61), .ZN(new_n1242));
  OR2_X1    g1042(.A1(new_n1233), .A2(new_n1240), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n924), .B(G390), .C1(new_n958), .C2(new_n975), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT127), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(G393), .A2(G396), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1246), .A2(new_n1208), .A3(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(G387), .A2(new_n1041), .A3(new_n1018), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n1244), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1248), .A2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1207), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1252), .A2(new_n1244), .A3(new_n1249), .A4(new_n1247), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1251), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1241), .A2(new_n1242), .A3(new_n1243), .A4(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1238), .ZN(new_n1258));
  AOI21_X1  g1058(.A(KEYINPUT61), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT62), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1222), .A2(new_n1223), .A3(new_n1260), .A4(new_n1232), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1233), .A2(KEYINPUT62), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1259), .A2(new_n1261), .A3(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n1254), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1256), .A2(new_n1264), .ZN(G405));
  INV_X1    g1065(.A(new_n1232), .ZN(new_n1266));
  AND3_X1   g1066(.A1(new_n1206), .A2(new_n1254), .A3(new_n1223), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1254), .B1(new_n1206), .B2(new_n1223), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1266), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1206), .A2(new_n1223), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1255), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1206), .A2(new_n1254), .A3(new_n1223), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1271), .A2(new_n1232), .A3(new_n1272), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1269), .A2(new_n1273), .ZN(G402));
endmodule


