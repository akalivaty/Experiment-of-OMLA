//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 0 1 1 1 0 1 0 1 1 0 0 1 1 1 1 0 1 0 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1264, new_n1265, new_n1266, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n209), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT1), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n209), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  INV_X1    g0019(.A(KEYINPUT0), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(G50), .B1(G58), .B2(G68), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(new_n219), .A2(new_n220), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n226), .B1(new_n220), .B2(new_n219), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n217), .A2(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT2), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n233), .B(new_n234), .Z(new_n235));
  XOR2_X1   g0035(.A(new_n232), .B(new_n235), .Z(G358));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT64), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G87), .B(G97), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n202), .A2(G68), .ZN(new_n241));
  INV_X1    g0041(.A(G68), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n240), .B(new_n246), .ZN(G351));
  XNOR2_X1  g0047(.A(KEYINPUT3), .B(G33), .ZN(new_n248));
  INV_X1    g0048(.A(G1698), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n248), .A2(G222), .A3(new_n249), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n248), .A2(G223), .A3(G1698), .ZN(new_n251));
  INV_X1    g0051(.A(G77), .ZN(new_n252));
  OAI211_X1 g0052(.A(new_n250), .B(new_n251), .C1(new_n252), .C2(new_n248), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n221), .B1(G33), .B2(G41), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n256), .B1(G41), .B2(G45), .ZN(new_n257));
  INV_X1    g0057(.A(G274), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(G1), .A3(G13), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n257), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n259), .B1(new_n263), .B2(G226), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n255), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT68), .ZN(new_n267));
  INV_X1    g0067(.A(G179), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n221), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT65), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT65), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n270), .A2(new_n273), .A3(new_n221), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n256), .A2(G13), .A3(G20), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n256), .A2(G20), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G50), .ZN(new_n279));
  XNOR2_X1  g0079(.A(new_n279), .B(KEYINPUT67), .ZN(new_n280));
  OAI22_X1  g0080(.A1(new_n277), .A2(new_n280), .B1(G50), .B2(new_n276), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT8), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(KEYINPUT66), .A3(G58), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT66), .ZN(new_n285));
  INV_X1    g0085(.A(G58), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n285), .B1(KEYINPUT8), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(KEYINPUT8), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n284), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G33), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(G20), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G20), .A2(G33), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n275), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n282), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(KEYINPUT68), .B1(new_n265), .B2(G179), .ZN(new_n298));
  INV_X1    g0098(.A(G169), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n265), .A2(new_n299), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n269), .A2(new_n297), .A3(new_n298), .A4(new_n300), .ZN(new_n301));
  OR2_X1    g0101(.A1(KEYINPUT70), .A2(KEYINPUT9), .ZN(new_n302));
  NAND2_X1  g0102(.A1(KEYINPUT70), .A2(KEYINPUT9), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n282), .A2(new_n302), .A3(new_n296), .A4(new_n303), .ZN(new_n304));
  OAI211_X1 g0104(.A(KEYINPUT70), .B(KEYINPUT9), .C1(new_n281), .C2(new_n295), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT10), .ZN(new_n307));
  INV_X1    g0107(.A(G200), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n308), .B1(new_n255), .B2(new_n264), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n309), .B1(new_n266), .B2(G190), .ZN(new_n310));
  AND3_X1   g0110(.A1(new_n306), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n307), .B1(new_n306), .B2(new_n310), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n301), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n290), .A2(KEYINPUT3), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT3), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G33), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n314), .A2(new_n316), .A3(G226), .A4(G1698), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n314), .A2(new_n316), .A3(G223), .A4(new_n249), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G33), .A2(G87), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n254), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n259), .B1(new_n263), .B2(G232), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n321), .A2(G190), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n308), .B1(new_n321), .B2(new_n322), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n275), .A2(new_n278), .A3(new_n289), .ZN(new_n326));
  INV_X1    g0126(.A(new_n276), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n327), .B(new_n284), .C1(new_n287), .C2(new_n288), .ZN(new_n328));
  AND3_X1   g0128(.A1(new_n326), .A2(KEYINPUT77), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(KEYINPUT77), .B1(new_n326), .B2(new_n328), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT7), .ZN(new_n332));
  NOR3_X1   g0132(.A1(new_n248), .A2(new_n332), .A3(G20), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n314), .A2(new_n316), .ZN(new_n334));
  AOI21_X1  g0134(.A(KEYINPUT7), .B1(new_n334), .B2(new_n222), .ZN(new_n335));
  OAI21_X1  g0135(.A(G68), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  AND2_X1   g0136(.A1(G58), .A2(G68), .ZN(new_n337));
  OAI21_X1  g0137(.A(G20), .B1(new_n337), .B2(new_n201), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT76), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI211_X1 g0140(.A(KEYINPUT76), .B(G20), .C1(new_n337), .C2(new_n201), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n293), .A2(G159), .ZN(new_n342));
  AND3_X1   g0142(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n336), .A2(new_n343), .A3(KEYINPUT16), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT16), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n332), .B1(new_n248), .B2(G20), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n334), .A2(KEYINPUT7), .A3(new_n222), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n242), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n345), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n344), .A2(new_n350), .A3(new_n271), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n325), .A2(new_n331), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT17), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n352), .A2(KEYINPUT17), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n331), .A2(new_n351), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n321), .A2(new_n322), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(G169), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n321), .A2(new_n322), .A3(G179), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AND3_X1   g0160(.A1(new_n356), .A2(KEYINPUT18), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(KEYINPUT18), .B1(new_n356), .B2(new_n360), .ZN(new_n362));
  OAI22_X1  g0162(.A1(new_n354), .A2(new_n355), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n313), .B1(new_n364), .B2(KEYINPUT78), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n248), .A2(G232), .A3(new_n249), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n248), .A2(G238), .A3(G1698), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n366), .B(new_n367), .C1(new_n206), .C2(new_n248), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n254), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT69), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n259), .B1(new_n263), .B2(G244), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n370), .B1(new_n369), .B2(new_n371), .ZN(new_n374));
  OAI21_X1  g0174(.A(G190), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n374), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n376), .A2(G200), .A3(new_n372), .ZN(new_n377));
  INV_X1    g0177(.A(new_n271), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n378), .A2(G77), .A3(new_n278), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(G77), .B2(new_n276), .ZN(new_n380));
  NAND2_X1  g0180(.A1(G20), .A2(G77), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n283), .A2(G58), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n288), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n293), .ZN(new_n384));
  XOR2_X1   g0184(.A(KEYINPUT15), .B(G87), .Z(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n222), .A2(G33), .ZN(new_n387));
  OAI221_X1 g0187(.A(new_n381), .B1(new_n383), .B2(new_n384), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n380), .B1(new_n388), .B2(new_n271), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n375), .A2(new_n377), .A3(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n268), .B1(new_n373), .B2(new_n374), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n376), .A2(new_n299), .A3(new_n372), .ZN(new_n392));
  INV_X1    g0192(.A(new_n389), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT78), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n395), .B1(new_n363), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(G190), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n314), .A2(new_n316), .A3(G232), .A4(G1698), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n314), .A2(new_n316), .A3(G226), .A4(new_n249), .ZN(new_n400));
  AND3_X1   g0200(.A1(KEYINPUT71), .A2(G33), .A3(G97), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT71), .B1(G33), .B2(G97), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n399), .A2(new_n400), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT72), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT72), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n399), .A2(new_n400), .A3(new_n406), .A4(new_n403), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n405), .A2(new_n407), .A3(new_n254), .ZN(new_n408));
  INV_X1    g0208(.A(G238), .ZN(new_n409));
  OAI22_X1  g0209(.A1(new_n262), .A2(new_n409), .B1(new_n258), .B2(new_n257), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT13), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT73), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT13), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n408), .A2(new_n415), .A3(new_n411), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n413), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n412), .A2(KEYINPUT73), .A3(KEYINPUT13), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n398), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n275), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n291), .A2(G77), .B1(G20), .B2(new_n242), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(new_n202), .B2(new_n384), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  XOR2_X1   g0223(.A(KEYINPUT74), .B(KEYINPUT11), .Z(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n420), .A2(new_n422), .A3(new_n424), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n378), .A2(G68), .A3(new_n278), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n327), .A2(KEYINPUT12), .A3(new_n242), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT12), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(new_n276), .B2(G68), .ZN(new_n431));
  AND3_X1   g0231(.A1(new_n428), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n426), .A2(new_n427), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT75), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n426), .A2(KEYINPUT75), .A3(new_n427), .A4(new_n432), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n261), .B1(new_n404), .B2(KEYINPUT72), .ZN(new_n438));
  AOI211_X1 g0238(.A(KEYINPUT13), .B(new_n410), .C1(new_n438), .C2(new_n407), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n415), .B1(new_n408), .B2(new_n411), .ZN(new_n440));
  OAI21_X1  g0240(.A(G200), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n419), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n416), .A2(new_n414), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n444), .A2(new_n440), .ZN(new_n445));
  INV_X1    g0245(.A(new_n418), .ZN(new_n446));
  OAI21_X1  g0246(.A(G179), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(G169), .B1(new_n439), .B2(new_n440), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT14), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT14), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n450), .B(G169), .C1(new_n439), .C2(new_n440), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n447), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n437), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n443), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AND3_X1   g0254(.A1(new_n365), .A2(new_n397), .A3(new_n454), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n314), .A2(new_n316), .A3(G244), .A4(new_n249), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT4), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n248), .A2(KEYINPUT4), .A3(G244), .A4(new_n249), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G33), .A2(G283), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n248), .A2(G250), .A3(G1698), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n458), .A2(new_n459), .A3(new_n460), .A4(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n254), .ZN(new_n463));
  INV_X1    g0263(.A(G41), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n256), .B(G45), .C1(new_n464), .C2(KEYINPUT5), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT5), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(G41), .ZN(new_n467));
  OAI211_X1 g0267(.A(G257), .B(new_n261), .C1(new_n465), .C2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(G45), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(G1), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n464), .A2(KEYINPUT5), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n466), .A2(G41), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n470), .A2(new_n471), .A3(new_n472), .A4(G274), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n463), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT82), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n474), .B1(new_n462), .B2(new_n254), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT82), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n481), .A2(G190), .B1(G200), .B2(new_n476), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT81), .ZN(new_n483));
  AND2_X1   g0283(.A1(G97), .A2(G107), .ZN(new_n484));
  NOR2_X1   g0284(.A1(G97), .A2(G107), .ZN(new_n485));
  OAI22_X1  g0285(.A1(new_n484), .A2(new_n485), .B1(KEYINPUT79), .B2(KEYINPUT6), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G97), .A2(G107), .ZN(new_n487));
  NOR2_X1   g0287(.A1(KEYINPUT79), .A2(KEYINPUT6), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n207), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n205), .A2(KEYINPUT6), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n486), .A2(new_n489), .A3(G20), .A4(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n293), .A2(G77), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT80), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n346), .A2(new_n347), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n493), .A2(new_n494), .B1(new_n495), .B2(G107), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n491), .A2(KEYINPUT80), .A3(new_n492), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n378), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n327), .A2(new_n205), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n256), .A2(G33), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n275), .A2(new_n276), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n499), .B1(new_n501), .B2(new_n205), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n483), .B1(new_n498), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n493), .A2(new_n494), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n495), .A2(G107), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n504), .A2(new_n497), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n271), .ZN(new_n507));
  INV_X1    g0307(.A(new_n502), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n507), .A2(KEYINPUT81), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n476), .A2(G179), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n479), .B1(new_n463), .B2(new_n475), .ZN(new_n512));
  AOI211_X1 g0312(.A(KEYINPUT82), .B(new_n474), .C1(new_n462), .C2(new_n254), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n511), .B1(new_n514), .B2(new_n299), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n507), .A2(new_n508), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n482), .A2(new_n510), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n314), .A2(new_n316), .A3(G244), .A4(G1698), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n314), .A2(new_n316), .A3(G238), .A4(new_n249), .ZN(new_n519));
  NAND2_X1  g0319(.A1(G33), .A2(G116), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n254), .ZN(new_n522));
  INV_X1    g0322(.A(G250), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n523), .B1(new_n256), .B2(G45), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n524), .A2(new_n261), .B1(new_n470), .B2(G274), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n525), .A2(KEYINPUT83), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n261), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n470), .A2(G274), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n527), .A2(KEYINPUT83), .A3(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n522), .B(G190), .C1(new_n526), .C2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT84), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n207), .A2(G87), .ZN(new_n533));
  OAI21_X1  g0333(.A(KEYINPUT19), .B1(new_n401), .B2(new_n402), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n533), .B1(new_n534), .B2(new_n222), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n314), .A2(new_n316), .A3(new_n222), .A4(G68), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n387), .A2(new_n205), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n536), .B1(KEYINPUT19), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n271), .B1(new_n535), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n386), .A2(new_n327), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n275), .A2(G87), .A3(new_n276), .A4(new_n500), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n522), .B1(new_n526), .B2(new_n529), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G200), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n527), .A2(new_n528), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT83), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n525), .A2(KEYINPUT83), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n549), .A2(KEYINPUT84), .A3(G190), .A4(new_n522), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n532), .A2(new_n542), .A3(new_n544), .A4(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n539), .B(new_n540), .C1(new_n386), .C2(new_n501), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n547), .A2(new_n548), .B1(new_n254), .B2(new_n521), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n268), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n552), .B(new_n554), .C1(G169), .C2(new_n553), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT91), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n314), .A2(new_n316), .A3(new_n222), .A4(G87), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT22), .ZN(new_n559));
  OR2_X1    g0359(.A1(new_n559), .A2(KEYINPUT88), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n248), .A2(new_n222), .A3(new_n560), .A4(G87), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(KEYINPUT89), .B1(new_n222), .B2(G107), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(KEYINPUT23), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT23), .ZN(new_n567));
  OAI211_X1 g0367(.A(KEYINPUT89), .B(new_n567), .C1(new_n222), .C2(G107), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n566), .A2(new_n568), .B1(G116), .B2(new_n291), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT24), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n564), .A2(KEYINPUT24), .A3(new_n569), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n572), .A2(new_n271), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n327), .A2(new_n206), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT25), .ZN(new_n576));
  XNOR2_X1  g0376(.A(new_n575), .B(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(new_n206), .B2(new_n501), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n314), .A2(new_n316), .A3(G250), .A4(new_n249), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n314), .A2(new_n316), .A3(G257), .A4(G1698), .ZN(new_n582));
  NAND2_X1  g0382(.A1(G33), .A2(G294), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n254), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n464), .A2(KEYINPUT5), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n256), .A2(G45), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n254), .B1(new_n588), .B2(new_n471), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(G264), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n585), .A2(new_n590), .A3(new_n473), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(G200), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n254), .A2(new_n584), .B1(new_n589), .B2(G264), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n593), .A2(G190), .A3(new_n473), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n557), .B1(new_n580), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n378), .B1(new_n570), .B2(new_n571), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n578), .B1(new_n597), .B2(new_n573), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n598), .A2(KEYINPUT91), .A3(new_n594), .A4(new_n592), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n556), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n276), .A2(G116), .A3(new_n500), .ZN(new_n601));
  INV_X1    g0401(.A(G116), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n601), .A2(new_n378), .B1(new_n602), .B2(new_n327), .ZN(new_n603));
  AOI21_X1  g0403(.A(G20), .B1(G33), .B2(G283), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n290), .A2(G97), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT86), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n604), .A2(new_n605), .A3(KEYINPUT86), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n270), .A2(new_n221), .B1(G20), .B2(new_n602), .ZN(new_n611));
  AOI21_X1  g0411(.A(KEYINPUT20), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n604), .A2(new_n605), .A3(KEYINPUT86), .ZN(new_n613));
  AOI21_X1  g0413(.A(KEYINPUT86), .B1(new_n604), .B2(new_n605), .ZN(new_n614));
  OAI211_X1 g0414(.A(KEYINPUT20), .B(new_n611), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n603), .B1(new_n612), .B2(new_n616), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n314), .A2(new_n316), .A3(G257), .A4(new_n249), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n314), .A2(new_n316), .A3(G264), .A4(G1698), .ZN(new_n619));
  INV_X1    g0419(.A(G303), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n618), .B(new_n619), .C1(new_n620), .C2(new_n248), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n254), .ZN(new_n622));
  OAI211_X1 g0422(.A(G270), .B(new_n261), .C1(new_n465), .C2(new_n467), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n623), .A2(KEYINPUT85), .A3(new_n473), .ZN(new_n624));
  AOI21_X1  g0424(.A(KEYINPUT85), .B1(new_n623), .B2(new_n473), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n622), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n617), .A2(KEYINPUT21), .A3(G169), .A4(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n623), .A2(new_n473), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT85), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n623), .A2(KEYINPUT85), .A3(new_n473), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n630), .A2(new_n631), .B1(new_n254), .B2(new_n621), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n617), .A2(new_n632), .A3(G179), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n627), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n630), .A2(new_n631), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n299), .B1(new_n635), .B2(new_n622), .ZN(new_n636));
  AOI21_X1  g0436(.A(KEYINPUT21), .B1(new_n636), .B2(new_n617), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n603), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n611), .B1(new_n613), .B2(new_n614), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT20), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n639), .B1(new_n642), .B2(new_n615), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n622), .B(G190), .C1(new_n624), .C2(new_n625), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n308), .B1(new_n635), .B2(new_n622), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT87), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n626), .A2(G200), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT87), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n648), .A2(new_n649), .A3(new_n644), .A4(new_n643), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n299), .B1(new_n593), .B2(new_n473), .ZN(new_n652));
  OAI22_X1  g0452(.A1(new_n652), .A2(KEYINPUT90), .B1(new_n268), .B2(new_n591), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n591), .A2(KEYINPUT90), .A3(G169), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n580), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n638), .A2(new_n651), .A3(new_n655), .ZN(new_n656));
  AND4_X1   g0456(.A1(new_n455), .A2(new_n517), .A3(new_n600), .A4(new_n656), .ZN(G372));
  OR2_X1    g0457(.A1(new_n311), .A2(new_n312), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n325), .A2(new_n331), .A3(new_n351), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT17), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n353), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n419), .B2(new_n442), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n449), .A2(new_n451), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n268), .B1(new_n417), .B2(new_n418), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n453), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n663), .B1(new_n666), .B2(new_n394), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n356), .A2(new_n360), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT18), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n356), .A2(KEYINPUT18), .A3(new_n360), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n658), .B1(new_n667), .B2(new_n673), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n674), .A2(new_n301), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n477), .A2(new_n299), .A3(new_n480), .ZN(new_n676));
  INV_X1    g0476(.A(new_n511), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(new_n516), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n482), .A2(new_n510), .ZN(new_n679));
  INV_X1    g0479(.A(new_n637), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n627), .A2(new_n633), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n655), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  AND4_X1   g0482(.A1(new_n678), .A2(new_n600), .A3(new_n679), .A4(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(KEYINPUT81), .B1(new_n507), .B2(new_n508), .ZN(new_n684));
  AOI211_X1 g0484(.A(new_n483), .B(new_n502), .C1(new_n506), .C2(new_n271), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n551), .A2(new_n555), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT26), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n686), .A2(new_n687), .A3(new_n688), .A4(new_n515), .ZN(new_n689));
  OAI21_X1  g0489(.A(KEYINPUT26), .B1(new_n678), .B2(new_n556), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(new_n555), .A3(new_n690), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n683), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n455), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n675), .A2(new_n693), .ZN(G369));
  INV_X1    g0494(.A(G330), .ZN(new_n695));
  INV_X1    g0495(.A(new_n638), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n256), .A2(new_n222), .A3(G13), .ZN(new_n697));
  OR3_X1    g0497(.A1(new_n697), .A2(KEYINPUT92), .A3(KEYINPUT27), .ZN(new_n698));
  OAI21_X1  g0498(.A(KEYINPUT92), .B1(new_n697), .B2(KEYINPUT27), .ZN(new_n699));
  INV_X1    g0499(.A(G213), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n700), .B1(new_n697), .B2(KEYINPUT27), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n698), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  XNOR2_X1  g0503(.A(KEYINPUT93), .B(G343), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n696), .A2(new_n617), .A3(new_n706), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n638), .B(new_n651), .C1(new_n643), .C2(new_n705), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n695), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n596), .A2(new_n599), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n655), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n598), .A2(new_n705), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n655), .ZN(new_n716));
  AOI22_X1  g0516(.A1(new_n713), .A2(new_n715), .B1(new_n716), .B2(new_n706), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n710), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n638), .A2(new_n706), .ZN(new_n720));
  AOI22_X1  g0520(.A1(new_n713), .A2(new_n720), .B1(new_n716), .B2(new_n705), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n719), .A2(new_n721), .ZN(G399));
  INV_X1    g0522(.A(new_n218), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G41), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n533), .A2(new_n602), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n724), .A2(new_n725), .A3(new_n256), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n726), .B1(new_n225), .B2(new_n724), .ZN(new_n727));
  XOR2_X1   g0527(.A(new_n727), .B(KEYINPUT28), .Z(new_n728));
  NAND4_X1  g0528(.A1(new_n600), .A2(new_n682), .A3(new_n679), .A4(new_n678), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n687), .A2(new_n688), .A3(new_n515), .A4(new_n516), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n676), .A2(new_n551), .A3(new_n677), .A4(new_n555), .ZN(new_n731));
  OAI21_X1  g0531(.A(KEYINPUT26), .B1(new_n731), .B2(new_n510), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n729), .A2(new_n555), .A3(new_n730), .A4(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(new_n705), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(KEYINPUT29), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n656), .A2(new_n517), .A3(new_n600), .A4(new_n705), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n632), .A2(G179), .A3(new_n553), .A4(new_n593), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n738), .A2(new_n481), .A3(KEYINPUT30), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n543), .B(KEYINPUT94), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n632), .A2(G179), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n740), .A2(new_n476), .A3(new_n591), .A4(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT30), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(new_n514), .B2(new_n737), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n739), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n745), .A2(KEYINPUT31), .A3(new_n706), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n706), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT31), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n736), .A2(new_n746), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G330), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT29), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n752), .B(new_n705), .C1(new_n683), .C2(new_n691), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n735), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n728), .B1(new_n755), .B2(G1), .ZN(G364));
  AOI21_X1  g0556(.A(new_n221), .B1(G20), .B2(new_n299), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n222), .A2(new_n398), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n268), .A2(G200), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n286), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n268), .A2(new_n308), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n763), .A2(new_n759), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n398), .A2(G20), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(new_n763), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n765), .A2(new_n202), .B1(new_n768), .B2(new_n242), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n308), .A2(G179), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n759), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n762), .B(new_n769), .C1(G87), .C2(new_n772), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n766), .A2(new_n268), .A3(G200), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n248), .B1(new_n775), .B2(new_n252), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n398), .A2(G179), .A3(G200), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n222), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n776), .B1(G97), .B2(new_n779), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n766), .B(KEYINPUT97), .Z(new_n781));
  NOR3_X1   g0581(.A1(new_n781), .A2(G179), .A3(new_n308), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n773), .B(new_n780), .C1(new_n206), .C2(new_n783), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n781), .A2(G179), .A3(G200), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G159), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT32), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n771), .A2(new_n620), .ZN(new_n788));
  INV_X1    g0588(.A(G326), .ZN(new_n789));
  XOR2_X1   g0589(.A(KEYINPUT33), .B(G317), .Z(new_n790));
  OAI22_X1  g0590(.A1(new_n765), .A2(new_n789), .B1(new_n768), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n761), .ZN(new_n792));
  AOI211_X1 g0592(.A(new_n788), .B(new_n791), .C1(G322), .C2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n248), .B1(new_n774), .B2(G311), .ZN(new_n794));
  INV_X1    g0594(.A(G294), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n793), .B(new_n794), .C1(new_n795), .C2(new_n778), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n785), .A2(G329), .ZN(new_n797));
  INV_X1    g0597(.A(G283), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n797), .B1(new_n783), .B2(new_n798), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n784), .A2(new_n787), .B1(new_n796), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT98), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n758), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(new_n801), .B2(new_n800), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n222), .A2(G13), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n256), .B1(new_n804), .B2(G45), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(new_n724), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n723), .A2(new_n334), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n207), .A2(KEYINPUT95), .A3(G87), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT95), .ZN(new_n810));
  NAND2_X1  g0610(.A1(G355), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n808), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n246), .A2(new_n469), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n723), .A2(new_n248), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n814), .B1(G45), .B2(new_n224), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n812), .B1(G116), .B2(new_n218), .C1(new_n813), .C2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT96), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n816), .A2(new_n817), .ZN(new_n819));
  NOR2_X1   g0619(.A1(G13), .A2(G33), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(G20), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(new_n757), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n803), .B(new_n807), .C1(new_n818), .C2(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT99), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n707), .A2(new_n708), .A3(new_n822), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n807), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n707), .A2(new_n695), .A3(new_n708), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n710), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(G396));
  AND2_X1   g0633(.A1(new_n692), .A2(new_n705), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n391), .A2(new_n392), .A3(new_n393), .A4(new_n705), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n389), .A2(new_n705), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT100), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n390), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n836), .B1(new_n839), .B2(new_n394), .ZN(new_n840));
  OR2_X1    g0640(.A1(new_n834), .A2(new_n840), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n705), .B(new_n840), .C1(new_n683), .C2(new_n691), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n807), .B1(new_n843), .B2(new_n751), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n751), .B2(new_n843), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n757), .A2(new_n820), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n829), .B1(new_n252), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n782), .A2(G87), .ZN(new_n848));
  INV_X1    g0648(.A(new_n785), .ZN(new_n849));
  INV_X1    g0649(.A(G311), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n772), .A2(G107), .B1(new_n774), .B2(G116), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n852), .B1(new_n798), .B2(new_n768), .C1(new_n795), .C2(new_n761), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n334), .B1(new_n205), .B2(new_n778), .C1(new_n765), .C2(new_n620), .ZN(new_n854));
  NOR3_X1   g0654(.A1(new_n851), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n764), .A2(G137), .B1(new_n774), .B2(G159), .ZN(new_n856));
  INV_X1    g0656(.A(G143), .ZN(new_n857));
  INV_X1    g0657(.A(G150), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n856), .B1(new_n857), .B2(new_n761), .C1(new_n858), .C2(new_n768), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT34), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n782), .A2(G68), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n785), .A2(G132), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n779), .A2(G58), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n334), .B1(new_n772), .B2(G50), .ZN(new_n864));
  AND4_X1   g0664(.A1(new_n861), .A2(new_n862), .A3(new_n863), .A4(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n855), .B1(new_n860), .B2(new_n865), .ZN(new_n866));
  OAI221_X1 g0666(.A(new_n847), .B1(new_n758), .B2(new_n866), .C1(new_n840), .C2(new_n821), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n845), .A2(new_n867), .ZN(G384));
  NAND3_X1  g0668(.A1(new_n486), .A2(new_n489), .A3(new_n490), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT35), .ZN(new_n870));
  OR2_X1    g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n869), .A2(new_n870), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n871), .A2(G116), .A3(new_n223), .A4(new_n872), .ZN(new_n873));
  XOR2_X1   g0673(.A(new_n873), .B(KEYINPUT36), .Z(new_n874));
  OAI211_X1 g0674(.A(new_n225), .B(G77), .C1(new_n286), .C2(new_n242), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n256), .B(G13), .C1(new_n875), .C2(new_n241), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n443), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n453), .A2(new_n706), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n878), .A2(new_n666), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n452), .A2(new_n453), .A3(new_n706), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n882), .A2(new_n750), .A3(new_n840), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n344), .A2(new_n350), .A3(new_n271), .ZN(new_n884));
  INV_X1    g0684(.A(new_n330), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n326), .A2(KEYINPUT77), .A3(new_n328), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n703), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n668), .A2(new_n888), .A3(new_n352), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT37), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n668), .A2(new_n888), .A3(new_n892), .A4(new_n352), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n363), .A2(new_n889), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  XNOR2_X1  g0694(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT103), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n344), .A2(new_n350), .A3(new_n420), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n702), .B1(new_n331), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n363), .A2(new_n898), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n331), .A2(new_n897), .B1(new_n358), .B2(new_n359), .ZN(new_n900));
  NOR3_X1   g0700(.A1(new_n659), .A2(new_n900), .A3(new_n898), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n893), .B1(new_n901), .B2(new_n892), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n899), .A2(KEYINPUT38), .A3(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT103), .ZN(new_n904));
  INV_X1    g0704(.A(new_n895), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n891), .A2(new_n893), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n888), .B1(new_n672), .B2(new_n662), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n904), .B(new_n905), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n896), .A2(new_n903), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n883), .A2(new_n909), .A3(KEYINPUT40), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT40), .ZN(new_n911));
  INV_X1    g0711(.A(new_n903), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT38), .B1(new_n899), .B2(new_n902), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n882), .A2(new_n750), .A3(new_n840), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n911), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n910), .A2(new_n916), .ZN(new_n917));
  XOR2_X1   g0717(.A(new_n917), .B(KEYINPUT105), .Z(new_n918));
  AND2_X1   g0718(.A1(new_n455), .A2(new_n750), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n695), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n919), .B2(new_n918), .ZN(new_n921));
  INV_X1    g0721(.A(new_n753), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n752), .B1(new_n733), .B2(new_n705), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n455), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n675), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n921), .B(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT39), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n896), .A2(new_n908), .A3(new_n927), .A4(new_n903), .ZN(new_n928));
  OAI21_X1  g0728(.A(KEYINPUT39), .B1(new_n912), .B2(new_n913), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n449), .A2(new_n451), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n437), .B1(new_n931), .B2(new_n447), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n705), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n930), .A2(new_n934), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n454), .A2(new_n879), .B1(new_n932), .B2(new_n706), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n835), .B(KEYINPUT101), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n936), .B1(new_n842), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n913), .B2(new_n912), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n673), .A2(new_n702), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n935), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n941), .B(KEYINPUT104), .Z(new_n942));
  NAND2_X1  g0742(.A1(new_n926), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n256), .B2(new_n804), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n926), .A2(new_n942), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n877), .B1(new_n944), .B2(new_n945), .ZN(G367));
  INV_X1    g0746(.A(new_n814), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n235), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n823), .B1(new_n218), .B2(new_n386), .ZN(new_n949));
  OAI221_X1 g0749(.A(new_n334), .B1(new_n761), .B2(new_n620), .C1(new_n778), .C2(new_n206), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n764), .A2(G311), .B1(new_n774), .B2(G283), .ZN(new_n951));
  INV_X1    g0751(.A(G317), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n951), .B1(new_n795), .B2(new_n768), .C1(new_n849), .C2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n771), .A2(new_n602), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT46), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n783), .A2(new_n205), .ZN(new_n956));
  OR4_X1    g0756(.A1(new_n950), .A2(new_n953), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n334), .B1(new_n782), .B2(G77), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT113), .Z(new_n959));
  INV_X1    g0759(.A(G137), .ZN(new_n960));
  INV_X1    g0760(.A(G159), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n775), .A2(new_n202), .B1(new_n961), .B2(new_n768), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n849), .A2(new_n960), .B1(KEYINPUT112), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(KEYINPUT112), .B2(new_n962), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n778), .A2(new_n242), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n286), .A2(new_n771), .B1(new_n761), .B2(new_n858), .ZN(new_n966));
  AOI211_X1 g0766(.A(new_n965), .B(new_n966), .C1(G143), .C2(new_n764), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n957), .B1(new_n959), .B2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT47), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n757), .B1(new_n969), .B2(new_n970), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n807), .B1(new_n948), .B2(new_n949), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT114), .ZN(new_n974));
  INV_X1    g0774(.A(new_n822), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n542), .A2(new_n705), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n687), .A2(new_n976), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n977), .A2(KEYINPUT106), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(KEYINPUT106), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n976), .A2(new_n555), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n974), .B1(new_n975), .B2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n981), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT43), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n981), .A2(KEYINPUT43), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n679), .B(new_n678), .C1(new_n510), .C2(new_n705), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n510), .A2(new_n705), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n515), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n678), .B1(new_n991), .B2(new_n655), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n696), .A2(new_n705), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n993), .A2(new_n712), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n990), .A2(new_n994), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n992), .A2(new_n705), .B1(KEYINPUT42), .B2(new_n995), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n996), .A2(KEYINPUT107), .B1(KEYINPUT42), .B2(new_n995), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n992), .A2(new_n705), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n995), .A2(KEYINPUT42), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT107), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n985), .B(new_n986), .C1(new_n997), .C2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n995), .A2(KEYINPUT42), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n996), .A2(KEYINPUT107), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1005), .A2(new_n984), .A3(new_n983), .A4(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n719), .A2(new_n991), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1003), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(KEYINPUT108), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n724), .B(KEYINPUT41), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n721), .A2(new_n990), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT45), .ZN(new_n1014));
  XOR2_X1   g0814(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  OR3_X1    g0816(.A1(new_n721), .A2(new_n990), .A3(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1016), .B1(new_n721), .B2(new_n990), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n718), .B1(new_n1014), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT45), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1013), .B(new_n1021), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1022), .A2(new_n719), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT110), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n993), .B1(new_n655), .B2(new_n705), .C1(new_n712), .C2(new_n714), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n994), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1024), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n994), .A2(KEYINPUT110), .ZN(new_n1028));
  OR3_X1    g0828(.A1(new_n1027), .A2(new_n709), .A3(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n709), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1020), .A2(new_n1023), .A3(new_n755), .A4(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1012), .B1(new_n1032), .B2(new_n755), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n1033), .A2(KEYINPUT111), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n805), .B1(new_n1033), .B2(KEYINPUT111), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1010), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1008), .B1(new_n1003), .B2(new_n1007), .ZN(new_n1037));
  AND3_X1   g0837(.A1(new_n1003), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT108), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1037), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n982), .B1(new_n1036), .B2(new_n1041), .ZN(G387));
  INV_X1    g0842(.A(new_n1031), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1043), .A2(KEYINPUT116), .A3(new_n754), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1031), .A2(new_n755), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT116), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n1031), .B2(new_n755), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1044), .A2(new_n724), .A3(new_n1045), .A4(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n334), .B1(new_n849), .B2(new_n789), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n764), .A2(G322), .B1(new_n774), .B2(G303), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n850), .B2(new_n768), .C1(new_n952), .C2(new_n761), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT48), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1052), .B1(new_n798), .B2(new_n778), .C1(new_n795), .C2(new_n771), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT49), .Z(new_n1054));
  AOI211_X1 g0854(.A(new_n1049), .B(new_n1054), .C1(G116), .C2(new_n782), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n768), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n289), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n849), .B2(new_n858), .ZN(new_n1058));
  OR3_X1    g0858(.A1(new_n765), .A2(KEYINPUT115), .A3(new_n961), .ZN(new_n1059));
  OAI21_X1  g0859(.A(KEYINPUT115), .B1(new_n765), .B2(new_n961), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n779), .A2(new_n385), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n771), .A2(new_n252), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(G68), .B2(new_n774), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1064), .B(new_n248), .C1(new_n202), .C2(new_n761), .ZN(new_n1065));
  NOR4_X1   g0865(.A1(new_n1058), .A2(new_n956), .A3(new_n1062), .A4(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n757), .B1(new_n1055), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n717), .A2(new_n822), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n947), .B1(new_n232), .B2(G45), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(new_n725), .B2(new_n808), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT50), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n383), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1071), .B1(new_n1072), .B2(new_n202), .ZN(new_n1073));
  NOR3_X1   g0873(.A1(new_n383), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n469), .B1(new_n242), .B2(new_n252), .ZN(new_n1075));
  NOR4_X1   g0875(.A1(new_n1073), .A2(new_n1074), .A3(new_n725), .A4(new_n1075), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n1070), .A2(new_n1076), .B1(G107), .B2(new_n218), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n829), .B1(new_n1077), .B2(new_n823), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1067), .A2(new_n1068), .A3(new_n1078), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1048), .B(new_n1079), .C1(new_n805), .C2(new_n1043), .ZN(G393));
  NAND2_X1  g0880(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n1045), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1082), .A2(new_n724), .A3(new_n1032), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1020), .A2(new_n1023), .A3(new_n806), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n823), .B1(new_n205), .B2(new_n218), .C1(new_n240), .C2(new_n947), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n807), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n774), .A2(new_n1072), .B1(new_n772), .B2(G68), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n779), .A2(G77), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n334), .B1(new_n1056), .B2(G50), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n765), .A2(new_n858), .B1(new_n761), .B2(new_n961), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT51), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1092), .B(new_n848), .C1(new_n857), .C2(new_n849), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n765), .A2(new_n952), .B1(new_n761), .B2(new_n850), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT52), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n785), .A2(G322), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n1096), .B1(new_n1095), .B2(new_n1094), .C1(new_n206), .C2(new_n783), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n248), .B1(new_n1056), .B2(G303), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n772), .A2(G283), .B1(new_n774), .B2(G294), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1098), .B(new_n1099), .C1(new_n602), .C2(new_n778), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n1090), .A2(new_n1093), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1086), .B1(new_n1101), .B2(new_n757), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n990), .B2(new_n975), .ZN(new_n1103));
  AND2_X1   g0903(.A1(new_n1084), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1083), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT117), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1083), .A2(KEYINPUT117), .A3(new_n1104), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(G390));
  NAND3_X1  g0909(.A1(new_n928), .A2(new_n929), .A3(new_n820), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n846), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n807), .B1(new_n1111), .B2(new_n289), .ZN(new_n1112));
  INV_X1    g0912(.A(G128), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n765), .A2(new_n1113), .B1(new_n768), .B2(new_n960), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(G132), .B2(new_n792), .ZN(new_n1115));
  INV_X1    g0915(.A(G125), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n1115), .B1(new_n783), .B2(new_n202), .C1(new_n1116), .C2(new_n849), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n771), .A2(new_n858), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1118), .B(KEYINPUT53), .ZN(new_n1119));
  XOR2_X1   g0919(.A(KEYINPUT54), .B(G143), .Z(new_n1120));
  AOI21_X1  g0920(.A(new_n334), .B1(new_n774), .B2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1119), .B(new_n1121), .C1(new_n961), .C2(new_n778), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n861), .B1(new_n849), .B2(new_n795), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1056), .A2(G107), .B1(G97), .B2(new_n774), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n792), .A2(G116), .B1(new_n764), .B2(G283), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n248), .B1(new_n772), .B2(G87), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1124), .A2(new_n1125), .A3(new_n1088), .A4(new_n1126), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n1117), .A2(new_n1122), .B1(new_n1123), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1112), .B1(new_n1128), .B2(new_n757), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1110), .A2(new_n1129), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n929), .B(new_n928), .C1(new_n938), .C2(new_n934), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n882), .A2(new_n750), .A3(G330), .A4(new_n840), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n937), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n732), .A2(new_n730), .A3(new_n555), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n706), .B1(new_n1134), .B2(new_n729), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1133), .B1(new_n1135), .B2(new_n840), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n909), .B(new_n933), .C1(new_n1136), .C2(new_n936), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n1131), .A2(new_n1132), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1132), .B1(new_n1131), .B2(new_n1137), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1130), .B1(new_n1141), .B2(new_n805), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n724), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n455), .A2(G330), .A3(new_n750), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n924), .A2(new_n1145), .A3(new_n675), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n750), .A2(G330), .A3(new_n840), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n936), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n1132), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n842), .A2(new_n937), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1148), .A2(new_n1132), .A3(new_n1136), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1146), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1144), .B1(new_n1140), .B2(new_n1154), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n1148), .A2(new_n1132), .A3(new_n1136), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1150), .B1(new_n1148), .B2(new_n1132), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n1138), .A2(new_n1139), .B1(new_n1158), .B2(new_n1146), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT118), .B1(new_n1155), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1131), .A2(new_n1137), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1132), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1131), .A2(new_n1137), .A3(new_n1132), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1154), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  AND4_X1   g0965(.A1(KEYINPUT118), .A2(new_n1159), .A3(new_n1165), .A4(new_n724), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1143), .B1(new_n1160), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT119), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1159), .A2(new_n1165), .A3(new_n724), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT118), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1159), .A2(new_n1165), .A3(KEYINPUT118), .A4(new_n724), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1174), .A2(KEYINPUT119), .A3(new_n1143), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1169), .A2(new_n1175), .ZN(G378));
  NAND2_X1  g0976(.A1(new_n297), .A2(new_n703), .ZN(new_n1177));
  XOR2_X1   g0977(.A(new_n313), .B(new_n1177), .Z(new_n1178));
  XNOR2_X1  g0978(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1178), .B(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1181), .A2(new_n821), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n785), .A2(G124), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(G33), .A2(G41), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1183), .B(new_n1184), .C1(new_n783), .C2(new_n961), .ZN(new_n1185));
  INV_X1    g0985(.A(G132), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n768), .A2(new_n1186), .B1(new_n761), .B2(new_n1113), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(G150), .B2(new_n779), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n772), .A2(new_n1120), .B1(new_n774), .B2(G137), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1188), .B(new_n1189), .C1(new_n1116), .C2(new_n765), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1185), .B1(new_n1190), .B2(KEYINPUT59), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(KEYINPUT59), .B2(new_n1190), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT58), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1063), .B(new_n965), .C1(new_n385), .C2(new_n774), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n782), .A2(G58), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n785), .A2(G283), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n765), .A2(new_n602), .B1(new_n761), .B2(new_n206), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n464), .B(new_n334), .C1(new_n768), .C2(new_n205), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .A4(new_n1199), .ZN(new_n1200));
  AOI211_X1 g1000(.A(G50), .B(new_n1184), .C1(new_n334), .C2(new_n464), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n1200), .B2(new_n1193), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT120), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1192), .B1(new_n1193), .B2(new_n1200), .C1(new_n1202), .C2(new_n1203), .ZN(new_n1204));
  AND2_X1   g1004(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n757), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT121), .ZN(new_n1207));
  OR2_X1    g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n829), .B1(new_n202), .B2(new_n846), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1182), .A2(new_n1211), .ZN(new_n1212));
  AND3_X1   g1012(.A1(new_n910), .A2(new_n916), .A3(G330), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n941), .A2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n910), .A2(new_n916), .A3(G330), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n930), .A2(new_n934), .B1(new_n673), .B2(new_n702), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1215), .B1(new_n1216), .B2(new_n939), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1181), .B1(new_n1214), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n941), .A2(new_n1213), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1216), .A2(new_n1215), .A3(new_n939), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1219), .A2(new_n1220), .A3(new_n1180), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1218), .A2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1212), .B1(new_n1222), .B2(new_n806), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1146), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1165), .A2(new_n1224), .ZN(new_n1225));
  AND3_X1   g1025(.A1(new_n1219), .A2(new_n1220), .A3(new_n1180), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1180), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1225), .B(KEYINPUT57), .C1(new_n1226), .C2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n724), .ZN(new_n1229));
  AOI21_X1  g1029(.A(KEYINPUT57), .B1(new_n1222), .B2(new_n1225), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1223), .B1(new_n1229), .B2(new_n1230), .ZN(G375));
  NOR2_X1   g1031(.A1(new_n1154), .A2(new_n1012), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1152), .A2(new_n1146), .A3(new_n1153), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1158), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n936), .A2(new_n820), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n807), .B1(new_n1111), .B2(G68), .ZN(new_n1237));
  XOR2_X1   g1037(.A(new_n1237), .B(KEYINPUT122), .Z(new_n1238));
  AOI21_X1  g1038(.A(new_n248), .B1(new_n782), .B2(G77), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1239), .B(KEYINPUT123), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n849), .A2(new_n620), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n772), .A2(G97), .B1(new_n764), .B2(G294), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1242), .B1(new_n798), .B2(new_n761), .ZN(new_n1243));
  OAI221_X1 g1043(.A(new_n1061), .B1(new_n206), .B2(new_n775), .C1(new_n602), .C2(new_n768), .ZN(new_n1244));
  NOR4_X1   g1044(.A1(new_n1240), .A2(new_n1241), .A3(new_n1243), .A4(new_n1244), .ZN(new_n1245));
  OR2_X1    g1045(.A1(new_n1245), .A2(KEYINPUT124), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(KEYINPUT124), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n778), .A2(new_n202), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n334), .B(new_n1248), .C1(new_n1056), .C2(new_n1120), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n785), .A2(G128), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n765), .A2(new_n1186), .B1(new_n771), .B2(new_n961), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n775), .A2(new_n858), .B1(new_n960), .B2(new_n761), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1249), .A2(new_n1195), .A3(new_n1250), .A4(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1246), .A2(new_n1247), .A3(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1238), .B1(new_n1255), .B2(new_n757), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1235), .A2(new_n806), .B1(new_n1236), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1234), .A2(new_n1257), .ZN(G381));
  INV_X1    g1058(.A(G375), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1142), .B1(new_n1159), .B2(new_n1155), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  OR4_X1    g1061(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1262));
  OR4_X1    g1062(.A1(G387), .A2(new_n1261), .A3(new_n1262), .A4(G381), .ZN(G407));
  NOR2_X1   g1063(.A1(new_n704), .A2(new_n700), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(new_n1264), .B(KEYINPUT125), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  OAI211_X1 g1066(.A(G407), .B(G213), .C1(new_n1261), .C2(new_n1266), .ZN(G409));
  NOR2_X1   g1067(.A1(new_n1154), .A2(new_n1144), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1158), .A2(KEYINPUT60), .A3(new_n1146), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT60), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1233), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1268), .A2(new_n1269), .A3(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(G384), .A2(new_n1257), .A3(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(G384), .B1(new_n1272), .B2(new_n1257), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(G375), .B1(new_n1169), .B2(new_n1175), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1222), .A2(new_n1011), .A3(new_n1225), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1223), .A2(new_n1278), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1279), .A2(new_n1260), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1266), .B(new_n1276), .C1(new_n1277), .C2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(KEYINPUT62), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT61), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1279), .A2(new_n1260), .ZN(new_n1284));
  AOI21_X1  g1084(.A(KEYINPUT119), .B1(new_n1174), .B2(new_n1143), .ZN(new_n1285));
  AOI211_X1 g1085(.A(new_n1168), .B(new_n1142), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1284), .B1(new_n1287), .B2(G375), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT62), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1288), .A2(new_n1289), .A3(new_n1266), .A4(new_n1276), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT126), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1291), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1272), .A2(new_n1257), .ZN(new_n1293));
  AND2_X1   g1093(.A1(new_n845), .A2(new_n867), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1295), .A2(KEYINPUT126), .A3(new_n1273), .ZN(new_n1296));
  AOI22_X1  g1096(.A1(new_n1292), .A2(new_n1296), .B1(G2897), .B2(new_n1265), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1296), .A2(G2897), .A3(new_n1265), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1280), .B1(G378), .B2(new_n1259), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1299), .B1(new_n1300), .B2(new_n1265), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1282), .A2(new_n1283), .A3(new_n1290), .A4(new_n1301), .ZN(new_n1302));
  OAI211_X1 g1102(.A(new_n982), .B(G390), .C1(new_n1036), .C2(new_n1041), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  OAI211_X1 g1104(.A(new_n1040), .B(new_n1010), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1305));
  AOI21_X1  g1105(.A(G390), .B1(new_n1305), .B2(new_n982), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(G393), .B(new_n832), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  NOR3_X1   g1108(.A1(new_n1304), .A2(new_n1306), .A3(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(G390), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(G387), .A2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1307), .B1(new_n1311), .B2(new_n1303), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1309), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1302), .A2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1288), .A2(new_n1266), .ZN(new_n1316));
  AOI21_X1  g1116(.A(KEYINPUT61), .B1(new_n1316), .B2(new_n1299), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1288), .A2(KEYINPUT63), .A3(new_n1266), .A4(new_n1276), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT63), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1281), .A2(new_n1319), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1317), .A2(new_n1313), .A3(new_n1318), .A4(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1315), .A2(new_n1321), .ZN(G405));
  NAND2_X1  g1122(.A1(G375), .A2(new_n1260), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1323), .B1(new_n1287), .B2(G375), .ZN(new_n1324));
  AND2_X1   g1124(.A1(new_n1324), .A2(new_n1276), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1324), .A2(new_n1276), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  OAI21_X1  g1127(.A(KEYINPUT127), .B1(new_n1309), .B2(new_n1312), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1308), .B1(new_n1304), .B2(new_n1306), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT127), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1311), .A2(new_n1307), .A3(new_n1303), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1329), .A2(new_n1330), .A3(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1328), .A2(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1327), .A2(new_n1333), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1328), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1335));
  AND2_X1   g1135(.A1(new_n1334), .A2(new_n1335), .ZN(G402));
endmodule


