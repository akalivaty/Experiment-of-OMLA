//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1 1 1 1 0 1 0 0 0 0 1 0 0 1 0 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 0 1 1 1 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT72), .ZN(new_n188));
  OR2_X1    g002(.A1(KEYINPUT64), .A2(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT64), .A2(G143), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(G146), .A3(new_n190), .ZN(new_n191));
  AND2_X1   g005(.A1(KEYINPUT0), .A2(G128), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(new_n192), .A3(new_n194), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n193), .A2(G143), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT64), .B(G143), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n196), .B1(new_n197), .B2(new_n193), .ZN(new_n198));
  NOR2_X1   g012(.A1(KEYINPUT0), .A2(G128), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n192), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n195), .B1(new_n198), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G137), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G134), .ZN(new_n204));
  AND2_X1   g018(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n205));
  NOR2_X1   g019(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n203), .A2(KEYINPUT11), .A3(G134), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT66), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n204), .B(KEYINPUT66), .C1(new_n205), .C2(new_n206), .ZN(new_n211));
  INV_X1    g025(.A(G134), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G137), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n210), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G131), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT67), .B(G131), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n210), .A2(new_n211), .A3(new_n213), .A4(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n202), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G128), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n191), .A2(new_n194), .A3(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n219), .B1(new_n194), .B2(KEYINPUT1), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n221), .B1(new_n198), .B2(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n203), .A2(G134), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT68), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n213), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n225), .A2(new_n204), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G131), .ZN(new_n229));
  AND3_X1   g043(.A1(new_n223), .A2(new_n217), .A3(new_n229), .ZN(new_n230));
  XOR2_X1   g044(.A(G116), .B(G119), .Z(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT69), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT2), .B(G113), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n232), .B(new_n234), .ZN(new_n235));
  NOR3_X1   g049(.A1(new_n218), .A2(new_n230), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT71), .ZN(new_n237));
  INV_X1    g051(.A(G953), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(KEYINPUT71), .A2(G953), .ZN(new_n240));
  AND2_X1   g054(.A1(KEYINPUT70), .A2(G237), .ZN(new_n241));
  NOR2_X1   g055(.A1(KEYINPUT70), .A2(G237), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n239), .B(new_n240), .C1(new_n241), .C2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G210), .ZN(new_n244));
  OR3_X1    g058(.A1(new_n243), .A2(KEYINPUT27), .A3(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT27), .B1(new_n243), .B2(new_n244), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT26), .B(G101), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n247), .B(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n188), .B1(new_n236), .B2(new_n250), .ZN(new_n251));
  NOR3_X1   g065(.A1(new_n218), .A2(new_n230), .A3(KEYINPUT30), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT30), .ZN(new_n253));
  INV_X1    g067(.A(new_n202), .ZN(new_n254));
  AND4_X1   g068(.A1(new_n211), .A2(new_n210), .A3(new_n213), .A4(new_n216), .ZN(new_n255));
  INV_X1    g069(.A(G131), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n224), .B1(new_n207), .B2(new_n209), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n256), .B1(new_n257), .B2(new_n211), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n254), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n223), .A2(new_n217), .A3(new_n229), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n253), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n235), .B1(new_n252), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT31), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n247), .B(new_n248), .ZN(new_n264));
  INV_X1    g078(.A(new_n235), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n259), .A2(new_n265), .A3(new_n260), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n264), .A2(new_n266), .A3(KEYINPUT72), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n251), .A2(new_n262), .A3(new_n263), .A4(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT73), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n268), .B(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n265), .B1(new_n259), .B2(new_n260), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT28), .B1(new_n236), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(KEYINPUT74), .B1(new_n236), .B2(KEYINPUT28), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT74), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT28), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n266), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n272), .A2(new_n273), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n250), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n251), .A2(new_n262), .A3(new_n267), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT31), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  OAI211_X1 g095(.A(KEYINPUT32), .B(new_n187), .C1(new_n270), .C2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT75), .ZN(new_n283));
  AND3_X1   g097(.A1(new_n264), .A2(new_n266), .A3(KEYINPUT72), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT30), .B1(new_n218), .B2(new_n230), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n259), .A2(new_n253), .A3(new_n260), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n265), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n288), .A2(new_n269), .A3(new_n263), .A4(new_n251), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n268), .A2(KEYINPUT73), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI22_X1  g105(.A1(KEYINPUT31), .A2(new_n279), .B1(new_n277), .B2(new_n250), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n187), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT32), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n272), .A2(new_n273), .A3(new_n264), .A4(new_n276), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT29), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n250), .B1(new_n287), .B2(new_n236), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G902), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n300), .B(new_n301), .C1(new_n298), .C2(new_n297), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G472), .ZN(new_n303));
  INV_X1    g117(.A(new_n187), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n304), .B1(new_n291), .B2(new_n292), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT75), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(new_n306), .A3(KEYINPUT32), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n283), .A2(new_n296), .A3(new_n303), .A4(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G125), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n309), .A2(G140), .ZN(new_n310));
  XNOR2_X1  g124(.A(G125), .B(G140), .ZN(new_n311));
  MUX2_X1   g125(.A(new_n310), .B(new_n311), .S(KEYINPUT16), .Z(new_n312));
  OR2_X1    g126(.A1(new_n312), .A2(new_n193), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT23), .ZN(new_n314));
  INV_X1    g128(.A(G119), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n314), .B1(new_n315), .B2(G128), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n219), .A2(KEYINPUT23), .A3(G119), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n316), .B(new_n317), .C1(G119), .C2(new_n219), .ZN(new_n318));
  XNOR2_X1  g132(.A(G119), .B(G128), .ZN(new_n319));
  XOR2_X1   g133(.A(KEYINPUT24), .B(G110), .Z(new_n320));
  OAI22_X1  g134(.A1(new_n318), .A2(G110), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n311), .A2(new_n193), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n313), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n312), .B(G146), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n318), .A2(G110), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n320), .A2(new_n319), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n323), .B1(new_n324), .B2(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT22), .B(G137), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n329), .B(KEYINPUT76), .ZN(new_n330));
  XOR2_X1   g144(.A(KEYINPUT71), .B(G953), .Z(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(G221), .A3(G234), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n330), .B(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n328), .B(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT77), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT25), .ZN(new_n337));
  AOI21_X1  g151(.A(G902), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n336), .A2(new_n337), .ZN(new_n340));
  OR2_X1    g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G234), .ZN(new_n342));
  OAI21_X1  g156(.A(G217), .B1(new_n342), .B2(G902), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n343), .B1(new_n339), .B2(new_n340), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n301), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  AOI22_X1  g160(.A1(new_n341), .A2(new_n344), .B1(new_n335), .B2(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT9), .B(G234), .ZN(new_n348));
  OAI21_X1  g162(.A(G221), .B1(new_n348), .B2(G902), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(KEYINPUT79), .B(G469), .ZN(new_n351));
  AND2_X1   g165(.A1(KEYINPUT64), .A2(G143), .ZN(new_n352));
  NOR2_X1   g166(.A1(KEYINPUT64), .A2(G143), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n193), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n219), .B1(new_n354), .B2(KEYINPUT1), .ZN(new_n355));
  INV_X1    g169(.A(new_n194), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n352), .A2(new_n353), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n356), .B1(new_n357), .B2(G146), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n221), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G104), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT3), .B1(new_n360), .B2(G107), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT3), .ZN(new_n362));
  INV_X1    g176(.A(G107), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(new_n363), .A3(G104), .ZN(new_n364));
  INV_X1    g178(.A(G101), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n360), .A2(G107), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n361), .A2(new_n364), .A3(new_n365), .A4(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n360), .A2(G107), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n363), .A2(G104), .ZN(new_n369));
  OAI21_X1  g183(.A(G101), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n359), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT10), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n255), .A2(new_n258), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n361), .A2(new_n364), .A3(new_n366), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G101), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n378), .A2(KEYINPUT4), .A3(new_n367), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n354), .B1(G143), .B2(new_n193), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n200), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT4), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n377), .A2(new_n382), .A3(G101), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n379), .A2(new_n195), .A3(new_n381), .A4(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n223), .A2(new_n372), .A3(KEYINPUT10), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n375), .A2(new_n376), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n215), .A2(new_n217), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n191), .A2(new_n194), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT1), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n389), .B1(new_n197), .B2(new_n193), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n388), .B1(new_n390), .B2(new_n219), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n371), .B1(new_n391), .B2(new_n221), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n223), .A2(new_n372), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n387), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT12), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT12), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n387), .B(new_n396), .C1(new_n392), .C2(new_n393), .ZN(new_n397));
  XNOR2_X1  g211(.A(G110), .B(G140), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n398), .B(KEYINPUT78), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n331), .A2(G227), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n399), .B(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  AND4_X1   g216(.A1(new_n386), .A2(new_n395), .A3(new_n397), .A4(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n384), .A2(new_n385), .ZN(new_n404));
  AOI21_X1  g218(.A(KEYINPUT10), .B1(new_n359), .B2(new_n372), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n387), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n402), .B1(new_n406), .B2(new_n386), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n301), .B(new_n351), .C1(new_n403), .C2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT80), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n406), .A2(new_n386), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n401), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n395), .A2(new_n386), .A3(new_n397), .A4(new_n402), .ZN(new_n413));
  AOI21_X1  g227(.A(G902), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n414), .A2(KEYINPUT80), .A3(new_n351), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n410), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n395), .A2(new_n386), .A3(new_n397), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n401), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n406), .A2(new_n386), .A3(new_n402), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n301), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G469), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n350), .B1(new_n416), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(G214), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n357), .B1(new_n243), .B2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT70), .B(G237), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n331), .A2(G143), .A3(G214), .A4(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n216), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(KEYINPUT84), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT17), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT84), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n428), .A2(new_n433), .A3(new_n429), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n425), .A2(new_n427), .A3(new_n216), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n431), .A2(new_n432), .A3(new_n434), .A4(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n433), .B1(new_n428), .B2(new_n429), .ZN(new_n437));
  AOI211_X1 g251(.A(KEYINPUT84), .B(new_n216), .C1(new_n425), .C2(new_n427), .ZN(new_n438));
  OAI21_X1  g252(.A(KEYINPUT17), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n436), .A2(new_n324), .A3(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(G113), .B(G122), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n441), .B(new_n360), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n311), .B(KEYINPUT83), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(G146), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n322), .ZN(new_n445));
  AND2_X1   g259(.A1(KEYINPUT18), .A2(G131), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n445), .B1(new_n428), .B2(new_n446), .ZN(new_n447));
  AND2_X1   g261(.A1(new_n428), .A2(new_n446), .ZN(new_n448));
  OR2_X1    g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n440), .A2(new_n442), .A3(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n442), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n443), .A2(KEYINPUT19), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT19), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n311), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n452), .A2(new_n193), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n313), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n437), .A2(new_n438), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n456), .B1(new_n457), .B2(new_n435), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n447), .A2(new_n448), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n451), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n450), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g275(.A1(G475), .A2(G902), .ZN(new_n462));
  NAND2_X1  g276(.A1(KEYINPUT85), .A2(KEYINPUT20), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n461), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n462), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n466), .B1(new_n450), .B2(new_n460), .ZN(new_n467));
  NOR2_X1   g281(.A1(KEYINPUT85), .A2(KEYINPUT20), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n465), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(G475), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n440), .A2(new_n449), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n451), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n450), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n472), .B1(new_n475), .B2(new_n301), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(G122), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G116), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT86), .B1(new_n478), .B2(G116), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT86), .ZN(new_n481));
  INV_X1    g295(.A(G116), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n481), .A2(new_n482), .A3(G122), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT14), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n480), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n484), .B1(new_n480), .B2(new_n483), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n479), .B(new_n485), .C1(new_n486), .C2(KEYINPUT88), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n486), .A2(KEYINPUT88), .ZN(new_n488));
  OAI21_X1  g302(.A(G107), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n480), .A2(new_n483), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n490), .A2(new_n363), .A3(new_n479), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n197), .A2(new_n219), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n219), .A2(G143), .ZN(new_n493));
  OAI21_X1  g307(.A(G134), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n493), .B1(new_n357), .B2(G128), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n212), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n491), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(KEYINPUT89), .B1(new_n489), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n489), .A2(new_n497), .A3(KEYINPUT89), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT87), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n495), .A2(KEYINPUT13), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT13), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n357), .A2(new_n504), .A3(G128), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n503), .A2(G134), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n363), .B1(new_n490), .B2(new_n479), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n496), .B1(new_n491), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n502), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  OR2_X1    g323(.A1(new_n491), .A2(new_n507), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n503), .A2(G134), .A3(new_n505), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n510), .A2(new_n511), .A3(KEYINPUT87), .A4(new_n496), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(G217), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n348), .A2(new_n514), .A3(G953), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n501), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n515), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n489), .A2(new_n497), .A3(KEYINPUT89), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n518), .A2(new_n498), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n509), .A2(new_n512), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(G902), .B1(new_n516), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(G478), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n523), .A2(KEYINPUT15), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  AOI211_X1 g340(.A(G902), .B(new_n524), .C1(new_n516), .C2(new_n521), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n238), .A2(G952), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n529), .B1(G234), .B2(G237), .ZN(new_n530));
  XNOR2_X1  g344(.A(KEYINPUT21), .B(G898), .ZN(new_n531));
  XOR2_X1   g345(.A(new_n531), .B(KEYINPUT90), .Z(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  AOI211_X1 g347(.A(new_n301), .B(new_n331), .C1(G234), .C2(G237), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n530), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(G214), .B1(G237), .B2(G902), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n254), .A2(G125), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n223), .A2(new_n309), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(G224), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n542), .A2(G953), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n541), .B(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT5), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(new_n315), .A3(G116), .ZN(new_n547));
  OAI211_X1 g361(.A(G113), .B(new_n547), .C1(new_n231), .C2(new_n546), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n548), .B1(new_n231), .B2(new_n233), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n549), .A2(new_n371), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n235), .A2(new_n383), .A3(new_n379), .ZN(new_n552));
  XNOR2_X1  g366(.A(G110), .B(G122), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n551), .A2(new_n552), .ZN(new_n555));
  XOR2_X1   g369(.A(new_n553), .B(KEYINPUT81), .Z(new_n556));
  AOI22_X1  g370(.A1(new_n554), .A2(KEYINPUT6), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n555), .A2(KEYINPUT6), .A3(new_n556), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n545), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n541), .A2(KEYINPUT7), .A3(new_n544), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n553), .B(KEYINPUT8), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n549), .A2(new_n371), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n561), .B1(new_n562), .B2(new_n550), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n544), .A2(KEYINPUT7), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n539), .A2(new_n540), .A3(new_n564), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n560), .A2(new_n554), .A3(new_n563), .A4(new_n565), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n566), .A2(new_n301), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n559), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(G210), .B1(G237), .B2(G902), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(KEYINPUT82), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n559), .A2(new_n567), .A3(new_n569), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n538), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n477), .A2(new_n528), .A3(new_n536), .A4(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n308), .A2(new_n347), .A3(new_n423), .A4(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(G101), .ZN(G3));
  NAND2_X1  g391(.A1(new_n516), .A2(new_n521), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n521), .A2(KEYINPUT91), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n578), .A2(new_n579), .A3(KEYINPUT33), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT33), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n516), .B(new_n521), .C1(KEYINPUT91), .C2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n580), .A2(G478), .A3(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n523), .A2(new_n301), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n584), .B1(new_n522), .B2(new_n523), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n583), .B(new_n585), .C1(new_n471), .C2(new_n476), .ZN(new_n586));
  INV_X1    g400(.A(new_n569), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n541), .B(new_n543), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n554), .A2(KEYINPUT6), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n555), .A2(new_n556), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n555), .A2(KEYINPUT6), .A3(new_n556), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n588), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n566), .A2(new_n301), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n587), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n538), .B1(new_n595), .B2(new_n572), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n536), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT92), .B1(new_n586), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n583), .A2(new_n585), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  AOI211_X1 g414(.A(new_n535), .B(new_n538), .C1(new_n595), .C2(new_n572), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT92), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n440), .A2(new_n442), .A3(new_n449), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n442), .B1(new_n440), .B2(new_n449), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n301), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(G475), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n461), .A2(new_n462), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n469), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n606), .A2(new_n608), .A3(new_n465), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n600), .A2(new_n601), .A3(new_n602), .A4(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n598), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(G472), .ZN(new_n612));
  AOI21_X1  g426(.A(G902), .B1(new_n291), .B2(new_n292), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n294), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n416), .A2(new_n422), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n615), .A2(new_n347), .A3(new_n349), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n611), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT34), .B(G104), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G6));
  INV_X1    g434(.A(new_n596), .ZN(new_n621));
  NOR4_X1   g435(.A1(new_n621), .A2(new_n609), .A3(new_n528), .A4(new_n535), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n617), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT35), .B(G107), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT93), .B(KEYINPUT94), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G9));
  NOR2_X1   g441(.A1(new_n333), .A2(KEYINPUT36), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n328), .B(new_n628), .ZN(new_n629));
  AOI22_X1  g443(.A1(new_n341), .A2(new_n344), .B1(new_n346), .B2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n423), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n614), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n575), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT37), .B(G110), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G12));
  NOR2_X1   g451(.A1(new_n467), .A2(new_n470), .ZN(new_n638));
  AOI211_X1 g452(.A(new_n466), .B(new_n463), .C1(new_n450), .C2(new_n460), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n578), .A2(new_n301), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n524), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n522), .A2(new_n525), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(G900), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n530), .B1(new_n534), .B2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n640), .A2(new_n644), .A3(new_n606), .A4(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(KEYINPUT95), .B1(new_n649), .B2(new_n596), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT95), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n648), .A2(new_n651), .A3(new_n621), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n308), .B(new_n633), .C1(new_n650), .C2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G128), .ZN(G30));
  NAND2_X1  g468(.A1(new_n615), .A2(new_n349), .ZN(new_n655));
  XOR2_X1   g469(.A(new_n646), .B(KEYINPUT39), .Z(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  OR2_X1    g473(.A1(new_n659), .A2(KEYINPUT40), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n250), .B1(new_n236), .B2(new_n271), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n279), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g476(.A(G472), .B1(new_n662), .B2(G902), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n283), .A2(new_n296), .A3(new_n307), .A4(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n659), .A2(KEYINPUT40), .ZN(new_n665));
  INV_X1    g479(.A(new_n572), .ZN(new_n666));
  INV_X1    g480(.A(new_n570), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n667), .B1(new_n559), .B2(new_n567), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT38), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n609), .A2(new_n644), .A3(new_n537), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n670), .A2(new_n631), .A3(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n660), .A2(new_n664), .A3(new_n665), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(new_n197), .ZN(G45));
  AND4_X1   g488(.A1(new_n306), .A2(new_n293), .A3(KEYINPUT32), .A4(new_n187), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n306), .B1(new_n305), .B2(KEYINPUT32), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI22_X1  g491(.A1(new_n294), .A2(new_n295), .B1(G472), .B2(new_n302), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n632), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT96), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n680), .B1(new_n586), .B2(new_n646), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n600), .A2(KEYINPUT96), .A3(new_n609), .A4(new_n647), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n681), .A2(new_n596), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT97), .B(G146), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G48));
  INV_X1    g500(.A(G469), .ZN(new_n687));
  OR2_X1    g501(.A1(new_n414), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n408), .A2(new_n409), .ZN(new_n689));
  AOI21_X1  g503(.A(KEYINPUT80), .B1(new_n414), .B2(new_n351), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n349), .B(new_n688), .C1(new_n689), .C2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n691), .A2(KEYINPUT98), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT98), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n414), .A2(new_n687), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n694), .B1(new_n410), .B2(new_n415), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n693), .B1(new_n695), .B2(new_n349), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n611), .A2(new_n308), .A3(new_n347), .A4(new_n697), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT41), .B(G113), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(KEYINPUT99), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n698), .B(new_n700), .ZN(G15));
  NAND4_X1  g515(.A1(new_n308), .A2(new_n347), .A3(new_n697), .A4(new_n622), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G116), .ZN(G18));
  NAND2_X1  g517(.A1(new_n691), .A2(KEYINPUT98), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n695), .A2(new_n693), .A3(new_n349), .ZN(new_n705));
  AND3_X1   g519(.A1(new_n704), .A2(new_n596), .A3(new_n705), .ZN(new_n706));
  NOR4_X1   g520(.A1(new_n630), .A2(new_n609), .A3(new_n644), .A4(new_n535), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n706), .A2(new_n308), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G119), .ZN(G21));
  NOR2_X1   g523(.A1(new_n613), .A2(new_n612), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n187), .B(KEYINPUT100), .ZN(new_n711));
  AOI21_X1  g525(.A(KEYINPUT101), .B1(new_n293), .B2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT101), .ZN(new_n713));
  INV_X1    g527(.A(new_n711), .ZN(new_n714));
  AOI211_X1 g528(.A(new_n713), .B(new_n714), .C1(new_n291), .C2(new_n292), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n710), .A2(new_n712), .A3(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n609), .A2(new_n644), .A3(new_n536), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n706), .A2(new_n716), .A3(new_n347), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G122), .ZN(G24));
  AOI21_X1  g534(.A(new_n714), .B1(new_n291), .B2(new_n292), .ZN(new_n721));
  OAI22_X1  g535(.A1(KEYINPUT101), .A2(new_n721), .B1(new_n613), .B2(new_n612), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n722), .A2(new_n630), .A3(new_n715), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n723), .A2(new_n681), .A3(new_n682), .A4(new_n706), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G125), .ZN(G27));
  AND2_X1   g539(.A1(new_n681), .A2(new_n682), .ZN(new_n726));
  INV_X1    g540(.A(new_n347), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n727), .B1(new_n678), .B2(new_n282), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n350), .A2(new_n538), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT103), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n419), .B(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n418), .A2(KEYINPUT102), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT102), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n417), .A2(new_n733), .A3(new_n401), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n731), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n687), .B1(new_n735), .B2(new_n301), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n689), .A2(new_n690), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n669), .B(new_n729), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n726), .A2(KEYINPUT42), .A3(new_n728), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n308), .A2(new_n347), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n739), .A2(new_n681), .A3(new_n682), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n740), .B1(new_n743), .B2(KEYINPUT42), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G131), .ZN(G33));
  NOR2_X1   g559(.A1(new_n738), .A2(new_n648), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n308), .A2(new_n746), .A3(new_n347), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G134), .ZN(G36));
  INV_X1    g562(.A(KEYINPUT45), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n735), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n687), .B1(new_n420), .B2(new_n749), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(G469), .A2(G902), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT46), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI22_X1  g570(.A1(new_n750), .A2(new_n751), .B1(G469), .B2(G902), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(KEYINPUT46), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n756), .A2(new_n416), .A3(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(new_n349), .A3(new_n656), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(KEYINPUT104), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n666), .A2(new_n538), .A3(new_n668), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g577(.A(KEYINPUT105), .B1(new_n609), .B2(new_n599), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT43), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n764), .A2(new_n765), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(new_n614), .A3(new_n631), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT44), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n763), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI211_X1 g585(.A(new_n761), .B(new_n771), .C1(new_n770), .C2(new_n769), .ZN(new_n772));
  XNOR2_X1  g586(.A(KEYINPUT106), .B(G137), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n772), .B(new_n773), .ZN(G39));
  OR2_X1    g588(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n775));
  NAND2_X1  g589(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n776));
  AOI22_X1  g590(.A1(new_n759), .A2(new_n349), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n416), .B1(new_n757), .B2(KEYINPUT46), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n752), .A2(KEYINPUT46), .A3(new_n753), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n349), .B(new_n776), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  AND3_X1   g596(.A1(new_n726), .A2(new_n727), .A3(new_n762), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n782), .A2(new_n678), .A3(new_n677), .A4(new_n783), .ZN(new_n784));
  XOR2_X1   g598(.A(KEYINPUT108), .B(G140), .Z(new_n785));
  XNOR2_X1  g599(.A(new_n784), .B(new_n785), .ZN(G42));
  NOR2_X1   g600(.A1(G952), .A2(G953), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n724), .A2(new_n653), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n595), .A2(new_n572), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n609), .A2(new_n644), .A3(new_n537), .A4(new_n789), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n647), .A2(KEYINPUT112), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n350), .B1(new_n647), .B2(KEYINPUT112), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n630), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n736), .A2(new_n737), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n790), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n664), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n308), .A2(new_n633), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n681), .A2(new_n596), .A3(new_n682), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT52), .ZN(new_n800));
  OR3_X1    g614(.A1(new_n788), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n802), .B(new_n800), .C1(new_n788), .C2(new_n799), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n684), .A2(new_n653), .A3(new_n724), .A4(new_n796), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n802), .B1(new_n805), .B2(new_n800), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n801), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n642), .A2(new_n643), .A3(new_n647), .ZN(new_n808));
  OAI21_X1  g622(.A(KEYINPUT110), .B1(new_n609), .B2(new_n808), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n526), .A2(new_n527), .A3(new_n646), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT110), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n810), .A2(new_n640), .A3(new_n811), .A4(new_n606), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n809), .A2(new_n762), .A3(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n813), .A2(new_n308), .A3(new_n633), .ZN(new_n814));
  INV_X1    g628(.A(new_n723), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n814), .B(new_n747), .C1(new_n815), .C2(new_n742), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT111), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n726), .A2(new_n723), .A3(new_n739), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n819), .A2(KEYINPUT111), .A3(new_n747), .A4(new_n814), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  AND4_X1   g635(.A1(new_n698), .A2(new_n719), .A3(new_n702), .A4(new_n708), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n574), .A2(new_n614), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n573), .A2(new_n536), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n640), .A2(new_n644), .A3(new_n606), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n824), .B1(new_n586), .B2(new_n825), .ZN(new_n826));
  AOI22_X1  g640(.A1(new_n633), .A2(new_n823), .B1(new_n617), .B2(new_n826), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n827), .A2(KEYINPUT109), .A3(new_n576), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT109), .B1(new_n827), .B2(new_n576), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n822), .B(new_n744), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n821), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n807), .A2(new_n831), .A3(KEYINPUT53), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT53), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n800), .B1(new_n788), .B2(new_n799), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n801), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n698), .A2(new_n719), .A3(new_n702), .A4(new_n708), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT109), .ZN(new_n837));
  INV_X1    g651(.A(new_n576), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n617), .A2(new_n826), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n635), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n837), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n827), .A2(KEYINPUT109), .A3(new_n576), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n836), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n818), .A2(new_n820), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n843), .A2(new_n844), .A3(new_n744), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n833), .B1(new_n835), .B2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n832), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n805), .A2(new_n800), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n834), .A2(KEYINPUT113), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n850), .B1(new_n851), .B2(new_n803), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n833), .B1(new_n852), .B2(new_n845), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT114), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n801), .A2(new_n834), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n831), .A2(new_n856), .A3(KEYINPUT53), .ZN(new_n857));
  OAI211_X1 g671(.A(KEYINPUT114), .B(new_n833), .C1(new_n852), .C2(new_n845), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n855), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n849), .B1(new_n859), .B2(KEYINPUT54), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n766), .A2(new_n530), .A3(new_n767), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n697), .A2(new_n762), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(KEYINPUT117), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n347), .A2(new_n530), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n862), .A2(new_n664), .A3(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n600), .A2(new_n609), .ZN(new_n867));
  AOI22_X1  g681(.A1(new_n864), .A2(new_n723), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n695), .A2(new_n350), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n869), .B1(new_n777), .B2(new_n781), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT118), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n861), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n722), .A2(new_n727), .A3(new_n715), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n873), .A2(new_n874), .A3(new_n762), .ZN(new_n875));
  OAI211_X1 g689(.A(KEYINPUT118), .B(new_n869), .C1(new_n777), .C2(new_n781), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n872), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n697), .A2(new_n538), .A3(new_n670), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n873), .A2(new_n874), .A3(new_n878), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n879), .B(KEYINPUT50), .Z(new_n880));
  NAND4_X1  g694(.A1(new_n868), .A2(new_n877), .A3(new_n880), .A4(KEYINPUT51), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n864), .A2(new_n728), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(KEYINPUT48), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT48), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n864), .A2(new_n884), .A3(new_n728), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n873), .A2(new_n706), .A3(new_n874), .ZN(new_n887));
  INV_X1    g701(.A(new_n586), .ZN(new_n888));
  AOI211_X1 g702(.A(new_n529), .B(new_n887), .C1(new_n888), .C2(new_n866), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n881), .A2(new_n886), .A3(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT115), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n782), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(KEYINPUT115), .B1(new_n777), .B2(new_n781), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n892), .A2(new_n893), .A3(new_n869), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(new_n875), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(KEYINPUT116), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT116), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n894), .A2(new_n897), .A3(new_n875), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n896), .A2(new_n898), .A3(new_n880), .A4(new_n868), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT51), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n890), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n787), .B1(new_n860), .B2(new_n901), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n670), .A2(new_n347), .A3(new_n729), .ZN(new_n903));
  INV_X1    g717(.A(new_n664), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n609), .A2(new_n599), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n695), .B(KEYINPUT49), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n903), .A2(new_n904), .A3(new_n905), .A4(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(KEYINPUT119), .B1(new_n902), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n858), .A2(new_n857), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n807), .A2(new_n831), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT114), .B1(new_n911), .B2(new_n833), .ZN(new_n912));
  OAI21_X1  g726(.A(KEYINPUT54), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n901), .A2(new_n913), .A3(new_n848), .ZN(new_n914));
  INV_X1    g728(.A(new_n787), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT119), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n916), .A2(new_n917), .A3(new_n907), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n909), .A2(new_n918), .ZN(G75));
  NOR2_X1   g733(.A1(new_n331), .A2(G952), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n557), .A2(new_n558), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(new_n588), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n559), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT55), .Z(new_n924));
  NAND2_X1  g738(.A1(new_n832), .A2(new_n846), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n925), .A2(G210), .A3(G902), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT56), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n924), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n925), .A2(G902), .A3(new_n570), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n924), .A2(new_n927), .ZN(new_n930));
  AOI211_X1 g744(.A(new_n920), .B(new_n928), .C1(new_n929), .C2(new_n930), .ZN(G51));
  NAND2_X1  g745(.A1(new_n925), .A2(KEYINPUT54), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n848), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n753), .B(KEYINPUT57), .ZN(new_n935));
  OAI22_X1  g749(.A1(new_n934), .A2(new_n935), .B1(new_n407), .B2(new_n403), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n925), .A2(G902), .ZN(new_n937));
  OR2_X1    g751(.A1(new_n937), .A2(new_n752), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n920), .B1(new_n936), .B2(new_n938), .ZN(G54));
  INV_X1    g753(.A(KEYINPUT58), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n937), .A2(new_n940), .A3(new_n472), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n941), .A2(new_n461), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n941), .A2(new_n461), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n942), .A2(new_n943), .A3(new_n920), .ZN(G60));
  XNOR2_X1  g758(.A(new_n584), .B(KEYINPUT59), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n945), .B1(new_n580), .B2(new_n582), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n920), .B1(new_n933), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n945), .B1(new_n913), .B2(new_n848), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n580), .A2(new_n582), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT120), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n947), .B(KEYINPUT120), .C1(new_n948), .C2(new_n949), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(G63));
  NAND2_X1  g768(.A1(G217), .A2(G902), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT121), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT60), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n925), .A2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n335), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n920), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n925), .A2(new_n629), .A3(new_n957), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT122), .ZN(new_n962));
  AOI22_X1  g776(.A1(new_n960), .A2(new_n961), .B1(new_n962), .B2(KEYINPUT61), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n962), .A2(KEYINPUT61), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n963), .B(new_n964), .ZN(G66));
  INV_X1    g779(.A(new_n843), .ZN(new_n966));
  AOI21_X1  g780(.A(KEYINPUT123), .B1(new_n966), .B2(new_n331), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n966), .A2(KEYINPUT123), .A3(new_n331), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n238), .B1(new_n532), .B2(G224), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT124), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n973), .B(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n921), .B1(G898), .B2(new_n331), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n975), .B(new_n976), .Z(G69));
  NOR2_X1   g791(.A1(new_n252), .A2(new_n261), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n452), .A2(new_n454), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n978), .B(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(new_n645), .B2(new_n331), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n772), .A2(new_n784), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n744), .A2(new_n747), .ZN(new_n983));
  INV_X1    g797(.A(new_n684), .ZN(new_n984));
  AOI211_X1 g798(.A(new_n727), .B(new_n790), .C1(new_n678), .C2(new_n282), .ZN(new_n985));
  AOI211_X1 g799(.A(new_n984), .B(new_n788), .C1(new_n761), .C2(new_n985), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n982), .A2(new_n983), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n981), .B1(new_n987), .B2(new_n331), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n673), .A2(new_n653), .A3(new_n684), .A4(new_n724), .ZN(new_n989));
  OR2_X1    g803(.A1(new_n989), .A2(KEYINPUT62), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(KEYINPUT62), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n763), .B1(new_n586), .B2(new_n825), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n308), .A2(new_n347), .A3(new_n658), .A4(new_n992), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n982), .A2(new_n990), .A3(new_n991), .A4(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n980), .B1(new_n994), .B2(new_n331), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n988), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n331), .B1(G227), .B2(G900), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n996), .B(new_n997), .Z(G72));
  NOR2_X1   g812(.A1(new_n287), .A2(new_n236), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(new_n250), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT127), .Z(new_n1001));
  NAND4_X1  g815(.A1(new_n982), .A2(new_n843), .A3(new_n983), .A4(new_n986), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT126), .ZN(new_n1003));
  NAND2_X1  g817(.A1(G472), .A2(G902), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1004), .B(KEYINPUT63), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT125), .ZN(new_n1006));
  AND3_X1   g820(.A1(new_n1002), .A2(new_n1003), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1003), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1001), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1006), .B1(new_n994), .B2(new_n966), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n999), .A2(new_n250), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n920), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1005), .B1(new_n279), .B2(new_n299), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1013), .B1(new_n859), .B2(new_n1014), .ZN(G57));
endmodule


