//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 1 1 1 1 1 1 1 0 0 1 0 1 0 1 0 1 1 1 0 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n827, new_n828,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  XOR2_X1   g001(.A(KEYINPUT71), .B(G211gat), .Z(new_n203));
  INV_X1    g002(.A(G218gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(KEYINPUT70), .B(KEYINPUT22), .Z(new_n206));
  OAI21_X1  g005(.A(new_n202), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n208), .B(new_n202), .C1(new_n205), .C2(new_n206), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT25), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT24), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n215), .A2(G183gat), .A3(G190gat), .ZN(new_n216));
  XNOR2_X1  g015(.A(G183gat), .B(G190gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n216), .B1(new_n217), .B2(new_n215), .ZN(new_n218));
  INV_X1    g017(.A(G169gat), .ZN(new_n219));
  INV_X1    g018(.A(G176gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(new_n220), .A3(KEYINPUT23), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT23), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n222), .B1(G169gat), .B2(G176gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n221), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n214), .B1(new_n218), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT65), .ZN(new_n227));
  INV_X1    g026(.A(G183gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G190gat), .ZN(new_n229));
  INV_X1    g028(.A(G190gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G183gat), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n215), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n216), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n227), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  OAI211_X1 g033(.A(KEYINPUT65), .B(new_n216), .C1(new_n217), .C2(new_n215), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n223), .A2(KEYINPUT25), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT64), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n221), .A2(new_n238), .A3(new_n224), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n238), .B1(new_n221), .B2(new_n224), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n237), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n226), .B1(new_n236), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(G226gat), .A2(G233gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n219), .A2(new_n220), .A3(KEYINPUT66), .ZN(new_n244));
  OR2_X1    g043(.A1(new_n244), .A2(KEYINPUT26), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(KEYINPUT26), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(new_n224), .A3(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT27), .B(G183gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n230), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT28), .ZN(new_n250));
  NAND2_X1  g049(.A1(G183gat), .A2(G190gat), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT28), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n248), .A2(new_n252), .A3(new_n230), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n247), .A2(new_n250), .A3(new_n251), .A4(new_n253), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n242), .A2(new_n243), .A3(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT29), .B1(G226gat), .B2(G233gat), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n256), .B1(new_n242), .B2(new_n254), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n213), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n242), .A2(new_n243), .A3(new_n254), .ZN(new_n259));
  INV_X1    g058(.A(new_n240), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n221), .A2(new_n238), .A3(new_n224), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n262), .A2(new_n234), .A3(new_n237), .A4(new_n235), .ZN(new_n263));
  AND3_X1   g062(.A1(new_n250), .A2(new_n251), .A3(new_n253), .ZN(new_n264));
  AOI22_X1  g063(.A1(new_n263), .A2(new_n226), .B1(new_n264), .B2(new_n247), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n259), .B(new_n212), .C1(new_n265), .C2(new_n256), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n258), .A2(KEYINPUT72), .A3(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT72), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n268), .B(new_n213), .C1(new_n255), .C2(new_n257), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G8gat), .B(G36gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT73), .ZN(new_n272));
  XNOR2_X1  g071(.A(G64gat), .B(G92gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT75), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT30), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n274), .B1(new_n267), .B2(new_n269), .ZN(new_n280));
  OAI21_X1  g079(.A(KEYINPUT75), .B1(new_n280), .B2(KEYINPUT30), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n270), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n274), .B(KEYINPUT74), .ZN(new_n284));
  AOI22_X1  g083(.A1(new_n283), .A2(new_n284), .B1(new_n280), .B2(KEYINPUT30), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G1gat), .B(G29gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n288), .B(KEYINPUT0), .ZN(new_n289));
  XNOR2_X1  g088(.A(G57gat), .B(G85gat), .ZN(new_n290));
  XOR2_X1   g089(.A(new_n289), .B(new_n290), .Z(new_n291));
  INV_X1    g090(.A(G120gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(G113gat), .ZN(new_n293));
  INV_X1    g092(.A(G113gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(G120gat), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT1), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G134gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(G127gat), .ZN(new_n298));
  INV_X1    g097(.A(G127gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G134gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT67), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT67), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n298), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n296), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G113gat), .B(G120gat), .ZN(new_n306));
  NOR3_X1   g105(.A1(new_n301), .A2(new_n306), .A3(KEYINPUT1), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(G141gat), .A2(G148gat), .ZN(new_n309));
  AND2_X1   g108(.A1(G141gat), .A2(G148gat), .ZN(new_n310));
  NOR2_X1   g109(.A1(G155gat), .A2(G162gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT2), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G155gat), .A2(G162gat), .ZN(new_n314));
  AOI211_X1 g113(.A(new_n309), .B(new_n310), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT76), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n317), .B1(new_n310), .B2(new_n309), .ZN(new_n318));
  INV_X1    g117(.A(G141gat), .ZN(new_n319));
  INV_X1    g118(.A(G148gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(G141gat), .A2(G148gat), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n321), .A2(KEYINPUT76), .A3(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n318), .A2(new_n323), .A3(new_n312), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT77), .ZN(new_n325));
  INV_X1    g124(.A(new_n314), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n326), .A2(new_n311), .ZN(new_n327));
  AND3_X1   g126(.A1(new_n324), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n325), .B1(new_n324), .B2(new_n327), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n308), .B(new_n316), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT4), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n324), .A2(new_n327), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT77), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n324), .A2(new_n325), .A3(new_n327), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT4), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n335), .A2(new_n336), .A3(new_n316), .A4(new_n308), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n331), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n316), .B1(new_n328), .B2(new_n329), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT3), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT3), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n335), .A2(new_n341), .A3(new_n316), .ZN(new_n342));
  OAI21_X1  g141(.A(KEYINPUT78), .B1(new_n305), .B2(new_n307), .ZN(new_n343));
  INV_X1    g142(.A(new_n304), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n303), .B1(new_n298), .B2(new_n300), .ZN(new_n345));
  OAI22_X1  g144(.A1(new_n344), .A2(new_n345), .B1(KEYINPUT1), .B2(new_n306), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT78), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n296), .A2(new_n298), .A3(new_n300), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n343), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n340), .A2(new_n342), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT5), .ZN(new_n352));
  NAND2_X1  g151(.A1(G225gat), .A2(G233gat), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n338), .A2(new_n351), .A3(new_n352), .A4(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT81), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT79), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n331), .A2(new_n356), .A3(new_n337), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n330), .A2(KEYINPUT79), .A3(KEYINPUT4), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n357), .A2(new_n351), .A3(new_n358), .A4(new_n353), .ZN(new_n359));
  INV_X1    g158(.A(new_n353), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT80), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n339), .A2(new_n350), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(new_n330), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n361), .B1(new_n339), .B2(new_n350), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n360), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  AND4_X1   g164(.A1(new_n355), .A2(new_n359), .A3(KEYINPUT5), .A4(new_n365), .ZN(new_n366));
  NOR3_X1   g165(.A1(new_n305), .A2(KEYINPUT78), .A3(new_n307), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n347), .B1(new_n346), .B2(new_n348), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n315), .B1(new_n333), .B2(new_n334), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT80), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n371), .A2(new_n330), .A3(new_n362), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n352), .B1(new_n372), .B2(new_n360), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n355), .B1(new_n373), .B2(new_n359), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n291), .B(new_n354), .C1(new_n366), .C2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT6), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n359), .A2(KEYINPUT5), .A3(new_n365), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT81), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n373), .A2(new_n355), .A3(new_n359), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n291), .B1(new_n381), .B2(new_n354), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n354), .B1(new_n366), .B2(new_n374), .ZN(new_n384));
  INV_X1    g183(.A(new_n291), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(KEYINPUT6), .A3(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n287), .B1(new_n383), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n242), .A2(new_n254), .ZN(new_n389));
  INV_X1    g188(.A(new_n308), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n389), .B(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(G227gat), .ZN(new_n392));
  INV_X1    g191(.A(G233gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT34), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT68), .ZN(new_n398));
  INV_X1    g197(.A(new_n394), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n265), .A2(new_n390), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n389), .A2(new_n308), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n396), .B(new_n399), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n397), .B1(new_n398), .B2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(G15gat), .B(G43gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(G71gat), .B(G99gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n404), .B(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n394), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT33), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n407), .A2(KEYINPUT32), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n407), .B(KEYINPUT32), .C1(new_n408), .C2(new_n406), .ZN(new_n412));
  OR2_X1    g211(.A1(new_n402), .A2(new_n398), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n403), .A2(new_n411), .A3(new_n412), .A4(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT69), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n411), .A2(new_n412), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n402), .A2(new_n398), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n413), .B(new_n417), .C1(new_n396), .C2(new_n395), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n414), .A2(new_n415), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n416), .A2(KEYINPUT69), .A3(new_n418), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(G78gat), .B(G106gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n424), .B(G22gat), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT29), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n212), .B1(new_n342), .B2(new_n427), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n428), .A2(KEYINPUT84), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(G228gat), .A2(G233gat), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n428), .A2(KEYINPUT84), .ZN(new_n432));
  INV_X1    g231(.A(new_n211), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT29), .B1(new_n433), .B2(KEYINPUT83), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT83), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n210), .A2(new_n435), .A3(new_n211), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT3), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  OR2_X1    g236(.A1(new_n437), .A2(new_n370), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n430), .A2(new_n431), .A3(new_n432), .A4(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n341), .B1(new_n213), .B2(KEYINPUT29), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n339), .ZN(new_n441));
  INV_X1    g240(.A(new_n428), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n431), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT31), .B(G50gat), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n439), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n446), .B1(new_n439), .B2(new_n444), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n426), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n449), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n451), .A2(new_n425), .A3(new_n447), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT35), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n450), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NOR3_X1   g253(.A1(new_n388), .A2(new_n423), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT82), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n388), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n384), .A2(new_n385), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n458), .A2(new_n376), .A3(new_n375), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n386), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n460), .A2(KEYINPUT82), .A3(new_n287), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n450), .A2(new_n452), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n414), .A2(new_n419), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n457), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n455), .B1(new_n465), .B2(KEYINPUT35), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT86), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n371), .A2(new_n330), .A3(new_n353), .A4(new_n362), .ZN(new_n468));
  AND2_X1   g267(.A1(new_n338), .A2(new_n351), .ZN(new_n469));
  OAI211_X1 g268(.A(KEYINPUT39), .B(new_n468), .C1(new_n469), .C2(new_n353), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n353), .B1(new_n338), .B2(new_n351), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT39), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n385), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT40), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n474), .B1(new_n384), .B2(new_n385), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n470), .A2(new_n473), .A3(KEYINPUT40), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT85), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT85), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n470), .A2(new_n473), .A3(new_n478), .A4(KEYINPUT40), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  AND4_X1   g279(.A1(new_n467), .A2(new_n475), .A3(new_n286), .A4(new_n480), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n282), .A2(new_n285), .B1(new_n477), .B2(new_n479), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n467), .B1(new_n482), .B2(new_n475), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT87), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n258), .A2(new_n266), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT37), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT38), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(new_n488), .A3(new_n284), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT37), .B1(new_n267), .B2(new_n269), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n276), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n283), .A2(KEYINPUT37), .ZN(new_n492));
  INV_X1    g291(.A(new_n490), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n492), .A2(new_n274), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n491), .B1(new_n494), .B2(KEYINPUT38), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n459), .A2(new_n386), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n462), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NOR3_X1   g297(.A1(new_n484), .A2(new_n485), .A3(new_n498), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n496), .A2(new_n497), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n475), .A2(new_n286), .A3(new_n480), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT86), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n482), .A2(new_n467), .A3(new_n475), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT87), .B1(new_n500), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n499), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT36), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n420), .A2(new_n507), .A3(new_n421), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n414), .A2(KEYINPUT36), .A3(new_n419), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n457), .A2(new_n461), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n511), .B1(new_n512), .B2(new_n462), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n466), .B1(new_n506), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT88), .ZN(new_n517));
  OR3_X1    g316(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT88), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n517), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT89), .ZN(new_n522));
  AOI22_X1  g321(.A1(new_n521), .A2(new_n522), .B1(G29gat), .B2(G36gat), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n523), .B1(new_n522), .B2(new_n521), .ZN(new_n524));
  XOR2_X1   g323(.A(G43gat), .B(G50gat), .Z(new_n525));
  INV_X1    g324(.A(KEYINPUT15), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n527), .B1(G29gat), .B2(G36gat), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT90), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n516), .B1(new_n518), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n531), .B1(new_n530), .B2(new_n518), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n525), .A2(new_n526), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n529), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n528), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(KEYINPUT17), .ZN(new_n536));
  XNOR2_X1  g335(.A(G15gat), .B(G22gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(KEYINPUT91), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT92), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(G8gat), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT16), .ZN(new_n541));
  AOI21_X1  g340(.A(G1gat), .B1(new_n538), .B2(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n540), .B(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n536), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(G229gat), .A2(G233gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n543), .A2(new_n535), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT18), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n545), .A2(KEYINPUT18), .A3(new_n546), .A4(new_n547), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n543), .B(new_n535), .ZN(new_n552));
  XOR2_X1   g351(.A(new_n546), .B(KEYINPUT13), .Z(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n550), .A2(new_n551), .A3(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G113gat), .B(G141gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(G197gat), .ZN(new_n557));
  XOR2_X1   g356(.A(KEYINPUT11), .B(G169gat), .Z(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n559), .B(KEYINPUT12), .Z(new_n560));
  NAND2_X1  g359(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n560), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n550), .A2(new_n562), .A3(new_n551), .A4(new_n554), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  XOR2_X1   g364(.A(G57gat), .B(G64gat), .Z(new_n566));
  AND2_X1   g365(.A1(G71gat), .A2(G78gat), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n566), .B1(KEYINPUT9), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT93), .ZN(new_n569));
  NOR2_X1   g368(.A1(G71gat), .A2(G78gat), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n567), .A2(new_n570), .ZN(new_n572));
  OR2_X1    g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n572), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT21), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(G231gat), .A2(G233gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(G127gat), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n544), .B1(new_n577), .B2(new_n576), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(G155gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(G183gat), .B(G211gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n583), .B(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(G232gat), .A2(G233gat), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n590), .A2(KEYINPUT41), .ZN(new_n591));
  XNOR2_X1  g390(.A(G134gat), .B(G162gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(KEYINPUT95), .B(KEYINPUT7), .Z(new_n595));
  INV_X1    g394(.A(KEYINPUT94), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n596), .A2(G85gat), .A3(G92gat), .ZN(new_n597));
  OR2_X1    g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(G99gat), .A2(G106gat), .ZN(new_n599));
  INV_X1    g398(.A(G85gat), .ZN(new_n600));
  INV_X1    g399(.A(G92gat), .ZN(new_n601));
  AOI22_X1  g400(.A1(KEYINPUT8), .A2(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(G99gat), .B(G106gat), .Z(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(KEYINPUT96), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n595), .A2(new_n597), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n598), .A2(new_n602), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n603), .A2(KEYINPUT96), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n606), .A2(new_n607), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n536), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT97), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT97), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n536), .A2(new_n613), .A3(new_n610), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(G190gat), .B(G218gat), .Z(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n535), .B1(new_n608), .B2(new_n609), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n590), .A2(KEYINPUT41), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n615), .A2(new_n617), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n617), .B1(new_n615), .B2(new_n621), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n594), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n624), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n626), .A2(new_n593), .A3(new_n622), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n576), .A2(new_n610), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT10), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n575), .B1(new_n608), .B2(new_n609), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(KEYINPUT98), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n631), .A2(new_n630), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT98), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n629), .A2(new_n635), .A3(new_n630), .A4(new_n631), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n633), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT99), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(G230gat), .A2(G233gat), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n633), .A2(KEYINPUT99), .A3(new_n634), .A4(new_n636), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n629), .A2(new_n631), .ZN(new_n643));
  INV_X1    g442(.A(new_n640), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(G120gat), .B(G148gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(G176gat), .B(G204gat), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n646), .B(new_n647), .Z(new_n648));
  NAND3_X1  g447(.A1(new_n642), .A2(new_n645), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n637), .A2(new_n640), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n645), .ZN(new_n651));
  INV_X1    g450(.A(new_n648), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n589), .A2(new_n628), .A3(new_n655), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n514), .A2(new_n565), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n460), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g459(.A1(new_n657), .A2(new_n286), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n661), .A2(KEYINPUT100), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(KEYINPUT100), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n662), .A2(G8gat), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT101), .ZN(new_n665));
  XOR2_X1   g464(.A(KEYINPUT16), .B(G8gat), .Z(new_n666));
  NAND4_X1  g465(.A1(new_n657), .A2(KEYINPUT42), .A3(new_n286), .A4(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n666), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n668), .B1(new_n662), .B2(new_n663), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n665), .B(new_n667), .C1(KEYINPUT42), .C2(new_n669), .ZN(G1325gat));
  NOR2_X1   g469(.A1(new_n514), .A2(new_n565), .ZN(new_n671));
  INV_X1    g470(.A(new_n656), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(G15gat), .B1(new_n673), .B2(new_n510), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n423), .A2(G15gat), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n674), .B1(new_n673), .B2(new_n675), .ZN(G1326gat));
  NAND2_X1  g475(.A1(new_n657), .A2(new_n462), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT43), .B(G22gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1327gat));
  NAND2_X1  g478(.A1(new_n588), .A2(new_n655), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n680), .A2(new_n628), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n671), .A2(new_n681), .ZN(new_n682));
  OR3_X1    g481(.A1(new_n682), .A2(G29gat), .A3(new_n460), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT45), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n685), .B1(new_n514), .B2(new_n628), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n485), .B1(new_n484), .B2(new_n498), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n500), .A2(new_n504), .A3(KEYINPUT87), .ZN(new_n688));
  AOI21_X1  g487(.A(KEYINPUT82), .B1(new_n460), .B2(new_n287), .ZN(new_n689));
  AOI211_X1 g488(.A(new_n456), .B(new_n286), .C1(new_n459), .C2(new_n386), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n462), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n687), .A2(new_n688), .A3(new_n691), .A4(new_n510), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n465), .A2(KEYINPUT35), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n692), .B1(new_n693), .B2(new_n455), .ZN(new_n694));
  INV_X1    g493(.A(new_n628), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n694), .A2(KEYINPUT44), .A3(new_n695), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n686), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n680), .A2(new_n565), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(G29gat), .B1(new_n699), .B2(new_n460), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(KEYINPUT102), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT102), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n684), .A2(new_n703), .A3(new_n700), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(G1328gat));
  OR2_X1    g504(.A1(new_n287), .A2(G36gat), .ZN(new_n706));
  OAI22_X1  g505(.A1(new_n682), .A2(new_n706), .B1(KEYINPUT103), .B2(KEYINPUT46), .ZN(new_n707));
  NAND2_X1  g506(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n708));
  XOR2_X1   g507(.A(new_n707), .B(new_n708), .Z(new_n709));
  OAI21_X1  g508(.A(G36gat), .B1(new_n699), .B2(new_n287), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(G1329gat));
  NAND2_X1  g510(.A1(new_n511), .A2(G43gat), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n682), .A2(new_n423), .ZN(new_n713));
  OAI22_X1  g512(.A1(new_n699), .A2(new_n712), .B1(G43gat), .B2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g514(.A1(KEYINPUT105), .A2(KEYINPUT48), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n462), .A2(G50gat), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT104), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n462), .B1(new_n682), .B2(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(KEYINPUT104), .B1(new_n671), .B2(new_n681), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OAI221_X1 g520(.A(new_n716), .B1(new_n699), .B2(new_n717), .C1(new_n721), .C2(G50gat), .ZN(new_n722));
  OR2_X1    g521(.A1(KEYINPUT105), .A2(KEYINPUT48), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1331gat));
  NOR4_X1   g523(.A1(new_n588), .A2(new_n695), .A3(new_n564), .A4(new_n655), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n694), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(new_n658), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g528(.A1(new_n726), .A2(new_n287), .ZN(new_n730));
  NOR2_X1   g529(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(KEYINPUT49), .B(G64gat), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n732), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT106), .ZN(G1333gat));
  OR3_X1    g534(.A1(new_n726), .A2(G71gat), .A3(new_n423), .ZN(new_n736));
  OAI21_X1  g535(.A(G71gat), .B1(new_n726), .B2(new_n510), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n738), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g538(.A1(new_n727), .A2(new_n462), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g540(.A1(new_n589), .A2(new_n564), .A3(new_n655), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n686), .A2(new_n696), .A3(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT107), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n686), .A2(new_n696), .A3(KEYINPUT107), .A4(new_n742), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n745), .A2(new_n658), .A3(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n589), .A2(new_n564), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n694), .A2(new_n695), .A3(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT51), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n749), .A2(KEYINPUT108), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n694), .A2(KEYINPUT51), .A3(new_n695), .A4(new_n748), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n751), .B1(new_n754), .B2(KEYINPUT108), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n658), .A2(new_n600), .A3(new_n654), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT109), .ZN(new_n757));
  OAI22_X1  g556(.A1(new_n747), .A2(new_n600), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT110), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n758), .B(new_n759), .ZN(G1336gat));
  NAND4_X1  g559(.A1(new_n686), .A2(new_n696), .A3(new_n286), .A4(new_n742), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT52), .B1(new_n761), .B2(G92gat), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n655), .A2(G92gat), .A3(new_n287), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n762), .B1(new_n755), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n764), .B1(new_n752), .B2(new_n753), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n745), .A2(new_n286), .A3(new_n746), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n766), .B1(new_n767), .B2(G92gat), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n765), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(KEYINPUT111), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT111), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n772), .B(new_n765), .C1(new_n768), .C2(new_n769), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(G1337gat));
  AND3_X1   g573(.A1(new_n745), .A2(new_n511), .A3(new_n746), .ZN(new_n775));
  XNOR2_X1  g574(.A(KEYINPUT112), .B(G99gat), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n422), .A2(new_n654), .A3(new_n776), .ZN(new_n777));
  OAI22_X1  g576(.A1(new_n775), .A2(new_n776), .B1(new_n755), .B2(new_n777), .ZN(G1338gat));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n779));
  OAI21_X1  g578(.A(G106gat), .B1(new_n743), .B2(new_n497), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n655), .A2(new_n497), .A3(G106gat), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n779), .B(new_n780), .C1(new_n755), .C2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT114), .ZN(new_n784));
  XOR2_X1   g583(.A(new_n781), .B(KEYINPUT113), .Z(new_n785));
  AOI21_X1  g584(.A(new_n784), .B1(new_n754), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n754), .A2(new_n785), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n787), .A2(KEYINPUT114), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n745), .A2(new_n462), .A3(new_n746), .ZN(new_n789));
  AOI211_X1 g588(.A(new_n786), .B(new_n788), .C1(G106gat), .C2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n783), .B1(new_n790), .B2(new_n779), .ZN(G1339gat));
  NOR2_X1   g590(.A1(new_n656), .A2(new_n564), .ZN(new_n792));
  INV_X1    g591(.A(new_n649), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT54), .ZN(new_n795));
  INV_X1    g594(.A(new_n637), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n795), .B1(new_n796), .B2(new_n644), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n642), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n652), .B1(new_n650), .B2(KEYINPUT54), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n794), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n799), .B1(new_n642), .B2(new_n797), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n804), .A2(KEYINPUT115), .A3(KEYINPUT55), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n793), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n552), .A2(new_n553), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n546), .B1(new_n545), .B2(new_n547), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n559), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n563), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n801), .A2(new_n802), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n806), .A2(new_n695), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  AOI22_X1  g611(.A1(new_n801), .A2(new_n802), .B1(new_n561), .B2(new_n563), .ZN(new_n813));
  AOI22_X1  g612(.A1(new_n806), .A2(new_n813), .B1(new_n654), .B2(new_n810), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n812), .B1(new_n814), .B2(new_n695), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n792), .B1(new_n815), .B2(new_n588), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n816), .A2(new_n462), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n817), .A2(new_n658), .A3(new_n287), .A4(new_n422), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n818), .A2(new_n294), .A3(new_n565), .ZN(new_n819));
  INV_X1    g618(.A(new_n464), .ZN(new_n820));
  NOR4_X1   g619(.A1(new_n816), .A2(new_n460), .A3(new_n286), .A4(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(G113gat), .B1(new_n821), .B2(new_n564), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n819), .A2(new_n822), .ZN(G1340gat));
  NOR3_X1   g622(.A1(new_n818), .A2(new_n292), .A3(new_n655), .ZN(new_n824));
  AOI21_X1  g623(.A(G120gat), .B1(new_n821), .B2(new_n654), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n824), .A2(new_n825), .ZN(G1341gat));
  OAI21_X1  g625(.A(G127gat), .B1(new_n818), .B2(new_n588), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n821), .A2(new_n299), .A3(new_n589), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(G1342gat));
  NAND3_X1  g628(.A1(new_n821), .A2(new_n297), .A3(new_n695), .ZN(new_n830));
  XOR2_X1   g629(.A(new_n830), .B(KEYINPUT56), .Z(new_n831));
  OAI21_X1  g630(.A(G134gat), .B1(new_n818), .B2(new_n628), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(G1343gat));
  NOR3_X1   g632(.A1(new_n511), .A2(new_n460), .A3(new_n286), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n801), .A2(new_n794), .A3(new_n802), .ZN(new_n836));
  AOI21_X1  g635(.A(KEYINPUT115), .B1(new_n804), .B2(KEYINPUT55), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n649), .B(new_n813), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n810), .A2(new_n654), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n695), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n840), .A2(KEYINPUT116), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n812), .B1(new_n840), .B2(KEYINPUT116), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n588), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n792), .ZN(new_n844));
  AOI211_X1 g643(.A(new_n835), .B(new_n497), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n835), .B1(new_n816), .B2(new_n497), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n834), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(G141gat), .B1(new_n848), .B2(new_n565), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n695), .A2(new_n810), .A3(new_n811), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n649), .B1(new_n836), .B2(new_n837), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n588), .B1(new_n840), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n844), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n462), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n856), .A2(new_n834), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(new_n319), .A3(new_n564), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n849), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT58), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT58), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n849), .A2(new_n861), .A3(new_n858), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(new_n862), .ZN(G1344gat));
  AND2_X1   g662(.A1(new_n834), .A2(new_n654), .ZN(new_n864));
  AOI211_X1 g663(.A(new_n835), .B(new_n497), .C1(new_n853), .C2(new_n844), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n846), .B1(new_n865), .B2(KEYINPUT117), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n855), .A2(new_n867), .A3(new_n835), .ZN(new_n868));
  OAI211_X1 g667(.A(KEYINPUT118), .B(new_n864), .C1(new_n866), .C2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(G148gat), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n867), .B1(new_n855), .B2(new_n835), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n865), .A2(KEYINPUT117), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n871), .A2(new_n872), .A3(new_n846), .ZN(new_n873));
  AOI21_X1  g672(.A(KEYINPUT118), .B1(new_n873), .B2(new_n864), .ZN(new_n874));
  OAI21_X1  g673(.A(KEYINPUT59), .B1(new_n870), .B2(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n320), .A2(KEYINPUT59), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n876), .B1(new_n848), .B2(new_n655), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n856), .A2(new_n320), .A3(new_n864), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(G1345gat));
  OAI21_X1  g679(.A(G155gat), .B1(new_n848), .B2(new_n588), .ZN(new_n881));
  INV_X1    g680(.A(new_n857), .ZN(new_n882));
  OR2_X1    g681(.A1(new_n588), .A2(G155gat), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(G1346gat));
  INV_X1    g683(.A(G162gat), .ZN(new_n885));
  OR3_X1    g684(.A1(new_n848), .A2(new_n885), .A3(new_n628), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n885), .B1(new_n882), .B2(new_n628), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(G1347gat));
  NOR2_X1   g687(.A1(new_n658), .A2(new_n287), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n817), .A2(new_n422), .A3(new_n889), .ZN(new_n890));
  OR2_X1    g689(.A1(new_n890), .A2(KEYINPUT121), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(KEYINPUT121), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(G169gat), .B1(new_n893), .B2(new_n565), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n816), .A2(new_n658), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n820), .A2(new_n287), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT119), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n897), .B(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n565), .A2(G169gat), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n900), .A2(KEYINPUT120), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(KEYINPUT120), .B1(new_n900), .B2(new_n901), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n894), .B1(new_n902), .B2(new_n903), .ZN(G1348gat));
  NOR3_X1   g703(.A1(new_n893), .A2(new_n220), .A3(new_n655), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n220), .B1(new_n899), .B2(new_n655), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(KEYINPUT122), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT122), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n908), .B(new_n220), .C1(new_n899), .C2(new_n655), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n905), .B1(new_n907), .B2(new_n909), .ZN(G1349gat));
  INV_X1    g709(.A(KEYINPUT121), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n890), .B(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n228), .B1(new_n912), .B2(new_n589), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n895), .A2(new_n248), .A3(new_n589), .A4(new_n896), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(KEYINPUT123), .ZN(new_n915));
  OAI21_X1  g714(.A(KEYINPUT60), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(G183gat), .B1(new_n893), .B2(new_n588), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT60), .ZN(new_n918));
  INV_X1    g717(.A(new_n915), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n916), .A2(new_n920), .ZN(G1350gat));
  NAND3_X1  g720(.A1(new_n900), .A2(new_n230), .A3(new_n695), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n891), .A2(new_n695), .A3(new_n892), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT61), .ZN(new_n924));
  AND3_X1   g723(.A1(new_n923), .A2(new_n924), .A3(G190gat), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n924), .B1(new_n923), .B2(G190gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n922), .B1(new_n925), .B2(new_n926), .ZN(G1351gat));
  NAND3_X1  g726(.A1(new_n510), .A2(new_n286), .A3(new_n462), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT124), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n816), .A2(new_n658), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(G197gat), .B1(new_n930), .B2(new_n564), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n889), .A2(new_n510), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT125), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n873), .A2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n564), .A2(G197gat), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n931), .B1(new_n935), .B2(new_n936), .ZN(G1352gat));
  OAI21_X1  g736(.A(G204gat), .B1(new_n934), .B2(new_n655), .ZN(new_n938));
  INV_X1    g737(.A(G204gat), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n930), .A2(new_n939), .A3(new_n654), .ZN(new_n940));
  XOR2_X1   g739(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n941));
  XNOR2_X1  g740(.A(new_n940), .B(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n938), .A2(new_n942), .ZN(G1353gat));
  NAND3_X1  g742(.A1(new_n930), .A2(new_n203), .A3(new_n589), .ZN(new_n944));
  INV_X1    g743(.A(G211gat), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n932), .A2(new_n588), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n945), .B1(new_n873), .B2(new_n946), .ZN(new_n947));
  OR2_X1    g746(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n950), .B1(new_n947), .B2(new_n948), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n944), .B1(new_n949), .B2(new_n951), .ZN(G1354gat));
  AOI21_X1  g751(.A(G218gat), .B1(new_n930), .B2(new_n695), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n628), .A2(new_n204), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n953), .B1(new_n935), .B2(new_n954), .ZN(G1355gat));
endmodule


