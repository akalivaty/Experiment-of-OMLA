

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582;

  XNOR2_X1 U321 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U322 ( .A(n452), .B(KEYINPUT117), .ZN(n563) );
  XNOR2_X1 U323 ( .A(n359), .B(n358), .ZN(n360) );
  NOR2_X1 U324 ( .A1(n562), .A2(n400), .ZN(n401) );
  XNOR2_X1 U325 ( .A(n428), .B(KEYINPUT116), .ZN(n429) );
  XNOR2_X1 U326 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U327 ( .A(n404), .B(KEYINPUT41), .Z(n531) );
  XNOR2_X1 U328 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U329 ( .A(n456), .B(n455), .ZN(G1349GAT) );
  XNOR2_X1 U330 ( .A(KEYINPUT85), .B(KEYINPUT84), .ZN(n289) );
  XNOR2_X1 U331 ( .A(n289), .B(KEYINPUT3), .ZN(n290) );
  XOR2_X1 U332 ( .A(n290), .B(KEYINPUT2), .Z(n292) );
  XNOR2_X1 U333 ( .A(G141GAT), .B(G148GAT), .ZN(n291) );
  XNOR2_X1 U334 ( .A(n292), .B(n291), .ZN(n329) );
  XOR2_X1 U335 ( .A(G106GAT), .B(G162GAT), .Z(n294) );
  XNOR2_X1 U336 ( .A(G50GAT), .B(KEYINPUT69), .ZN(n293) );
  XNOR2_X1 U337 ( .A(n294), .B(n293), .ZN(n334) );
  XOR2_X1 U338 ( .A(n334), .B(KEYINPUT80), .Z(n296) );
  NAND2_X1 U339 ( .A1(G228GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U340 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U341 ( .A(n329), .B(n297), .ZN(n311) );
  XOR2_X1 U342 ( .A(KEYINPUT22), .B(G204GAT), .Z(n299) );
  XNOR2_X1 U343 ( .A(KEYINPUT86), .B(KEYINPUT81), .ZN(n298) );
  XNOR2_X1 U344 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U345 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n301) );
  XNOR2_X1 U346 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n300) );
  XNOR2_X1 U347 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U348 ( .A(G197GAT), .B(n302), .Z(n416) );
  XOR2_X1 U349 ( .A(n303), .B(n416), .Z(n309) );
  XOR2_X1 U350 ( .A(KEYINPUT23), .B(G218GAT), .Z(n306) );
  XNOR2_X1 U351 ( .A(G22GAT), .B(G155GAT), .ZN(n304) );
  XNOR2_X1 U352 ( .A(n304), .B(G78GAT), .ZN(n382) );
  XNOR2_X1 U353 ( .A(KEYINPUT87), .B(n382), .ZN(n305) );
  XNOR2_X1 U354 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U355 ( .A(KEYINPUT24), .B(n307), .ZN(n308) );
  XNOR2_X1 U356 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U357 ( .A(n311), .B(n310), .ZN(n467) );
  XOR2_X1 U358 ( .A(G120GAT), .B(G57GAT), .Z(n348) );
  XOR2_X1 U359 ( .A(G1GAT), .B(G127GAT), .Z(n386) );
  XOR2_X1 U360 ( .A(n348), .B(n386), .Z(n313) );
  XNOR2_X1 U361 ( .A(G162GAT), .B(G155GAT), .ZN(n312) );
  XNOR2_X1 U362 ( .A(n313), .B(n312), .ZN(n325) );
  XOR2_X1 U363 ( .A(KEYINPUT90), .B(KEYINPUT4), .Z(n315) );
  XNOR2_X1 U364 ( .A(KEYINPUT88), .B(KEYINPUT5), .ZN(n314) );
  XNOR2_X1 U365 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U366 ( .A(KEYINPUT91), .B(KEYINPUT6), .Z(n317) );
  XNOR2_X1 U367 ( .A(KEYINPUT1), .B(KEYINPUT89), .ZN(n316) );
  XNOR2_X1 U368 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U369 ( .A(n319), .B(n318), .Z(n323) );
  XNOR2_X1 U370 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n320) );
  XNOR2_X1 U371 ( .A(n320), .B(KEYINPUT75), .ZN(n441) );
  XNOR2_X1 U372 ( .A(G29GAT), .B(G134GAT), .ZN(n321) );
  XNOR2_X1 U373 ( .A(n321), .B(G85GAT), .ZN(n342) );
  XNOR2_X1 U374 ( .A(n441), .B(n342), .ZN(n322) );
  XNOR2_X1 U375 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U376 ( .A(n325), .B(n324), .Z(n327) );
  NAND2_X1 U377 ( .A1(G225GAT), .A2(G233GAT), .ZN(n326) );
  XNOR2_X1 U378 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U379 ( .A(n329), .B(n328), .ZN(n464) );
  XNOR2_X1 U380 ( .A(KEYINPUT92), .B(n464), .ZN(n489) );
  XOR2_X1 U381 ( .A(KEYINPUT64), .B(KEYINPUT11), .Z(n331) );
  NAND2_X1 U382 ( .A1(G232GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U383 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U384 ( .A(n332), .B(KEYINPUT10), .Z(n336) );
  XNOR2_X1 U385 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n333) );
  XNOR2_X1 U386 ( .A(n333), .B(KEYINPUT7), .ZN(n363) );
  XNOR2_X1 U387 ( .A(n363), .B(n334), .ZN(n335) );
  XNOR2_X1 U388 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U389 ( .A(G92GAT), .B(KEYINPUT9), .Z(n338) );
  XNOR2_X1 U390 ( .A(G99GAT), .B(KEYINPUT70), .ZN(n337) );
  XNOR2_X1 U391 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U392 ( .A(n340), .B(n339), .Z(n344) );
  XNOR2_X1 U393 ( .A(G36GAT), .B(G190GAT), .ZN(n341) );
  XNOR2_X1 U394 ( .A(n341), .B(G218GAT), .ZN(n422) );
  XNOR2_X1 U395 ( .A(n342), .B(n422), .ZN(n343) );
  XNOR2_X1 U396 ( .A(n344), .B(n343), .ZN(n562) );
  XOR2_X1 U397 ( .A(G78GAT), .B(KEYINPUT31), .Z(n346) );
  XNOR2_X1 U398 ( .A(G99GAT), .B(G148GAT), .ZN(n345) );
  XNOR2_X1 U399 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U400 ( .A(n348), .B(n347), .ZN(n350) );
  AND2_X1 U401 ( .A1(G230GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U402 ( .A(n350), .B(n349), .ZN(n352) );
  INV_X1 U403 ( .A(KEYINPUT33), .ZN(n351) );
  XNOR2_X1 U404 ( .A(n352), .B(n351), .ZN(n359) );
  XOR2_X1 U405 ( .A(G64GAT), .B(G92GAT), .Z(n354) );
  XNOR2_X1 U406 ( .A(G176GAT), .B(G204GAT), .ZN(n353) );
  XNOR2_X1 U407 ( .A(n354), .B(n353), .ZN(n419) );
  XNOR2_X1 U408 ( .A(n419), .B(KEYINPUT32), .ZN(n357) );
  XNOR2_X1 U409 ( .A(G106GAT), .B(G85GAT), .ZN(n355) );
  XNOR2_X1 U410 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n385) );
  XNOR2_X1 U411 ( .A(n355), .B(n385), .ZN(n356) );
  INV_X1 U412 ( .A(n360), .ZN(n404) );
  INV_X1 U413 ( .A(n531), .ZN(n503) );
  XOR2_X1 U414 ( .A(G29GAT), .B(G36GAT), .Z(n362) );
  XNOR2_X1 U415 ( .A(G50GAT), .B(G197GAT), .ZN(n361) );
  XNOR2_X1 U416 ( .A(n362), .B(n361), .ZN(n364) );
  XOR2_X1 U417 ( .A(n364), .B(n363), .Z(n369) );
  XOR2_X1 U418 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n366) );
  NAND2_X1 U419 ( .A1(G229GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U420 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U421 ( .A(KEYINPUT30), .B(n367), .ZN(n368) );
  XNOR2_X1 U422 ( .A(n369), .B(n368), .ZN(n377) );
  XOR2_X1 U423 ( .A(G15GAT), .B(G22GAT), .Z(n371) );
  XNOR2_X1 U424 ( .A(G169GAT), .B(G141GAT), .ZN(n370) );
  XNOR2_X1 U425 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U426 ( .A(KEYINPUT68), .B(G8GAT), .Z(n373) );
  XNOR2_X1 U427 ( .A(G113GAT), .B(G1GAT), .ZN(n372) );
  XNOR2_X1 U428 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U429 ( .A(n375), .B(n374), .Z(n376) );
  XNOR2_X1 U430 ( .A(n377), .B(n376), .ZN(n554) );
  INV_X1 U431 ( .A(n554), .ZN(n568) );
  NOR2_X1 U432 ( .A1(n503), .A2(n568), .ZN(n378) );
  XNOR2_X1 U433 ( .A(n378), .B(KEYINPUT46), .ZN(n398) );
  XOR2_X1 U434 ( .A(G64GAT), .B(KEYINPUT73), .Z(n380) );
  XNOR2_X1 U435 ( .A(G57GAT), .B(KEYINPUT15), .ZN(n379) );
  XNOR2_X1 U436 ( .A(n380), .B(n379), .ZN(n397) );
  XNOR2_X1 U437 ( .A(G8GAT), .B(G183GAT), .ZN(n381) );
  XNOR2_X1 U438 ( .A(n381), .B(KEYINPUT71), .ZN(n421) );
  XNOR2_X1 U439 ( .A(n382), .B(n421), .ZN(n395) );
  XOR2_X1 U440 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n384) );
  XNOR2_X1 U441 ( .A(KEYINPUT72), .B(KEYINPUT74), .ZN(n383) );
  XNOR2_X1 U442 ( .A(n384), .B(n383), .ZN(n391) );
  INV_X1 U443 ( .A(n385), .ZN(n387) );
  XOR2_X1 U444 ( .A(n387), .B(n386), .Z(n389) );
  XNOR2_X1 U445 ( .A(G15GAT), .B(G211GAT), .ZN(n388) );
  XNOR2_X1 U446 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U447 ( .A(n391), .B(n390), .Z(n393) );
  NAND2_X1 U448 ( .A1(G231GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U449 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U450 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U451 ( .A(n397), .B(n396), .ZN(n402) );
  INV_X1 U452 ( .A(n402), .ZN(n548) );
  XNOR2_X1 U453 ( .A(KEYINPUT106), .B(n548), .ZN(n558) );
  NOR2_X1 U454 ( .A1(n398), .A2(n558), .ZN(n399) );
  XNOR2_X1 U455 ( .A(n399), .B(KEYINPUT107), .ZN(n400) );
  XNOR2_X1 U456 ( .A(n401), .B(KEYINPUT47), .ZN(n409) );
  XOR2_X1 U457 ( .A(n562), .B(KEYINPUT36), .Z(n580) );
  NOR2_X1 U458 ( .A1(n580), .A2(n402), .ZN(n403) );
  XNOR2_X1 U459 ( .A(KEYINPUT45), .B(n403), .ZN(n405) );
  NAND2_X1 U460 ( .A1(n405), .A2(n360), .ZN(n406) );
  NOR2_X1 U461 ( .A1(n554), .A2(n406), .ZN(n407) );
  XOR2_X1 U462 ( .A(KEYINPUT108), .B(n407), .Z(n408) );
  NAND2_X1 U463 ( .A1(n409), .A2(n408), .ZN(n411) );
  XNOR2_X1 U464 ( .A(KEYINPUT48), .B(KEYINPUT109), .ZN(n410) );
  XNOR2_X1 U465 ( .A(n411), .B(n410), .ZN(n526) );
  XNOR2_X1 U466 ( .A(KEYINPUT78), .B(KEYINPUT19), .ZN(n412) );
  XNOR2_X1 U467 ( .A(n412), .B(KEYINPUT17), .ZN(n413) );
  XOR2_X1 U468 ( .A(n413), .B(KEYINPUT77), .Z(n415) );
  XNOR2_X1 U469 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n414) );
  XOR2_X1 U470 ( .A(n415), .B(n414), .Z(n449) );
  XOR2_X1 U471 ( .A(n449), .B(n416), .Z(n426) );
  XOR2_X1 U472 ( .A(KEYINPUT94), .B(KEYINPUT93), .Z(n418) );
  NAND2_X1 U473 ( .A1(G226GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U474 ( .A(n418), .B(n417), .ZN(n420) );
  XOR2_X1 U475 ( .A(n420), .B(n419), .Z(n424) );
  XNOR2_X1 U476 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U477 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U478 ( .A(n426), .B(n425), .ZN(n493) );
  XNOR2_X1 U479 ( .A(n493), .B(KEYINPUT115), .ZN(n427) );
  NOR2_X1 U480 ( .A1(n526), .A2(n427), .ZN(n430) );
  INV_X1 U481 ( .A(KEYINPUT54), .ZN(n428) );
  NOR2_X1 U482 ( .A1(n489), .A2(n431), .ZN(n567) );
  NAND2_X1 U483 ( .A1(n467), .A2(n567), .ZN(n432) );
  XNOR2_X1 U484 ( .A(n432), .B(KEYINPUT55), .ZN(n451) );
  XOR2_X1 U485 ( .A(G127GAT), .B(G176GAT), .Z(n434) );
  XNOR2_X1 U486 ( .A(G15GAT), .B(G183GAT), .ZN(n433) );
  XNOR2_X1 U487 ( .A(n434), .B(n433), .ZN(n448) );
  XOR2_X1 U488 ( .A(KEYINPUT65), .B(G71GAT), .Z(n436) );
  XNOR2_X1 U489 ( .A(G43GAT), .B(G99GAT), .ZN(n435) );
  XNOR2_X1 U490 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U491 ( .A(KEYINPUT76), .B(KEYINPUT20), .Z(n438) );
  XNOR2_X1 U492 ( .A(KEYINPUT79), .B(G120GAT), .ZN(n437) );
  XNOR2_X1 U493 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U494 ( .A(n440), .B(n439), .Z(n446) );
  XOR2_X1 U495 ( .A(G134GAT), .B(n441), .Z(n443) );
  NAND2_X1 U496 ( .A1(G227GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U498 ( .A(G190GAT), .B(n444), .ZN(n445) );
  XNOR2_X1 U499 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U500 ( .A(n448), .B(n447), .ZN(n450) );
  XNOR2_X1 U501 ( .A(n450), .B(n449), .ZN(n495) );
  NAND2_X1 U502 ( .A1(n451), .A2(n495), .ZN(n452) );
  NAND2_X1 U503 ( .A1(n563), .A2(n531), .ZN(n456) );
  XOR2_X1 U504 ( .A(G176GAT), .B(KEYINPUT56), .Z(n454) );
  XNOR2_X1 U505 ( .A(KEYINPUT57), .B(KEYINPUT120), .ZN(n453) );
  INV_X1 U506 ( .A(n489), .ZN(n516) );
  NOR2_X1 U507 ( .A1(n568), .A2(n404), .ZN(n486) );
  NAND2_X1 U508 ( .A1(n493), .A2(n495), .ZN(n457) );
  NAND2_X1 U509 ( .A1(n467), .A2(n457), .ZN(n458) );
  XNOR2_X1 U510 ( .A(KEYINPUT25), .B(n458), .ZN(n463) );
  NOR2_X1 U511 ( .A1(n495), .A2(n467), .ZN(n459) );
  XNOR2_X1 U512 ( .A(n459), .B(KEYINPUT26), .ZN(n566) );
  XOR2_X1 U513 ( .A(n493), .B(KEYINPUT27), .Z(n460) );
  XNOR2_X1 U514 ( .A(KEYINPUT95), .B(n460), .ZN(n466) );
  NAND2_X1 U515 ( .A1(n566), .A2(n466), .ZN(n461) );
  XOR2_X1 U516 ( .A(KEYINPUT96), .B(n461), .Z(n462) );
  NOR2_X1 U517 ( .A1(n463), .A2(n462), .ZN(n465) );
  NOR2_X1 U518 ( .A1(n465), .A2(n464), .ZN(n471) );
  NAND2_X1 U519 ( .A1(n466), .A2(n489), .ZN(n525) );
  XNOR2_X1 U520 ( .A(n467), .B(KEYINPUT66), .ZN(n468) );
  XNOR2_X1 U521 ( .A(n468), .B(KEYINPUT28), .ZN(n527) );
  INV_X1 U522 ( .A(n527), .ZN(n501) );
  OR2_X1 U523 ( .A1(n525), .A2(n501), .ZN(n469) );
  NOR2_X1 U524 ( .A1(n469), .A2(n495), .ZN(n470) );
  NOR2_X1 U525 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X1 U526 ( .A(KEYINPUT97), .B(n472), .ZN(n484) );
  INV_X1 U527 ( .A(n562), .ZN(n552) );
  NAND2_X1 U528 ( .A1(n548), .A2(n552), .ZN(n473) );
  XOR2_X1 U529 ( .A(KEYINPUT16), .B(n473), .Z(n474) );
  AND2_X1 U530 ( .A1(n484), .A2(n474), .ZN(n504) );
  NAND2_X1 U531 ( .A1(n486), .A2(n504), .ZN(n481) );
  NOR2_X1 U532 ( .A1(n516), .A2(n481), .ZN(n475) );
  XOR2_X1 U533 ( .A(KEYINPUT34), .B(n475), .Z(n476) );
  XNOR2_X1 U534 ( .A(G1GAT), .B(n476), .ZN(G1324GAT) );
  INV_X1 U535 ( .A(n493), .ZN(n519) );
  NOR2_X1 U536 ( .A1(n519), .A2(n481), .ZN(n477) );
  XOR2_X1 U537 ( .A(G8GAT), .B(n477), .Z(G1325GAT) );
  INV_X1 U538 ( .A(n495), .ZN(n529) );
  NOR2_X1 U539 ( .A1(n529), .A2(n481), .ZN(n479) );
  XNOR2_X1 U540 ( .A(KEYINPUT98), .B(KEYINPUT35), .ZN(n478) );
  XNOR2_X1 U541 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U542 ( .A(G15GAT), .B(n480), .ZN(G1326GAT) );
  NOR2_X1 U543 ( .A1(n527), .A2(n481), .ZN(n482) );
  XOR2_X1 U544 ( .A(G22GAT), .B(n482), .Z(G1327GAT) );
  XOR2_X1 U545 ( .A(G29GAT), .B(KEYINPUT100), .Z(n491) );
  NOR2_X1 U546 ( .A1(n548), .A2(n580), .ZN(n483) );
  NAND2_X1 U547 ( .A1(n484), .A2(n483), .ZN(n485) );
  XNOR2_X1 U548 ( .A(KEYINPUT37), .B(n485), .ZN(n513) );
  NAND2_X1 U549 ( .A1(n486), .A2(n513), .ZN(n487) );
  XNOR2_X1 U550 ( .A(n487), .B(KEYINPUT99), .ZN(n488) );
  XNOR2_X1 U551 ( .A(KEYINPUT38), .B(n488), .ZN(n500) );
  NAND2_X1 U552 ( .A1(n489), .A2(n500), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U554 ( .A(KEYINPUT39), .B(n492), .ZN(G1328GAT) );
  NAND2_X1 U555 ( .A1(n500), .A2(n493), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n494), .B(G36GAT), .ZN(G1329GAT) );
  XNOR2_X1 U557 ( .A(G43GAT), .B(KEYINPUT102), .ZN(n499) );
  XOR2_X1 U558 ( .A(KEYINPUT101), .B(KEYINPUT40), .Z(n497) );
  NAND2_X1 U559 ( .A1(n500), .A2(n495), .ZN(n496) );
  XNOR2_X1 U560 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U561 ( .A(n499), .B(n498), .ZN(G1330GAT) );
  NAND2_X1 U562 ( .A1(n501), .A2(n500), .ZN(n502) );
  XNOR2_X1 U563 ( .A(G50GAT), .B(n502), .ZN(G1331GAT) );
  NOR2_X1 U564 ( .A1(n503), .A2(n554), .ZN(n514) );
  NAND2_X1 U565 ( .A1(n514), .A2(n504), .ZN(n510) );
  NOR2_X1 U566 ( .A1(n516), .A2(n510), .ZN(n505) );
  XOR2_X1 U567 ( .A(G57GAT), .B(n505), .Z(n506) );
  XNOR2_X1 U568 ( .A(KEYINPUT42), .B(n506), .ZN(G1332GAT) );
  NOR2_X1 U569 ( .A1(n519), .A2(n510), .ZN(n507) );
  XOR2_X1 U570 ( .A(G64GAT), .B(n507), .Z(G1333GAT) );
  NOR2_X1 U571 ( .A1(n529), .A2(n510), .ZN(n509) );
  XNOR2_X1 U572 ( .A(G71GAT), .B(KEYINPUT103), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n509), .B(n508), .ZN(G1334GAT) );
  NOR2_X1 U574 ( .A1(n527), .A2(n510), .ZN(n512) );
  XNOR2_X1 U575 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n511) );
  XNOR2_X1 U576 ( .A(n512), .B(n511), .ZN(G1335GAT) );
  NAND2_X1 U577 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X1 U578 ( .A(n515), .B(KEYINPUT104), .ZN(n522) );
  NOR2_X1 U579 ( .A1(n522), .A2(n516), .ZN(n518) );
  XNOR2_X1 U580 ( .A(G85GAT), .B(KEYINPUT105), .ZN(n517) );
  XNOR2_X1 U581 ( .A(n518), .B(n517), .ZN(G1336GAT) );
  NOR2_X1 U582 ( .A1(n522), .A2(n519), .ZN(n520) );
  XOR2_X1 U583 ( .A(G92GAT), .B(n520), .Z(G1337GAT) );
  NOR2_X1 U584 ( .A1(n529), .A2(n522), .ZN(n521) );
  XOR2_X1 U585 ( .A(G99GAT), .B(n521), .Z(G1338GAT) );
  NOR2_X1 U586 ( .A1(n527), .A2(n522), .ZN(n523) );
  XOR2_X1 U587 ( .A(KEYINPUT44), .B(n523), .Z(n524) );
  XNOR2_X1 U588 ( .A(G106GAT), .B(n524), .ZN(G1339GAT) );
  NOR2_X1 U589 ( .A1(n526), .A2(n525), .ZN(n543) );
  NAND2_X1 U590 ( .A1(n527), .A2(n543), .ZN(n528) );
  NOR2_X1 U591 ( .A1(n529), .A2(n528), .ZN(n540) );
  NAND2_X1 U592 ( .A1(n540), .A2(n554), .ZN(n530) );
  XNOR2_X1 U593 ( .A(G113GAT), .B(n530), .ZN(G1340GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT49), .B(KEYINPUT110), .Z(n533) );
  NAND2_X1 U595 ( .A1(n540), .A2(n531), .ZN(n532) );
  XNOR2_X1 U596 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U597 ( .A(G120GAT), .B(n534), .ZN(G1341GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT50), .B(KEYINPUT113), .Z(n536) );
  XNOR2_X1 U599 ( .A(G127GAT), .B(KEYINPUT112), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U601 ( .A(KEYINPUT111), .B(n537), .Z(n539) );
  NAND2_X1 U602 ( .A1(n540), .A2(n558), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(G1342GAT) );
  XOR2_X1 U604 ( .A(G134GAT), .B(KEYINPUT51), .Z(n542) );
  NAND2_X1 U605 ( .A1(n540), .A2(n562), .ZN(n541) );
  XNOR2_X1 U606 ( .A(n542), .B(n541), .ZN(G1343GAT) );
  NAND2_X1 U607 ( .A1(n543), .A2(n566), .ZN(n551) );
  NOR2_X1 U608 ( .A1(n568), .A2(n551), .ZN(n544) );
  XOR2_X1 U609 ( .A(G141GAT), .B(n544), .Z(G1344GAT) );
  NOR2_X1 U610 ( .A1(n503), .A2(n551), .ZN(n546) );
  XNOR2_X1 U611 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(n547), .ZN(G1345GAT) );
  NOR2_X1 U614 ( .A1(n402), .A2(n551), .ZN(n549) );
  XOR2_X1 U615 ( .A(KEYINPUT114), .B(n549), .Z(n550) );
  XNOR2_X1 U616 ( .A(G155GAT), .B(n550), .ZN(G1346GAT) );
  NOR2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U618 ( .A(G162GAT), .B(n553), .Z(G1347GAT) );
  NAND2_X1 U619 ( .A1(n554), .A2(n563), .ZN(n557) );
  XOR2_X1 U620 ( .A(G169GAT), .B(KEYINPUT118), .Z(n555) );
  XNOR2_X1 U621 ( .A(KEYINPUT119), .B(n555), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(G1348GAT) );
  NAND2_X1 U623 ( .A1(n563), .A2(n558), .ZN(n560) );
  XOR2_X1 U624 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n559) );
  XNOR2_X1 U625 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U626 ( .A(n561), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U627 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U628 ( .A(n564), .B(KEYINPUT58), .ZN(n565) );
  XNOR2_X1 U629 ( .A(n565), .B(G190GAT), .ZN(G1351GAT) );
  NAND2_X1 U630 ( .A1(n567), .A2(n566), .ZN(n579) );
  NOR2_X1 U631 ( .A1(n579), .A2(n568), .ZN(n572) );
  XOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n570) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n569) );
  XNOR2_X1 U634 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U635 ( .A(n572), .B(n571), .ZN(G1352GAT) );
  NOR2_X1 U636 ( .A1(n579), .A2(n360), .ZN(n576) );
  XOR2_X1 U637 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n574) );
  XNOR2_X1 U638 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n576), .B(n575), .ZN(G1353GAT) );
  NOR2_X1 U641 ( .A1(n402), .A2(n579), .ZN(n577) );
  XOR2_X1 U642 ( .A(KEYINPUT126), .B(n577), .Z(n578) );
  XNOR2_X1 U643 ( .A(G211GAT), .B(n578), .ZN(G1354GAT) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U645 ( .A(KEYINPUT62), .B(n581), .Z(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

