//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 0 0 1 1 1 1 0 0 1 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 1 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G29gat), .A2(G36gat), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT14), .ZN(new_n208));
  INV_X1    g007(.A(G29gat), .ZN(new_n209));
  INV_X1    g008(.A(G36gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT92), .ZN(new_n212));
  NOR2_X1   g011(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT92), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n213), .A2(new_n214), .A3(new_n210), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n207), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n205), .B1(new_n216), .B2(KEYINPUT93), .ZN(new_n217));
  NOR4_X1   g016(.A1(KEYINPUT92), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n214), .B1(new_n213), .B2(new_n210), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n206), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT93), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n204), .B1(new_n217), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n211), .A2(new_n206), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(KEYINPUT15), .B2(new_n202), .ZN(new_n225));
  INV_X1    g024(.A(new_n205), .ZN(new_n226));
  NOR3_X1   g025(.A1(new_n225), .A2(new_n204), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n223), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G8gat), .ZN(new_n230));
  XNOR2_X1  g029(.A(G15gat), .B(G22gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n231), .A2(G1gat), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n230), .B1(new_n232), .B2(KEYINPUT94), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT16), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n231), .B1(new_n234), .B2(G1gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n235), .B1(G1gat), .B2(new_n231), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n233), .B(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n229), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(G229gat), .A2(G233gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT18), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT95), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n226), .B1(new_n220), .B2(new_n221), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n216), .A2(KEYINPUT93), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n203), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(KEYINPUT17), .B1(new_n246), .B2(new_n227), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT17), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n223), .A2(new_n248), .A3(new_n228), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n237), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n243), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  AOI211_X1 g051(.A(KEYINPUT95), .B(new_n237), .C1(new_n247), .C2(new_n249), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n242), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT96), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n242), .B(KEYINPUT96), .C1(new_n252), .C2(new_n253), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G113gat), .B(G141gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(G197gat), .ZN(new_n260));
  XOR2_X1   g059(.A(KEYINPUT11), .B(G169gat), .Z(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(new_n262), .B(KEYINPUT12), .Z(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n251), .B(new_n229), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n239), .B(KEYINPUT13), .Z(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n238), .B(new_n239), .C1(new_n252), .C2(new_n253), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n268), .B1(new_n269), .B2(new_n241), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n258), .A2(new_n264), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n264), .B1(new_n258), .B2(new_n270), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(G211gat), .A2(G218gat), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT22), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(G197gat), .ZN(new_n277));
  INV_X1    g076(.A(G204gat), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g078(.A1(G197gat), .A2(G204gat), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n276), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G211gat), .B(G218gat), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  OR3_X1    g083(.A1(new_n282), .A2(KEYINPUT76), .A3(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n284), .B1(new_n282), .B2(KEYINPUT76), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT78), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT29), .ZN(new_n289));
  NOR2_X1   g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290));
  AND2_X1   g089(.A1(KEYINPUT69), .A2(KEYINPUT26), .ZN(new_n291));
  NOR2_X1   g090(.A1(KEYINPUT69), .A2(KEYINPUT26), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n293), .B(KEYINPUT70), .ZN(new_n294));
  NAND2_X1  g093(.A1(G169gat), .A2(G176gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT26), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n295), .B1(new_n290), .B2(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G183gat), .ZN(new_n299));
  INV_X1    g098(.A(G190gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT68), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT27), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n302), .B1(new_n303), .B2(G183gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(KEYINPUT27), .B(G183gat), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n300), .B(new_n304), .C1(new_n305), .C2(new_n302), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT28), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n307), .A2(G190gat), .ZN(new_n308));
  AOI22_X1  g107(.A1(new_n306), .A2(new_n307), .B1(new_n305), .B2(new_n308), .ZN(new_n309));
  NOR3_X1   g108(.A1(new_n298), .A2(new_n301), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G169gat), .ZN(new_n312));
  INV_X1    g111(.A(G176gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT23), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n295), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n316), .B(KEYINPUT65), .ZN(new_n317));
  NOR3_X1   g116(.A1(new_n299), .A2(new_n300), .A3(KEYINPUT24), .ZN(new_n318));
  XOR2_X1   g117(.A(G183gat), .B(G190gat), .Z(new_n319));
  AOI21_X1  g118(.A(new_n318), .B1(new_n319), .B2(KEYINPUT24), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n314), .A2(new_n315), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n317), .A2(KEYINPUT25), .A3(new_n320), .A4(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT66), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AND3_X1   g123(.A1(new_n320), .A2(KEYINPUT25), .A3(new_n321), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n325), .A2(KEYINPUT66), .A3(new_n317), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT25), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n290), .A2(KEYINPUT23), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n321), .A2(new_n295), .A3(new_n328), .ZN(new_n329));
  OR2_X1    g128(.A1(new_n329), .A2(KEYINPUT64), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(KEYINPUT64), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n330), .A2(new_n320), .A3(new_n331), .ZN(new_n332));
  AOI22_X1  g131(.A1(new_n324), .A2(new_n326), .B1(new_n327), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n311), .B1(new_n333), .B2(KEYINPUT67), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n332), .A2(new_n327), .ZN(new_n335));
  INV_X1    g134(.A(new_n326), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT66), .B1(new_n325), .B2(new_n317), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n335), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT67), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n289), .B1(new_n334), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(G226gat), .A2(G233gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n342), .B(KEYINPUT77), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n333), .A2(new_n310), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n346), .A2(new_n344), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n288), .B1(new_n345), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(KEYINPUT78), .B1(new_n341), .B2(new_n344), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n287), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n338), .A2(new_n339), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n333), .A2(KEYINPUT67), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n352), .A2(new_n353), .A3(new_n311), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(new_n343), .ZN(new_n355));
  INV_X1    g154(.A(new_n287), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n344), .B1(new_n346), .B2(KEYINPUT29), .ZN(new_n357));
  AND3_X1   g156(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  XOR2_X1   g158(.A(G8gat), .B(G36gat), .Z(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(KEYINPUT79), .ZN(new_n361));
  XNOR2_X1  g160(.A(G64gat), .B(G92gat), .ZN(new_n362));
  XOR2_X1   g161(.A(new_n361), .B(new_n362), .Z(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n351), .A2(KEYINPUT30), .A3(new_n359), .A4(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n343), .B1(new_n354), .B2(new_n289), .ZN(new_n366));
  OAI21_X1  g165(.A(KEYINPUT78), .B1(new_n366), .B2(new_n347), .ZN(new_n367));
  INV_X1    g166(.A(new_n350), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n356), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n363), .B1(new_n369), .B2(new_n358), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n365), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT80), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  XOR2_X1   g172(.A(G1gat), .B(G29gat), .Z(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT85), .B(KEYINPUT0), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(G57gat), .B(G85gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n376), .B(new_n377), .ZN(new_n378));
  XOR2_X1   g177(.A(G113gat), .B(G120gat), .Z(new_n379));
  NOR2_X1   g178(.A1(KEYINPUT71), .A2(KEYINPUT1), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(G127gat), .B(G134gat), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n381), .B(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(G155gat), .ZN(new_n385));
  INV_X1    g184(.A(G162gat), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT2), .ZN(new_n388));
  NOR2_X1   g187(.A1(G155gat), .A2(G162gat), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  XOR2_X1   g189(.A(KEYINPUT82), .B(G141gat), .Z(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(G148gat), .ZN(new_n392));
  INV_X1    g191(.A(G148gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(G141gat), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n390), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  XOR2_X1   g194(.A(G141gat), .B(G148gat), .Z(new_n396));
  XOR2_X1   g195(.A(KEYINPUT81), .B(KEYINPUT2), .Z(new_n397));
  AOI211_X1 g196(.A(new_n387), .B(new_n389), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n384), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n398), .A2(new_n395), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n381), .B(new_n382), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(G225gat), .A2(G233gat), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT84), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n406), .A2(new_n407), .A3(KEYINPUT5), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n404), .B1(new_n399), .B2(new_n402), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT5), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT84), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT3), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n400), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(KEYINPUT3), .B1(new_n398), .B2(new_n395), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n413), .A2(new_n414), .A3(new_n384), .ZN(new_n415));
  AND2_X1   g214(.A1(new_n415), .A2(new_n404), .ZN(new_n416));
  XOR2_X1   g215(.A(KEYINPUT83), .B(KEYINPUT4), .Z(new_n417));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n400), .A2(new_n401), .A3(KEYINPUT4), .ZN(new_n419));
  AND2_X1   g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n408), .A2(new_n411), .B1(new_n416), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT4), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n402), .A2(new_n422), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n423), .B(new_n410), .C1(new_n402), .C2(new_n417), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n415), .A2(new_n404), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n378), .B1(new_n421), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT87), .ZN(new_n428));
  OR2_X1    g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n427), .A2(new_n428), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n416), .A2(new_n420), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n407), .B1(new_n406), .B2(KEYINPUT5), .ZN(new_n432));
  NOR3_X1   g231(.A1(new_n409), .A2(KEYINPUT84), .A3(new_n410), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n431), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n378), .ZN(new_n435));
  INV_X1    g234(.A(new_n426), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT6), .ZN(new_n438));
  AND3_X1   g237(.A1(new_n437), .A2(KEYINPUT86), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT86), .B1(new_n437), .B2(new_n438), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n429), .B(new_n430), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT88), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n427), .B(KEYINPUT87), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n444), .B(KEYINPUT88), .C1(new_n440), .C2(new_n439), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n427), .A2(new_n438), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n443), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n367), .A2(new_n368), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n358), .B1(new_n449), .B2(new_n287), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT30), .B1(new_n450), .B2(new_n364), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n365), .A2(new_n370), .A3(KEYINPUT80), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n373), .A2(new_n448), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(G22gat), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT89), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT29), .B1(new_n400), .B2(new_n412), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n282), .A2(new_n284), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT29), .B1(new_n281), .B2(new_n283), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT3), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OAI22_X1  g259(.A1(new_n457), .A2(new_n356), .B1(new_n400), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(G228gat), .A2(G233gat), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n456), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n461), .A2(new_n456), .A3(new_n462), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n457), .A2(new_n356), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n285), .A2(new_n289), .A3(new_n286), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n400), .B1(new_n468), .B2(new_n412), .ZN(new_n469));
  NOR3_X1   g268(.A1(new_n467), .A2(new_n462), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n455), .B1(new_n466), .B2(new_n471), .ZN(new_n472));
  AOI211_X1 g271(.A(G22gat), .B(new_n470), .C1(new_n464), .C2(new_n465), .ZN(new_n473));
  OAI21_X1  g272(.A(G78gat), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n465), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n471), .B1(new_n475), .B2(new_n463), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(G22gat), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n466), .A2(new_n455), .A3(new_n471), .ZN(new_n478));
  INV_X1    g277(.A(G78gat), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(KEYINPUT31), .B(G50gat), .ZN(new_n481));
  INV_X1    g280(.A(G106gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n481), .B(new_n482), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n474), .A2(new_n480), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n483), .B1(new_n474), .B2(new_n480), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n384), .B1(new_n334), .B2(new_n340), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n352), .A2(new_n353), .A3(new_n311), .A4(new_n401), .ZN(new_n488));
  NAND2_X1  g287(.A1(G227gat), .A2(G233gat), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT73), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n490), .A2(new_n491), .A3(KEYINPUT34), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n491), .B1(new_n490), .B2(KEYINPUT34), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT34), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n487), .A2(new_n488), .A3(new_n496), .A4(new_n489), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT74), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n497), .B(new_n498), .ZN(new_n499));
  XOR2_X1   g298(.A(G15gat), .B(G43gat), .Z(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(KEYINPUT72), .ZN(new_n501));
  XNOR2_X1  g300(.A(G71gat), .B(G99gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n489), .B1(new_n487), .B2(new_n488), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n503), .B1(new_n504), .B2(KEYINPUT33), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT32), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n487), .A2(new_n488), .ZN(new_n509));
  INV_X1    g308(.A(new_n489), .ZN(new_n510));
  AOI221_X4 g309(.A(new_n506), .B1(KEYINPUT33), .B2(new_n503), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  OAI22_X1  g310(.A1(new_n495), .A2(new_n499), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n509), .A2(new_n510), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT32), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT33), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n514), .A2(new_n516), .A3(new_n503), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n490), .A2(KEYINPUT34), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT73), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(new_n492), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n497), .B(KEYINPUT74), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n507), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n517), .A2(new_n520), .A3(new_n521), .A4(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n486), .A2(new_n512), .A3(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT35), .B1(new_n454), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n427), .A2(new_n437), .A3(new_n438), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT35), .B1(new_n447), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n486), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT75), .ZN(new_n529));
  OAI221_X1 g328(.A(new_n529), .B1(new_n508), .B2(new_n511), .C1(new_n495), .C2(new_n499), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n512), .A2(new_n523), .A3(KEYINPUT75), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n371), .A2(new_n451), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n525), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n486), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n454), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT36), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n538), .B1(new_n512), .B2(new_n523), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n531), .A2(new_n530), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n539), .B1(new_n540), .B2(new_n538), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n415), .B(new_n423), .C1(new_n402), .C2(new_n417), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n405), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(KEYINPUT90), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT39), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n378), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT90), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n543), .B(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT39), .B1(new_n403), .B2(new_n405), .ZN(new_n549));
  XOR2_X1   g348(.A(new_n549), .B(KEYINPUT91), .Z(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n546), .A2(KEYINPUT40), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n427), .ZN(new_n553));
  AOI21_X1  g352(.A(KEYINPUT40), .B1(new_n546), .B2(new_n551), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(new_n371), .B2(new_n451), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT38), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT37), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n364), .B1(new_n450), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g358(.A(KEYINPUT37), .B1(new_n369), .B2(new_n358), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n557), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n351), .A2(new_n558), .A3(new_n359), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n355), .A2(new_n357), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n558), .B1(new_n563), .B2(new_n287), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n345), .A2(new_n348), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n350), .B1(new_n565), .B2(KEYINPUT78), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n564), .B1(new_n566), .B2(new_n287), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n562), .A2(new_n567), .A3(new_n557), .A4(new_n363), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n447), .A2(new_n526), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n569), .B1(new_n450), .B2(new_n364), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n556), .B(new_n486), .C1(new_n561), .C2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n537), .A2(new_n541), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n273), .B1(new_n535), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n448), .ZN(new_n575));
  XOR2_X1   g374(.A(G57gat), .B(G64gat), .Z(new_n576));
  INV_X1    g375(.A(KEYINPUT97), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT9), .ZN(new_n578));
  INV_X1    g377(.A(G71gat), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n578), .B1(new_n579), .B2(new_n479), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n576), .A2(new_n577), .A3(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G71gat), .B(G78gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n583), .A2(KEYINPUT21), .ZN(new_n584));
  AND2_X1   g383(.A1(G231gat), .A2(G233gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(G127gat), .B(G155gat), .Z(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT20), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n586), .B(new_n588), .ZN(new_n589));
  XOR2_X1   g388(.A(G183gat), .B(G211gat), .Z(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT99), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n589), .B(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n237), .B1(KEYINPUT21), .B2(new_n583), .ZN(new_n593));
  XNOR2_X1  g392(.A(KEYINPUT98), .B(KEYINPUT19), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n592), .A2(new_n596), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(KEYINPUT100), .B1(G85gat), .B2(G92gat), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT8), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n601), .B1(G99gat), .B2(G106gat), .ZN(new_n602));
  INV_X1    g401(.A(G85gat), .ZN(new_n603));
  INV_X1    g402(.A(G92gat), .ZN(new_n604));
  AOI211_X1 g403(.A(new_n600), .B(new_n602), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G99gat), .B(G106gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n607));
  NAND3_X1  g406(.A1(KEYINPUT101), .A2(G85gat), .A3(G92gat), .ZN(new_n608));
  MUX2_X1   g407(.A(new_n607), .B(KEYINPUT7), .S(new_n608), .Z(new_n609));
  NAND3_X1  g408(.A1(new_n605), .A2(new_n606), .A3(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n606), .B1(new_n605), .B2(new_n609), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AND2_X1   g412(.A1(G232gat), .A2(G233gat), .ZN(new_n614));
  AOI22_X1  g413(.A1(new_n229), .A2(new_n613), .B1(KEYINPUT41), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n250), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n615), .B1(new_n616), .B2(new_n613), .ZN(new_n617));
  XNOR2_X1  g416(.A(G190gat), .B(G218gat), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT102), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n614), .A2(KEYINPUT41), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(G134gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(new_n386), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n617), .A2(new_n618), .ZN(new_n625));
  AOI22_X1  g424(.A1(new_n621), .A2(new_n624), .B1(new_n625), .B2(new_n619), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n625), .A2(KEYINPUT102), .A3(new_n619), .A4(new_n624), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G230gat), .A2(G233gat), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n581), .B(new_n582), .Z(new_n632));
  OAI21_X1  g431(.A(new_n632), .B1(new_n611), .B2(new_n612), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT10), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n605), .A2(new_n609), .ZN(new_n635));
  INV_X1    g434(.A(new_n606), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n637), .A2(new_n610), .A3(new_n583), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n633), .A2(new_n634), .A3(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n613), .A2(KEYINPUT10), .A3(new_n583), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n631), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n633), .A2(new_n638), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n641), .B1(new_n642), .B2(new_n631), .ZN(new_n643));
  XNOR2_X1  g442(.A(G120gat), .B(G148gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(G176gat), .B(G204gat), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n644), .B(new_n645), .Z(new_n646));
  OR2_X1    g445(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n643), .A2(new_n646), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n599), .A2(new_n629), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n574), .A2(new_n575), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g452(.A(KEYINPUT103), .B(G1gat), .Z(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(G1324gat));
  INV_X1    g454(.A(new_n533), .ZN(new_n656));
  AND3_X1   g455(.A1(new_n574), .A2(new_n656), .A3(new_n652), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n657), .A2(new_n230), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n658), .B(KEYINPUT104), .Z(new_n659));
  XOR2_X1   g458(.A(KEYINPUT16), .B(G8gat), .Z(new_n660));
  NAND2_X1  g459(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT42), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n659), .A2(new_n662), .ZN(G1325gat));
  AND2_X1   g462(.A1(new_n574), .A2(new_n652), .ZN(new_n664));
  INV_X1    g463(.A(new_n541), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(G15gat), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n651), .A2(G15gat), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n574), .A2(new_n540), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(G1326gat));
  NAND2_X1  g469(.A1(new_n664), .A2(new_n536), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT43), .B(G22gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(G1327gat));
  NOR3_X1   g472(.A1(new_n599), .A2(new_n629), .A3(new_n649), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n574), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n675), .A2(new_n209), .A3(new_n575), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT45), .ZN(new_n677));
  INV_X1    g476(.A(new_n628), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n678), .A2(new_n626), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n537), .A2(new_n541), .A3(new_n572), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n486), .A2(new_n512), .A3(new_n523), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n446), .B1(new_n441), .B2(new_n442), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n451), .B1(new_n682), .B2(new_n445), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n681), .A2(new_n373), .A3(new_n683), .A4(new_n453), .ZN(new_n684));
  AOI22_X1  g483(.A1(new_n684), .A2(KEYINPUT35), .B1(new_n532), .B2(new_n533), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n679), .B1(new_n680), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n629), .B1(new_n535), .B2(new_n573), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(KEYINPUT44), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n599), .B(KEYINPUT105), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n692), .A2(new_n273), .A3(new_n649), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n691), .A2(new_n448), .A3(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n677), .B1(new_n209), .B2(new_n695), .ZN(G1328gat));
  NAND3_X1  g495(.A1(new_n675), .A2(new_n210), .A3(new_n656), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n697), .B(KEYINPUT46), .Z(new_n698));
  NOR3_X1   g497(.A1(new_n691), .A2(new_n533), .A3(new_n694), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n698), .B1(new_n210), .B2(new_n699), .ZN(G1329gat));
  NAND4_X1  g499(.A1(new_n688), .A2(new_n665), .A3(new_n690), .A4(new_n693), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT106), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n535), .A2(new_n573), .ZN(new_n704));
  AOI21_X1  g503(.A(KEYINPUT44), .B1(new_n704), .B2(new_n679), .ZN(new_n705));
  AOI211_X1 g504(.A(new_n687), .B(new_n629), .C1(new_n535), .C2(new_n573), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n707), .A2(KEYINPUT106), .A3(new_n665), .A4(new_n693), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n703), .A2(new_n708), .A3(G43gat), .ZN(new_n709));
  INV_X1    g508(.A(G43gat), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n675), .A2(new_n710), .A3(new_n540), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(KEYINPUT47), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n701), .A2(G43gat), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n711), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT47), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n714), .A2(new_n715), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n710), .B1(new_n701), .B2(new_n702), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n712), .B1(new_n721), .B2(new_n708), .ZN(new_n722));
  AOI21_X1  g521(.A(KEYINPUT47), .B1(new_n716), .B2(new_n711), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT107), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n720), .A2(new_n724), .ZN(G1330gat));
  INV_X1    g524(.A(G50gat), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n675), .A2(new_n726), .A3(new_n536), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n691), .A2(new_n486), .A3(new_n694), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n727), .B1(new_n728), .B2(new_n726), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT48), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(G1331gat));
  AND4_X1   g530(.A1(new_n704), .A2(new_n273), .A3(new_n629), .A4(new_n599), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n732), .A2(new_n649), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n575), .ZN(new_n734));
  XNOR2_X1  g533(.A(KEYINPUT108), .B(G57gat), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1332gat));
  NAND2_X1  g535(.A1(new_n733), .A2(new_n656), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n738));
  XOR2_X1   g537(.A(KEYINPUT49), .B(G64gat), .Z(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n737), .B2(new_n739), .ZN(G1333gat));
  NAND2_X1  g539(.A1(new_n733), .A2(new_n665), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n540), .A2(new_n649), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(G71gat), .ZN(new_n743));
  AOI22_X1  g542(.A1(new_n741), .A2(G71gat), .B1(new_n732), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g544(.A1(new_n733), .A2(new_n536), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(G78gat), .ZN(G1335gat));
  INV_X1    g546(.A(new_n273), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n748), .A2(new_n599), .A3(new_n650), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n707), .A2(new_n749), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n750), .A2(new_n575), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n748), .A2(new_n599), .ZN(new_n752));
  AND4_X1   g551(.A1(KEYINPUT51), .A2(new_n704), .A3(new_n679), .A4(new_n752), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT51), .B1(new_n689), .B2(new_n752), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n575), .A2(new_n603), .A3(new_n649), .ZN(new_n756));
  OAI22_X1  g555(.A1(new_n751), .A2(new_n603), .B1(new_n755), .B2(new_n756), .ZN(G1336gat));
  NAND3_X1  g556(.A1(new_n707), .A2(new_n656), .A3(new_n749), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(G92gat), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n656), .A2(new_n604), .A3(new_n649), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n759), .B1(new_n755), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT52), .ZN(G1337gat));
  AND2_X1   g561(.A1(new_n750), .A2(new_n665), .ZN(new_n763));
  XNOR2_X1  g562(.A(KEYINPUT109), .B(G99gat), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n540), .A2(new_n649), .A3(new_n764), .ZN(new_n765));
  OAI22_X1  g564(.A1(new_n763), .A2(new_n764), .B1(new_n755), .B2(new_n765), .ZN(G1338gat));
  NAND3_X1  g565(.A1(new_n707), .A2(new_n536), .A3(new_n749), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(G106gat), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT110), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n486), .A2(G106gat), .A3(new_n650), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(new_n753), .B2(new_n754), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n768), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g572(.A1(new_n652), .A2(new_n273), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n639), .A2(new_n640), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n630), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n639), .A2(new_n640), .A3(new_n631), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n776), .A2(KEYINPUT54), .A3(new_n777), .ZN(new_n778));
  XOR2_X1   g577(.A(KEYINPUT111), .B(KEYINPUT54), .Z(new_n779));
  AOI21_X1  g578(.A(new_n646), .B1(new_n641), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n778), .A2(KEYINPUT55), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n648), .ZN(new_n782));
  AOI21_X1  g581(.A(KEYINPUT55), .B1(new_n778), .B2(new_n780), .ZN(new_n783));
  OR2_X1    g582(.A1(new_n783), .A2(KEYINPUT112), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT112), .ZN(new_n785));
  AOI211_X1 g584(.A(new_n785), .B(KEYINPUT55), .C1(new_n778), .C2(new_n780), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n782), .B1(new_n784), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n258), .A2(new_n264), .A3(new_n270), .ZN(new_n789));
  OR2_X1    g588(.A1(new_n252), .A2(new_n253), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n239), .B1(new_n790), .B2(new_n238), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n265), .A2(new_n267), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n262), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n789), .A2(new_n793), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n788), .A2(new_n794), .A3(new_n679), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n789), .A2(new_n793), .A3(new_n649), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(KEYINPUT113), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n789), .A2(new_n793), .A3(new_n649), .A4(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n783), .A2(KEYINPUT112), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n648), .B(new_n781), .C1(new_n800), .C2(new_n786), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n797), .B(new_n799), .C1(new_n273), .C2(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n795), .B1(new_n802), .B2(new_n629), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n774), .B1(new_n803), .B2(new_n692), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(KEYINPUT114), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT114), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n774), .B(new_n806), .C1(new_n803), .C2(new_n692), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n808), .A2(new_n448), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n681), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n810), .A2(new_n656), .ZN(new_n811));
  AOI21_X1  g610(.A(G113gat), .B1(new_n811), .B2(new_n748), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n808), .A2(new_n536), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n540), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n575), .A2(new_n533), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n748), .A2(G113gat), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n812), .B1(new_n816), .B2(new_n817), .ZN(G1340gat));
  AOI21_X1  g617(.A(G120gat), .B1(new_n811), .B2(new_n649), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n649), .A2(G120gat), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n819), .B1(new_n816), .B2(new_n820), .ZN(G1341gat));
  AND3_X1   g620(.A1(new_n816), .A2(G127gat), .A3(new_n692), .ZN(new_n822));
  INV_X1    g621(.A(new_n599), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n810), .A2(new_n656), .A3(new_n823), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n824), .A2(KEYINPUT115), .ZN(new_n825));
  AOI21_X1  g624(.A(G127gat), .B1(new_n824), .B2(KEYINPUT115), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n822), .B1(new_n825), .B2(new_n826), .ZN(G1342gat));
  NAND2_X1  g626(.A1(new_n533), .A2(new_n679), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(KEYINPUT116), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n810), .A2(G134gat), .A3(new_n829), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(KEYINPUT56), .ZN(new_n831));
  INV_X1    g630(.A(G134gat), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n814), .A2(new_n629), .A3(new_n815), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(G1343gat));
  NOR2_X1   g633(.A1(new_n665), .A2(new_n486), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n809), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n836), .A2(new_n656), .ZN(new_n837));
  INV_X1    g636(.A(G141gat), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n837), .A2(new_n838), .A3(new_n748), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(KEYINPUT118), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n805), .A2(new_n536), .A3(new_n807), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT57), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n782), .A2(new_n783), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n843), .B1(new_n271), .B2(new_n272), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT117), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n844), .A2(new_n845), .A3(new_n796), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n629), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n845), .B1(new_n844), .B2(new_n796), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n823), .B1(new_n849), .B2(new_n795), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n774), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n486), .A2(new_n842), .ZN(new_n852));
  AOI22_X1  g651(.A1(new_n841), .A2(new_n842), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n541), .A2(new_n533), .A3(new_n575), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n853), .A2(new_n273), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n855), .A2(new_n391), .ZN(new_n856));
  OR3_X1    g655(.A1(new_n840), .A2(KEYINPUT58), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT58), .B1(new_n840), .B2(new_n856), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(G1344gat));
  NAND3_X1  g658(.A1(new_n837), .A2(new_n393), .A3(new_n649), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n853), .A2(new_n650), .A3(new_n854), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n861), .A2(KEYINPUT59), .A3(new_n393), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT59), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n805), .A2(new_n807), .A3(new_n852), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT119), .B1(new_n801), .B2(new_n629), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n788), .A2(new_n866), .A3(new_n679), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n865), .A2(new_n867), .A3(new_n794), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n868), .B1(new_n847), .B2(new_n848), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(KEYINPUT120), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT120), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n868), .B(new_n871), .C1(new_n847), .C2(new_n848), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n870), .A2(new_n823), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n486), .B1(new_n873), .B2(new_n774), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n864), .B1(new_n874), .B2(KEYINPUT57), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n854), .A2(new_n650), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n863), .B1(new_n877), .B2(G148gat), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n860), .B1(new_n862), .B2(new_n878), .ZN(G1345gat));
  NAND3_X1  g678(.A1(new_n837), .A2(new_n385), .A3(new_n599), .ZN(new_n880));
  INV_X1    g679(.A(new_n692), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n853), .A2(new_n881), .A3(new_n854), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n880), .B1(new_n882), .B2(new_n385), .ZN(G1346gat));
  NOR3_X1   g682(.A1(new_n853), .A2(new_n629), .A3(new_n854), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n829), .A2(G162gat), .ZN(new_n885));
  OAI22_X1  g684(.A1(new_n884), .A2(new_n386), .B1(new_n836), .B2(new_n885), .ZN(G1347gat));
  NAND3_X1  g685(.A1(new_n805), .A2(new_n448), .A3(new_n807), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n533), .B1(new_n887), .B2(KEYINPUT121), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT121), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n805), .A2(new_n889), .A3(new_n448), .A4(new_n807), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n888), .A2(new_n681), .A3(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(G169gat), .B1(new_n892), .B2(new_n748), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n656), .A2(new_n448), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n814), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n273), .A2(new_n312), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n893), .B1(new_n895), .B2(new_n896), .ZN(G1348gat));
  AOI21_X1  g696(.A(G176gat), .B1(new_n892), .B2(new_n649), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n894), .A2(new_n742), .A3(new_n313), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n898), .B1(new_n813), .B2(new_n899), .ZN(G1349gat));
  INV_X1    g699(.A(new_n895), .ZN(new_n901));
  OAI21_X1  g700(.A(G183gat), .B1(new_n901), .B2(new_n881), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n599), .A2(new_n305), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n892), .A2(KEYINPUT122), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT122), .B1(new_n892), .B2(new_n903), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n902), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(KEYINPUT60), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT60), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n902), .B(new_n908), .C1(new_n904), .C2(new_n905), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(G1350gat));
  NAND2_X1  g709(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n911));
  NOR2_X1   g710(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n895), .A2(new_n679), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n913), .B1(new_n914), .B2(G190gat), .ZN(new_n915));
  AOI211_X1 g714(.A(new_n300), .B(new_n912), .C1(new_n895), .C2(new_n679), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n911), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n891), .A2(G190gat), .A3(new_n629), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT123), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(G1351gat));
  AND2_X1   g719(.A1(new_n888), .A2(new_n890), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n921), .A2(new_n835), .ZN(new_n922));
  AOI21_X1  g721(.A(G197gat), .B1(new_n922), .B2(new_n748), .ZN(new_n923));
  OAI211_X1 g722(.A(KEYINPUT125), .B(new_n864), .C1(new_n874), .C2(KEYINPUT57), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n665), .A2(new_n894), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n599), .B1(new_n869), .B2(KEYINPUT120), .ZN(new_n927));
  AOI22_X1  g726(.A1(new_n927), .A2(new_n872), .B1(new_n273), .B2(new_n652), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n842), .B1(new_n928), .B2(new_n486), .ZN(new_n929));
  AOI21_X1  g728(.A(KEYINPUT125), .B1(new_n929), .B2(new_n864), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n273), .A2(new_n277), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n923), .B1(new_n931), .B2(new_n932), .ZN(G1352gat));
  NAND4_X1  g732(.A1(new_n921), .A2(new_n278), .A3(new_n649), .A4(new_n835), .ZN(new_n934));
  XOR2_X1   g733(.A(new_n934), .B(KEYINPUT62), .Z(new_n935));
  NAND2_X1  g734(.A1(new_n931), .A2(new_n649), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(G204gat), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n935), .A2(new_n937), .ZN(G1353gat));
  INV_X1    g737(.A(G211gat), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n922), .A2(new_n939), .A3(new_n599), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n665), .A2(new_n823), .A3(new_n894), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n939), .B1(new_n875), .B2(new_n941), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n942), .B(KEYINPUT63), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n940), .A2(new_n943), .ZN(G1354gat));
  OAI21_X1  g743(.A(KEYINPUT126), .B1(new_n926), .B2(new_n930), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT125), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n875), .A2(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT126), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n947), .A2(new_n948), .A3(new_n925), .A4(new_n924), .ZN(new_n949));
  INV_X1    g748(.A(G218gat), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n629), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n945), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n921), .A2(new_n679), .A3(new_n835), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(new_n950), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT127), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n952), .A2(KEYINPUT127), .A3(new_n954), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1355gat));
endmodule


