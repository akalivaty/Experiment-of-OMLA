//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 0 0 0 1 1 1 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n832, new_n833, new_n834, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950;
  XOR2_X1   g000(.A(G15gat), .B(G22gat), .Z(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G15gat), .B(G22gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n205), .B1(new_n206), .B2(G1gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT88), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n204), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G8gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n209), .B(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G57gat), .B(G64gat), .ZN(new_n212));
  AOI21_X1  g011(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G71gat), .B(G78gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n214), .B(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT21), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n211), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n219), .B(G183gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(G127gat), .B(G155gat), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n220), .B(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(G231gat), .A2(G233gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n223), .B(KEYINPUT91), .ZN(new_n224));
  XOR2_X1   g023(.A(KEYINPUT92), .B(G211gat), .Z(new_n225));
  XOR2_X1   g024(.A(new_n224), .B(new_n225), .Z(new_n226));
  XNOR2_X1  g025(.A(new_n222), .B(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n217), .A2(new_n218), .ZN(new_n228));
  XNOR2_X1  g027(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n229));
  XOR2_X1   g028(.A(new_n228), .B(new_n229), .Z(new_n230));
  NAND2_X1  g029(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n226), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n222), .B(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n230), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n231), .A2(new_n235), .ZN(new_n236));
  XOR2_X1   g035(.A(G134gat), .B(G162gat), .Z(new_n237));
  AND2_X1   g036(.A1(G232gat), .A2(G233gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n238), .A2(KEYINPUT41), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n237), .B(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(G29gat), .ZN(new_n241));
  INV_X1    g040(.A(G36gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NOR2_X1   g042(.A1(G29gat), .A2(G36gat), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT14), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT87), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n243), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n244), .B(KEYINPUT14), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT87), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(G43gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(G50gat), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT15), .B1(new_n253), .B2(KEYINPUT86), .ZN(new_n254));
  INV_X1    g053(.A(G50gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(G43gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(new_n253), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n254), .B(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(KEYINPUT15), .B1(new_n249), .B2(new_n243), .ZN(new_n259));
  OAI22_X1  g058(.A1(new_n251), .A2(new_n258), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n260), .B(KEYINPUT17), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT93), .ZN(new_n262));
  INV_X1    g061(.A(G99gat), .ZN(new_n263));
  INV_X1    g062(.A(G106gat), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(KEYINPUT93), .A2(G99gat), .A3(G106gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(KEYINPUT8), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(G85gat), .A2(G92gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(KEYINPUT7), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n267), .B(new_n269), .C1(G85gat), .C2(G92gat), .ZN(new_n270));
  XOR2_X1   g069(.A(G99gat), .B(G106gat), .Z(new_n271));
  OR2_X1    g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(new_n271), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n261), .A2(new_n274), .ZN(new_n275));
  XOR2_X1   g074(.A(G190gat), .B(G218gat), .Z(new_n276));
  NAND2_X1  g075(.A1(new_n238), .A2(KEYINPUT41), .ZN(new_n277));
  INV_X1    g076(.A(new_n274), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(new_n260), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n275), .A2(new_n276), .A3(new_n277), .A4(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT94), .ZN(new_n281));
  AOI22_X1  g080(.A1(new_n261), .A2(new_n274), .B1(KEYINPUT41), .B2(new_n238), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT94), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n282), .A2(new_n283), .A3(new_n276), .A4(new_n279), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT95), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n240), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AND2_X1   g086(.A1(new_n282), .A2(new_n279), .ZN(new_n288));
  OR2_X1    g087(.A1(new_n288), .A2(new_n276), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(new_n285), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n289), .B(new_n285), .C1(new_n286), .C2(new_n240), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n236), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n216), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n274), .A2(new_n217), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(G230gat), .A2(G233gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n298), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT10), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n295), .A2(new_n301), .A3(new_n296), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n278), .A2(KEYINPUT10), .A3(new_n216), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n300), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT96), .ZN(new_n305));
  NOR3_X1   g104(.A1(new_n299), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n299), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n307), .A2(KEYINPUT96), .ZN(new_n308));
  XOR2_X1   g107(.A(G120gat), .B(G148gat), .Z(new_n309));
  XNOR2_X1  g108(.A(G176gat), .B(G204gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n309), .B(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT97), .B(KEYINPUT98), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  OR3_X1    g112(.A1(new_n306), .A2(new_n308), .A3(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n313), .B1(new_n308), .B2(new_n306), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n211), .ZN(new_n318));
  AND2_X1   g117(.A1(new_n318), .A2(new_n260), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n319), .B1(new_n261), .B2(new_n211), .ZN(new_n320));
  NAND2_X1  g119(.A1(G229gat), .A2(G233gat), .ZN(new_n321));
  AND3_X1   g120(.A1(new_n320), .A2(KEYINPUT18), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(KEYINPUT18), .B1(new_n320), .B2(new_n321), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(KEYINPUT11), .B(G169gat), .ZN(new_n325));
  INV_X1    g124(.A(G197gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n325), .B(new_n326), .ZN(new_n327));
  XOR2_X1   g126(.A(G113gat), .B(G141gat), .Z(new_n328));
  XNOR2_X1  g127(.A(new_n327), .B(new_n328), .ZN(new_n329));
  XOR2_X1   g128(.A(new_n329), .B(KEYINPUT12), .Z(new_n330));
  INV_X1    g129(.A(KEYINPUT89), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n211), .B(new_n260), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n321), .B(KEYINPUT13), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n333), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n318), .A2(new_n260), .ZN(new_n336));
  OAI211_X1 g135(.A(KEYINPUT89), .B(new_n335), .C1(new_n319), .C2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n324), .A2(KEYINPUT90), .A3(new_n330), .A4(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n320), .A2(new_n321), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT18), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n320), .A2(KEYINPUT18), .A3(new_n321), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n342), .A2(new_n330), .A3(new_n338), .A4(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT90), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n339), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n324), .A2(new_n338), .ZN(new_n348));
  INV_X1    g147(.A(new_n330), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n317), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT79), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT71), .ZN(new_n354));
  XOR2_X1   g153(.A(G211gat), .B(G218gat), .Z(new_n355));
  INV_X1    g154(.A(G204gat), .ZN(new_n356));
  AND2_X1   g155(.A1(KEYINPUT68), .A2(G197gat), .ZN(new_n357));
  NOR2_X1   g156(.A1(KEYINPUT68), .A2(G197gat), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT68), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(new_n326), .ZN(new_n361));
  NAND2_X1  g160(.A1(KEYINPUT68), .A2(G197gat), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n361), .A2(G204gat), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT70), .ZN(new_n365));
  OR2_X1    g164(.A1(KEYINPUT69), .A2(KEYINPUT22), .ZN(new_n366));
  NAND2_X1  g165(.A1(G211gat), .A2(G218gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(KEYINPUT69), .A2(KEYINPUT22), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  AND3_X1   g168(.A1(new_n364), .A2(new_n365), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n365), .B1(new_n364), .B2(new_n369), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n354), .B(new_n355), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n355), .ZN(new_n373));
  NOR3_X1   g172(.A1(new_n357), .A2(new_n358), .A3(new_n356), .ZN(new_n374));
  AOI21_X1  g173(.A(G204gat), .B1(new_n361), .B2(new_n362), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n369), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT70), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n364), .A2(new_n365), .A3(new_n369), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n373), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT71), .B1(new_n376), .B2(new_n355), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n372), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT74), .ZN(new_n382));
  INV_X1    g181(.A(G141gat), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n383), .A2(G148gat), .ZN(new_n384));
  INV_X1    g183(.A(G148gat), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n385), .A2(G141gat), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n382), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(G155gat), .A2(G162gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT2), .ZN(new_n389));
  NOR2_X1   g188(.A1(G155gat), .A2(G162gat), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(new_n388), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n385), .A2(G141gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n383), .A2(G148gat), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(new_n394), .A3(KEYINPUT74), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n387), .A2(new_n389), .A3(new_n392), .A4(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT3), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n389), .B1(new_n384), .B2(new_n386), .ZN(new_n398));
  INV_X1    g197(.A(new_n388), .ZN(new_n399));
  OAI21_X1  g198(.A(KEYINPUT73), .B1(new_n399), .B2(new_n390), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT73), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n391), .A2(new_n401), .A3(new_n388), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n398), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n396), .A2(new_n397), .A3(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(KEYINPUT72), .B(KEYINPUT29), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n396), .A2(new_n403), .ZN(new_n408));
  AND3_X1   g207(.A1(new_n364), .A2(new_n373), .A3(new_n369), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n373), .B1(new_n364), .B2(new_n369), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n406), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(new_n397), .ZN(new_n412));
  AOI22_X1  g211(.A1(new_n381), .A2(new_n407), .B1(new_n408), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(G228gat), .A2(G233gat), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n353), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n355), .B1(new_n370), .B2(new_n371), .ZN(new_n417));
  INV_X1    g216(.A(new_n380), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n419), .A2(new_n372), .B1(new_n404), .B2(new_n406), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n396), .A2(new_n403), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n421), .B1(new_n411), .B2(new_n397), .ZN(new_n422));
  OAI211_X1 g221(.A(KEYINPUT79), .B(new_n414), .C1(new_n420), .C2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n416), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n408), .A2(KEYINPUT3), .ZN(new_n425));
  OR2_X1    g224(.A1(new_n421), .A2(KEYINPUT29), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n425), .B1(new_n381), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT80), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI211_X1 g228(.A(KEYINPUT80), .B(new_n425), .C1(new_n381), .C2(new_n426), .ZN(new_n430));
  INV_X1    g229(.A(new_n420), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n429), .A2(new_n415), .A3(new_n430), .A4(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(G22gat), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n424), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n433), .B1(new_n424), .B2(new_n432), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT81), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n424), .A2(new_n432), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(G22gat), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT81), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n424), .A2(new_n432), .A3(new_n433), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(G78gat), .B(G106gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(KEYINPUT31), .B(G50gat), .ZN(new_n443));
  XOR2_X1   g242(.A(new_n442), .B(new_n443), .Z(new_n444));
  NAND3_X1  g243(.A1(new_n436), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n444), .ZN(new_n446));
  OAI211_X1 g245(.A(KEYINPUT81), .B(new_n446), .C1(new_n434), .C2(new_n435), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT82), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(KEYINPUT77), .B(KEYINPUT5), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(G120gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(G113gat), .ZN(new_n454));
  INV_X1    g253(.A(G113gat), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(G120gat), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT66), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT1), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(G127gat), .B(G134gat), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n457), .A2(new_n461), .A3(new_n458), .A4(new_n459), .ZN(new_n464));
  AND2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n421), .A2(new_n465), .A3(KEYINPUT76), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n463), .A2(new_n464), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n408), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n396), .A2(new_n463), .A3(new_n403), .A4(new_n464), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT76), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n466), .A2(new_n468), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(G225gat), .A2(G233gat), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n452), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  XOR2_X1   g274(.A(KEYINPUT75), .B(KEYINPUT4), .Z(new_n476));
  AND2_X1   g275(.A1(new_n469), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n466), .A2(new_n471), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT4), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n425), .A2(new_n467), .A3(new_n404), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(new_n473), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n475), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  XNOR2_X1  g282(.A(KEYINPUT0), .B(G57gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n484), .B(G85gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(G1gat), .B(G29gat), .ZN(new_n486));
  XOR2_X1   g285(.A(new_n485), .B(new_n486), .Z(new_n487));
  OAI22_X1  g286(.A1(new_n478), .A2(new_n479), .B1(new_n469), .B2(new_n476), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n482), .A2(new_n451), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n483), .A2(new_n487), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT78), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n483), .A2(new_n490), .ZN(new_n493));
  INV_X1    g292(.A(new_n487), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT6), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT78), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n483), .A2(new_n497), .A3(new_n487), .A4(new_n490), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n492), .A2(new_n495), .A3(new_n496), .A4(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n493), .A2(KEYINPUT6), .A3(new_n494), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  XOR2_X1   g300(.A(G8gat), .B(G36gat), .Z(new_n502));
  XNOR2_X1  g301(.A(new_n502), .B(G64gat), .ZN(new_n503));
  INV_X1    g302(.A(G92gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n503), .B(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(KEYINPUT64), .A2(KEYINPUT25), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(G169gat), .ZN(new_n509));
  INV_X1    g308(.A(G176gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT23), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT24), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n514), .A2(G183gat), .A3(G190gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(G183gat), .A2(G190gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT24), .ZN(new_n517));
  NOR2_X1   g316(.A1(G183gat), .A2(G190gat), .ZN(new_n518));
  OAI221_X1 g317(.A(new_n515), .B1(new_n509), .B2(new_n510), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n508), .B1(new_n513), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n517), .A2(new_n518), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n509), .A2(new_n510), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n511), .B(KEYINPUT23), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n523), .A2(new_n524), .A3(new_n507), .A4(new_n515), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT64), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT25), .ZN(new_n527));
  AOI22_X1  g326(.A1(new_n520), .A2(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(KEYINPUT27), .B(G183gat), .ZN(new_n529));
  INV_X1    g328(.A(G190gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT28), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n529), .A2(KEYINPUT28), .A3(new_n530), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NOR3_X1   g334(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(KEYINPUT65), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n522), .B1(KEYINPUT26), .B2(new_n511), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AND3_X1   g338(.A1(new_n535), .A2(new_n539), .A3(new_n516), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n528), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G226gat), .A2(G233gat), .ZN(new_n542));
  OR2_X1    g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n542), .B1(new_n541), .B2(new_n405), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n543), .A2(new_n381), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n542), .B1(new_n541), .B2(KEYINPUT29), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n381), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n506), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n543), .A2(new_n547), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n545), .B(new_n505), .C1(new_n550), .C2(new_n381), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n549), .A2(new_n551), .A3(KEYINPUT30), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n545), .B1(new_n550), .B2(new_n381), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT30), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n553), .A2(new_n554), .A3(new_n506), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n501), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n445), .A2(KEYINPUT82), .A3(new_n447), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n450), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n448), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT37), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n553), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g361(.A(KEYINPUT37), .B(new_n545), .C1(new_n550), .C2(new_n381), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(new_n505), .A3(new_n563), .ZN(new_n564));
  XOR2_X1   g363(.A(KEYINPUT85), .B(KEYINPUT38), .Z(new_n565));
  AOI22_X1  g364(.A1(new_n564), .A2(new_n565), .B1(new_n553), .B2(new_n506), .ZN(new_n566));
  AOI21_X1  g365(.A(KEYINPUT84), .B1(new_n493), .B2(new_n494), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT84), .ZN(new_n568));
  AOI211_X1 g367(.A(new_n568), .B(new_n487), .C1(new_n483), .C2(new_n490), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n492), .A2(new_n498), .A3(new_n496), .ZN(new_n571));
  OR2_X1    g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n550), .A2(new_n381), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n543), .A2(new_n544), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n573), .B(KEYINPUT37), .C1(new_n381), .C2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n565), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n575), .A2(new_n562), .A3(new_n505), .A4(new_n576), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n566), .A2(new_n572), .A3(new_n500), .A4(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT83), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n473), .B1(new_n488), .B2(new_n481), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT39), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n472), .A2(new_n474), .ZN(new_n582));
  OR3_X1    g381(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n494), .B1(new_n580), .B2(new_n581), .ZN(new_n584));
  AOI21_X1  g383(.A(KEYINPUT40), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n570), .B1(new_n579), .B2(new_n585), .ZN(new_n586));
  OR2_X1    g385(.A1(new_n585), .A2(new_n579), .ZN(new_n587));
  INV_X1    g386(.A(new_n556), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n583), .A2(KEYINPUT40), .A3(new_n584), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n586), .A2(new_n587), .A3(new_n588), .A4(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n560), .A2(new_n578), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n535), .A2(new_n539), .A3(new_n516), .ZN(new_n592));
  AND2_X1   g391(.A1(new_n520), .A2(new_n525), .ZN(new_n593));
  NOR2_X1   g392(.A1(KEYINPUT64), .A2(KEYINPUT25), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n465), .B(new_n592), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n467), .B1(new_n528), .B2(new_n540), .ZN(new_n596));
  INV_X1    g395(.A(G227gat), .ZN(new_n597));
  INV_X1    g396(.A(G233gat), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n595), .A2(new_n596), .A3(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n601), .B(KEYINPUT34), .Z(new_n602));
  AOI21_X1  g401(.A(new_n600), .B1(new_n595), .B2(new_n596), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT32), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G15gat), .B(G43gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(G71gat), .B(G99gat), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n607), .B(new_n608), .Z(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n596), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(new_n599), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT33), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n610), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n606), .A2(new_n614), .ZN(new_n615));
  AOI221_X4 g414(.A(new_n604), .B1(KEYINPUT33), .B2(new_n609), .C1(new_n611), .C2(new_n599), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT67), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n602), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n609), .B1(new_n603), .B2(KEYINPUT33), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n621), .A2(new_n605), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n602), .B(new_n619), .C1(new_n622), .C2(new_n616), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(KEYINPUT36), .B1(new_n620), .B2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n601), .B(KEYINPUT34), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n615), .A2(new_n626), .A3(new_n617), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n602), .B1(new_n622), .B2(new_n616), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT36), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n625), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n559), .A2(new_n591), .A3(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT35), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n500), .B1(new_n570), .B2(new_n571), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n627), .A2(new_n628), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n635), .A2(new_n556), .A3(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n634), .B1(new_n448), .B2(new_n637), .ZN(new_n638));
  AND3_X1   g437(.A1(new_n501), .A2(KEYINPUT35), .A3(new_n556), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n619), .B1(new_n622), .B2(new_n616), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(new_n626), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(new_n623), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n639), .A2(new_n445), .A3(new_n642), .A4(new_n447), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  AOI211_X1 g443(.A(new_n294), .B(new_n352), .C1(new_n633), .C2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n501), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g447(.A1(new_n645), .A2(new_n588), .ZN(new_n649));
  NAND2_X1  g448(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n206), .A2(new_n210), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT42), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n653), .B1(new_n210), .B2(new_n649), .ZN(G1325gat));
  AOI21_X1  g453(.A(G15gat), .B1(new_n645), .B2(new_n636), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT99), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n656), .B1(new_n625), .B2(new_n631), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n629), .B1(new_n641), .B2(new_n623), .ZN(new_n658));
  NOR3_X1   g457(.A1(new_n658), .A2(KEYINPUT99), .A3(new_n630), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(G15gat), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n662), .B(KEYINPUT100), .Z(new_n663));
  AOI21_X1  g462(.A(new_n655), .B1(new_n645), .B2(new_n663), .ZN(G1326gat));
  NAND2_X1  g463(.A1(new_n450), .A2(new_n558), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n645), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT43), .B(G22gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1327gat));
  AOI21_X1  g468(.A(new_n293), .B1(new_n633), .B2(new_n644), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n352), .A2(new_n236), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n670), .A2(new_n241), .A3(new_n646), .A4(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT45), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n559), .A2(new_n591), .A3(new_n660), .ZN(new_n674));
  AND3_X1   g473(.A1(new_n638), .A2(new_n643), .A3(KEYINPUT101), .ZN(new_n675));
  AOI21_X1  g474(.A(KEYINPUT101), .B1(new_n638), .B2(new_n643), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n674), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n291), .A2(new_n292), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT44), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AOI211_X1 g480(.A(new_n680), .B(new_n293), .C1(new_n633), .C2(new_n644), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n681), .A2(new_n671), .A3(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n684), .A2(new_n501), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n673), .B1(new_n685), .B2(new_n241), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT102), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OAI211_X1 g487(.A(new_n673), .B(KEYINPUT102), .C1(new_n685), .C2(new_n241), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(G1328gat));
  INV_X1    g489(.A(KEYINPUT104), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n691), .B1(new_n684), .B2(new_n556), .ZN(new_n692));
  AOI21_X1  g491(.A(KEYINPUT44), .B1(new_n677), .B2(new_n678), .ZN(new_n693));
  INV_X1    g492(.A(new_n671), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n693), .A2(new_n682), .A3(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n695), .A2(KEYINPUT104), .A3(new_n588), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n692), .A2(G36gat), .A3(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT103), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n556), .B1(new_n698), .B2(KEYINPUT46), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n670), .A2(new_n242), .A3(new_n671), .A4(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n698), .A2(KEYINPUT46), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n697), .A2(new_n702), .ZN(G1329gat));
  INV_X1    g502(.A(KEYINPUT105), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n704), .B1(new_n684), .B2(new_n660), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n695), .A2(KEYINPUT105), .A3(new_n661), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n705), .A2(G43gat), .A3(new_n706), .ZN(new_n707));
  AND4_X1   g506(.A1(new_n252), .A2(new_n670), .A3(new_n636), .A4(new_n671), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT47), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n252), .B1(new_n695), .B2(new_n661), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n709), .B1(new_n712), .B2(new_n708), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(new_n713), .ZN(G1330gat));
  OAI21_X1  g513(.A(G50gat), .B1(new_n684), .B2(new_n560), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n670), .A2(new_n255), .A3(new_n666), .A4(new_n671), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n715), .A2(KEYINPUT48), .A3(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n716), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n695), .A2(new_n666), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n718), .B1(new_n719), .B2(G50gat), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n717), .B1(new_n720), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR3_X1   g520(.A1(new_n294), .A2(new_n317), .A3(new_n351), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n677), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n501), .B(KEYINPUT106), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XOR2_X1   g524(.A(new_n725), .B(G57gat), .Z(G1332gat));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n677), .A2(KEYINPUT107), .A3(new_n722), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n556), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n731));
  AND2_X1   g530(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n733), .B1(new_n730), .B2(new_n731), .ZN(G1333gat));
  INV_X1    g533(.A(G71gat), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n627), .A2(new_n628), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n735), .B1(new_n723), .B2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT108), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n728), .A2(new_n729), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n660), .A2(new_n735), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n677), .A2(KEYINPUT107), .A3(new_n722), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT107), .B1(new_n677), .B2(new_n722), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n738), .B(new_n740), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n737), .B1(new_n741), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(KEYINPUT50), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT50), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n748), .B(new_n737), .C1(new_n741), .C2(new_n745), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n749), .ZN(G1334gat));
  NAND2_X1  g549(.A1(new_n739), .A2(new_n666), .ZN(new_n751));
  XNOR2_X1  g550(.A(KEYINPUT109), .B(G78gat), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n751), .B(new_n752), .ZN(G1335gat));
  NOR2_X1   g552(.A1(new_n236), .A2(new_n351), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(KEYINPUT51), .B1(new_n679), .B2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT51), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n677), .A2(new_n757), .A3(new_n678), .A4(new_n754), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n756), .A2(new_n646), .A3(new_n316), .A4(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(G85gat), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n693), .A2(new_n682), .A3(new_n755), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n762), .A2(G85gat), .A3(new_n646), .A4(new_n316), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT110), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n761), .A2(new_n763), .A3(KEYINPUT110), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(G1336gat));
  NAND4_X1  g567(.A1(new_n756), .A2(new_n588), .A3(new_n316), .A4(new_n758), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n504), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n762), .A2(G92gat), .A3(new_n588), .A4(new_n316), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n770), .A2(new_n771), .A3(KEYINPUT52), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(G1337gat));
  AND3_X1   g575(.A1(new_n756), .A2(new_n316), .A3(new_n758), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n777), .A2(new_n263), .A3(new_n636), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n681), .A2(new_n683), .A3(new_n316), .A4(new_n754), .ZN(new_n779));
  OAI21_X1  g578(.A(G99gat), .B1(new_n779), .B2(new_n660), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(G1338gat));
  NOR2_X1   g580(.A1(new_n560), .A2(G106gat), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n777), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(G106gat), .B1(new_n779), .B2(new_n560), .ZN(new_n784));
  XOR2_X1   g583(.A(KEYINPUT111), .B(KEYINPUT53), .Z(new_n785));
  NAND3_X1  g584(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n762), .A2(new_n666), .A3(new_n316), .ZN(new_n787));
  AOI22_X1  g586(.A1(G106gat), .A2(new_n787), .B1(new_n777), .B2(new_n782), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT53), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n786), .B1(new_n788), .B2(new_n789), .ZN(G1339gat));
  INV_X1    g589(.A(KEYINPUT113), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n347), .A2(new_n350), .ZN(new_n792));
  AND4_X1   g591(.A1(new_n293), .A2(new_n792), .A3(new_n236), .A4(new_n317), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n332), .A2(new_n333), .ZN(new_n794));
  XOR2_X1   g593(.A(new_n794), .B(KEYINPUT112), .Z(new_n795));
  OR2_X1    g594(.A1(new_n320), .A2(new_n321), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n329), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n797), .B1(new_n339), .B2(new_n346), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n313), .B1(new_n304), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n302), .A2(new_n300), .A3(new_n303), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(KEYINPUT54), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n800), .B1(new_n304), .B2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n800), .B(KEYINPUT55), .C1(new_n304), .C2(new_n802), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n805), .A2(new_n315), .A3(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n678), .A2(new_n798), .A3(new_n808), .ZN(new_n809));
  AOI22_X1  g608(.A1(new_n351), .A2(new_n808), .B1(new_n798), .B2(new_n316), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n809), .B1(new_n810), .B2(new_n678), .ZN(new_n811));
  INV_X1    g610(.A(new_n236), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n793), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n813), .A2(new_n666), .A3(new_n736), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n588), .A2(new_n501), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n351), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n791), .B1(new_n818), .B2(G113gat), .ZN(new_n819));
  AOI211_X1 g618(.A(KEYINPUT113), .B(new_n455), .C1(new_n817), .C2(new_n351), .ZN(new_n820));
  INV_X1    g619(.A(new_n813), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n724), .A2(new_n588), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n560), .A2(new_n642), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT114), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n351), .A2(new_n455), .ZN(new_n827));
  OAI22_X1  g626(.A1(new_n819), .A2(new_n820), .B1(new_n826), .B2(new_n827), .ZN(G1340gat));
  OAI21_X1  g627(.A(G120gat), .B1(new_n816), .B2(new_n317), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n316), .A2(new_n453), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n829), .B1(new_n826), .B2(new_n830), .ZN(G1341gat));
  AOI21_X1  g630(.A(G127gat), .B1(new_n825), .B2(new_n236), .ZN(new_n832));
  INV_X1    g631(.A(G127gat), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n816), .A2(new_n833), .A3(new_n812), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n832), .A2(new_n834), .ZN(G1342gat));
  NOR2_X1   g634(.A1(new_n293), .A2(G134gat), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n825), .A2(new_n836), .ZN(new_n837));
  OR3_X1    g636(.A1(new_n837), .A2(KEYINPUT115), .A3(KEYINPUT56), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(KEYINPUT56), .ZN(new_n839));
  OAI21_X1  g638(.A(G134gat), .B1(new_n816), .B2(new_n293), .ZN(new_n840));
  OAI21_X1  g639(.A(KEYINPUT115), .B1(new_n837), .B2(KEYINPUT56), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n838), .A2(new_n839), .A3(new_n840), .A4(new_n841), .ZN(G1343gat));
  OAI21_X1  g641(.A(KEYINPUT57), .B1(new_n813), .B2(new_n665), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n660), .A2(new_n815), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n821), .A2(new_n846), .A3(new_n448), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n351), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(G141gat), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n823), .A2(new_n560), .A3(new_n661), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(new_n383), .A3(new_n351), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT58), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT58), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n849), .A2(new_n854), .A3(new_n851), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n853), .A2(new_n855), .ZN(G1344gat));
  OAI21_X1  g655(.A(KEYINPUT57), .B1(new_n813), .B2(new_n560), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT117), .B1(new_n293), .B2(new_n807), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n808), .A2(new_n859), .A3(new_n292), .A4(new_n291), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n858), .A2(new_n860), .A3(new_n798), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n798), .A2(new_n316), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n807), .B1(new_n347), .B2(new_n350), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n293), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n236), .B1(new_n861), .B2(new_n864), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n846), .B(new_n666), .C1(new_n865), .C2(new_n793), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n857), .A2(new_n866), .A3(new_n316), .A4(new_n844), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(G148gat), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(KEYINPUT59), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n868), .A2(KEYINPUT118), .A3(KEYINPUT59), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n845), .A2(new_n847), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n873), .B(G148gat), .C1(new_n874), .C2(new_n317), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n871), .A2(new_n872), .A3(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n850), .A2(new_n385), .A3(new_n316), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT116), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n877), .B(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n876), .A2(new_n879), .ZN(G1345gat));
  AOI21_X1  g679(.A(G155gat), .B1(new_n850), .B2(new_n236), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n874), .A2(new_n812), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n881), .B1(new_n882), .B2(G155gat), .ZN(G1346gat));
  INV_X1    g682(.A(G162gat), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n850), .A2(new_n884), .A3(new_n678), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT119), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT120), .B1(new_n874), .B2(new_n293), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT120), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n845), .A2(new_n888), .A3(new_n678), .A4(new_n847), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n887), .A2(G162gat), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n886), .A2(new_n890), .ZN(G1347gat));
  NAND2_X1  g690(.A1(new_n724), .A2(new_n588), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n814), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(G169gat), .B1(new_n894), .B2(new_n792), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n813), .A2(new_n646), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n896), .A2(new_n588), .A3(new_n560), .A4(new_n642), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n897), .A2(G169gat), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n895), .B1(new_n898), .B2(new_n792), .ZN(G1348gat));
  OAI21_X1  g698(.A(new_n510), .B1(new_n897), .B2(new_n317), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT121), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n894), .A2(new_n510), .A3(new_n317), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n901), .A2(new_n902), .ZN(G1349gat));
  OAI21_X1  g702(.A(G183gat), .B1(new_n894), .B2(new_n812), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n236), .A2(new_n529), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n897), .B2(new_n905), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g706(.A(G190gat), .B1(new_n894), .B2(new_n293), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n908), .A2(KEYINPUT61), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n908), .A2(KEYINPUT61), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n678), .A2(new_n530), .ZN(new_n911));
  OAI22_X1  g710(.A1(new_n909), .A2(new_n910), .B1(new_n897), .B2(new_n911), .ZN(G1351gat));
  NAND3_X1  g711(.A1(new_n660), .A2(new_n588), .A3(new_n448), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(KEYINPUT122), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n896), .A2(new_n915), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n914), .A2(KEYINPUT122), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n916), .A2(new_n326), .A3(new_n351), .A4(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n893), .A2(new_n660), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT123), .ZN(new_n920));
  AND4_X1   g719(.A1(new_n351), .A2(new_n857), .A3(new_n920), .A4(new_n866), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n918), .B1(new_n326), .B2(new_n921), .ZN(G1352gat));
  NAND4_X1  g721(.A1(new_n916), .A2(new_n356), .A3(new_n316), .A4(new_n917), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT124), .ZN(new_n924));
  OR3_X1    g723(.A1(new_n923), .A2(new_n924), .A3(KEYINPUT62), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n857), .A2(new_n920), .A3(new_n866), .A4(new_n316), .ZN(new_n926));
  AOI22_X1  g725(.A1(new_n923), .A2(KEYINPUT62), .B1(G204gat), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n924), .B1(new_n923), .B2(KEYINPUT62), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n925), .A2(new_n927), .A3(new_n928), .ZN(G1353gat));
  NAND4_X1  g728(.A1(new_n857), .A2(new_n920), .A3(new_n866), .A4(new_n236), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(G211gat), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n931), .A2(KEYINPUT125), .A3(KEYINPUT63), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n812), .A2(G211gat), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n916), .A2(new_n917), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(KEYINPUT125), .A2(KEYINPUT63), .ZN(new_n935));
  OR2_X1    g734(.A1(KEYINPUT125), .A2(KEYINPUT63), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n930), .A2(G211gat), .A3(new_n935), .A4(new_n936), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n932), .A2(new_n934), .A3(new_n937), .ZN(G1354gat));
  NAND4_X1  g737(.A1(new_n917), .A2(new_n896), .A3(new_n678), .A4(new_n915), .ZN(new_n939));
  INV_X1    g738(.A(G218gat), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(KEYINPUT126), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT126), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n939), .A2(new_n943), .A3(new_n940), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n293), .A2(new_n940), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n857), .A2(new_n920), .A3(new_n866), .A4(new_n945), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n942), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT127), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g748(.A1(new_n942), .A2(KEYINPUT127), .A3(new_n944), .A4(new_n946), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(G1355gat));
endmodule


