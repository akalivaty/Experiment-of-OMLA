

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731;

  XNOR2_X1 U373 ( .A(n720), .B(G146), .ZN(n397) );
  XNOR2_X1 U374 ( .A(G110), .B(G107), .ZN(n370) );
  NOR2_X1 U375 ( .A1(n527), .A2(n526), .ZN(n529) );
  XNOR2_X1 U376 ( .A(n649), .B(KEYINPUT2), .ZN(n584) );
  NAND2_X2 U377 ( .A1(n486), .A2(n350), .ZN(n488) );
  INV_X1 U378 ( .A(n670), .ZN(n399) );
  NOR2_X2 U379 ( .A1(n559), .A2(n475), .ZN(n386) );
  OR2_X2 U380 ( .A1(n615), .A2(G902), .ZN(n378) );
  AND2_X2 U381 ( .A1(n584), .A2(n583), .ZN(n625) );
  AND2_X1 U382 ( .A1(n664), .A2(n665), .ZN(n562) );
  NOR2_X2 U383 ( .A1(n623), .A2(KEYINPUT44), .ZN(n542) );
  XNOR2_X2 U384 ( .A(n540), .B(KEYINPUT35), .ZN(n623) );
  XNOR2_X2 U385 ( .A(n471), .B(KEYINPUT39), .ZN(n486) );
  XNOR2_X1 U386 ( .A(n534), .B(KEYINPUT33), .ZN(n686) );
  XNOR2_X1 U387 ( .A(n653), .B(n652), .ZN(n654) );
  NAND2_X1 U388 ( .A1(n686), .A2(n560), .ZN(n536) );
  INV_X1 U389 ( .A(KEYINPUT34), .ZN(n535) );
  XNOR2_X1 U390 ( .A(n380), .B(n379), .ZN(n559) );
  INV_X1 U391 ( .A(KEYINPUT95), .ZN(n379) );
  NOR2_X1 U392 ( .A1(n474), .A2(n473), .ZN(n350) );
  AND2_X1 U393 ( .A1(n366), .A2(G217), .ZN(n351) );
  XNOR2_X1 U394 ( .A(KEYINPUT107), .B(KEYINPUT30), .ZN(n352) );
  XNOR2_X1 U395 ( .A(KEYINPUT15), .B(G902), .ZN(n582) );
  INV_X1 U396 ( .A(KEYINPUT86), .ZN(n551) );
  INV_X1 U397 ( .A(G104), .ZN(n372) );
  XNOR2_X1 U398 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U399 ( .A(n718), .B(n374), .ZN(n375) );
  INV_X1 U400 ( .A(KEYINPUT85), .ZN(n652) );
  INV_X1 U401 ( .A(KEYINPUT48), .ZN(n528) );
  INV_X1 U402 ( .A(KEYINPUT84), .ZN(n657) );
  AND2_X1 U403 ( .A1(n543), .A2(n661), .ZN(n665) );
  OR2_X1 U404 ( .A1(n590), .A2(G902), .ZN(n398) );
  XNOR2_X1 U405 ( .A(n529), .B(n528), .ZN(n533) );
  BUF_X1 U406 ( .A(n686), .Z(n698) );
  INV_X1 U407 ( .A(n582), .ZN(n583) );
  OR2_X1 U408 ( .A1(n600), .A2(n583), .ZN(n451) );
  XNOR2_X1 U409 ( .A(n536), .B(n535), .ZN(n539) );
  XNOR2_X1 U410 ( .A(n405), .B(KEYINPUT77), .ZN(n470) );
  NOR2_X1 U411 ( .A1(n703), .A2(G953), .ZN(n704) );
  XOR2_X1 U412 ( .A(KEYINPUT70), .B(KEYINPUT8), .Z(n354) );
  INV_X2 U413 ( .A(G953), .ZN(n725) );
  NAND2_X1 U414 ( .A1(G234), .A2(n725), .ZN(n353) );
  XNOR2_X1 U415 ( .A(n354), .B(n353), .ZN(n424) );
  NAND2_X1 U416 ( .A1(G221), .A2(n424), .ZN(n355) );
  XNOR2_X1 U417 ( .A(G146), .B(G125), .ZN(n440) );
  XNOR2_X1 U418 ( .A(n440), .B(KEYINPUT10), .ZN(n717) );
  XNOR2_X1 U419 ( .A(n355), .B(n717), .ZN(n362) );
  XNOR2_X1 U420 ( .A(G119), .B(G110), .ZN(n356) );
  XNOR2_X1 U421 ( .A(G137), .B(G140), .ZN(n371) );
  XNOR2_X1 U422 ( .A(n356), .B(n371), .ZN(n360) );
  XOR2_X1 U423 ( .A(KEYINPUT94), .B(KEYINPUT23), .Z(n358) );
  XNOR2_X1 U424 ( .A(G128), .B(KEYINPUT24), .ZN(n357) );
  XNOR2_X1 U425 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U426 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U427 ( .A(n362), .B(n361), .ZN(n586) );
  INV_X1 U428 ( .A(G902), .ZN(n401) );
  NAND2_X1 U429 ( .A1(n586), .A2(n401), .ZN(n365) );
  NAND2_X1 U430 ( .A1(G234), .A2(n582), .ZN(n363) );
  XNOR2_X1 U431 ( .A(n363), .B(KEYINPUT20), .ZN(n366) );
  XNOR2_X1 U432 ( .A(KEYINPUT25), .B(n351), .ZN(n364) );
  XNOR2_X2 U433 ( .A(n365), .B(n364), .ZN(n543) );
  AND2_X1 U434 ( .A1(n366), .A2(G221), .ZN(n367) );
  XNOR2_X1 U435 ( .A(n367), .B(KEYINPUT21), .ZN(n661) );
  XNOR2_X1 U436 ( .A(KEYINPUT71), .B(G131), .ZN(n412) );
  XNOR2_X1 U437 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n442) );
  XNOR2_X1 U438 ( .A(n412), .B(n442), .ZN(n369) );
  XNOR2_X2 U439 ( .A(G143), .B(G128), .ZN(n443) );
  INV_X1 U440 ( .A(G134), .ZN(n368) );
  XNOR2_X1 U441 ( .A(n443), .B(n368), .ZN(n422) );
  XNOR2_X1 U442 ( .A(n369), .B(n422), .ZN(n720) );
  XNOR2_X1 U443 ( .A(n370), .B(G101), .ZN(n432) );
  XNOR2_X1 U444 ( .A(KEYINPUT93), .B(n371), .ZN(n718) );
  NAND2_X1 U445 ( .A1(G227), .A2(n725), .ZN(n373) );
  XNOR2_X1 U446 ( .A(n432), .B(n375), .ZN(n376) );
  XNOR2_X1 U447 ( .A(n397), .B(n376), .ZN(n615) );
  XOR2_X1 U448 ( .A(KEYINPUT73), .B(G469), .Z(n377) );
  XNOR2_X2 U449 ( .A(n378), .B(n377), .ZN(n493) );
  NAND2_X1 U450 ( .A1(n665), .A2(n493), .ZN(n380) );
  NAND2_X1 U451 ( .A1(G234), .A2(G237), .ZN(n381) );
  XNOR2_X1 U452 ( .A(n381), .B(KEYINPUT14), .ZN(n382) );
  NAND2_X1 U453 ( .A1(G952), .A2(n382), .ZN(n694) );
  NOR2_X1 U454 ( .A1(G953), .A2(n694), .ZN(n458) );
  AND2_X1 U455 ( .A1(G953), .A2(n382), .ZN(n383) );
  NAND2_X1 U456 ( .A1(G902), .A2(n383), .ZN(n456) );
  XNOR2_X1 U457 ( .A(KEYINPUT106), .B(n456), .ZN(n384) );
  NOR2_X1 U458 ( .A1(G900), .A2(n384), .ZN(n385) );
  NOR2_X1 U459 ( .A1(n458), .A2(n385), .ZN(n475) );
  XNOR2_X1 U460 ( .A(n386), .B(KEYINPUT78), .ZN(n404) );
  XNOR2_X1 U461 ( .A(G119), .B(G116), .ZN(n388) );
  XNOR2_X1 U462 ( .A(KEYINPUT74), .B(KEYINPUT3), .ZN(n387) );
  XNOR2_X1 U463 ( .A(n388), .B(n387), .ZN(n435) );
  XNOR2_X1 U464 ( .A(G101), .B(G113), .ZN(n389) );
  XNOR2_X1 U465 ( .A(n389), .B(KEYINPUT96), .ZN(n390) );
  XNOR2_X1 U466 ( .A(n435), .B(n390), .ZN(n395) );
  NOR2_X1 U467 ( .A1(G237), .A2(G953), .ZN(n391) );
  XNOR2_X1 U468 ( .A(KEYINPUT76), .B(n391), .ZN(n408) );
  AND2_X1 U469 ( .A1(n408), .A2(G210), .ZN(n393) );
  XNOR2_X1 U470 ( .A(KEYINPUT5), .B(G137), .ZN(n392) );
  XNOR2_X1 U471 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U472 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U473 ( .A(n397), .B(n396), .ZN(n590) );
  XNOR2_X2 U474 ( .A(n398), .B(G472), .ZN(n670) );
  XNOR2_X2 U475 ( .A(n399), .B(KEYINPUT105), .ZN(n491) );
  INV_X1 U476 ( .A(G237), .ZN(n400) );
  NAND2_X1 U477 ( .A1(n401), .A2(n400), .ZN(n447) );
  AND2_X1 U478 ( .A1(n447), .A2(G214), .ZN(n453) );
  INV_X1 U479 ( .A(n453), .ZN(n677) );
  NAND2_X1 U480 ( .A1(n491), .A2(n677), .ZN(n402) );
  XNOR2_X1 U481 ( .A(n402), .B(n352), .ZN(n403) );
  NAND2_X1 U482 ( .A1(n404), .A2(n403), .ZN(n405) );
  XNOR2_X1 U483 ( .A(KEYINPUT99), .B(KEYINPUT13), .ZN(n418) );
  XOR2_X1 U484 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n407) );
  XNOR2_X1 U485 ( .A(G143), .B(G140), .ZN(n406) );
  XNOR2_X1 U486 ( .A(n407), .B(n406), .ZN(n410) );
  NAND2_X1 U487 ( .A1(n408), .A2(G214), .ZN(n409) );
  XNOR2_X1 U488 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U489 ( .A(n411), .B(n717), .ZN(n416) );
  XOR2_X1 U490 ( .A(KEYINPUT98), .B(n412), .Z(n414) );
  XNOR2_X1 U491 ( .A(G122), .B(G113), .ZN(n413) );
  XNOR2_X1 U492 ( .A(n413), .B(G104), .ZN(n434) );
  XNOR2_X1 U493 ( .A(n414), .B(n434), .ZN(n415) );
  XNOR2_X1 U494 ( .A(n416), .B(n415), .ZN(n609) );
  NOR2_X1 U495 ( .A1(G902), .A2(n609), .ZN(n417) );
  XNOR2_X1 U496 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U497 ( .A(n419), .B(G475), .ZN(n474) );
  XOR2_X1 U498 ( .A(KEYINPUT100), .B(G122), .Z(n421) );
  XNOR2_X1 U499 ( .A(G116), .B(G107), .ZN(n420) );
  XNOR2_X1 U500 ( .A(n421), .B(n420), .ZN(n423) );
  XNOR2_X1 U501 ( .A(n423), .B(n422), .ZN(n428) );
  NAND2_X1 U502 ( .A1(G217), .A2(n424), .ZN(n426) );
  XNOR2_X1 U503 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n425) );
  XNOR2_X1 U504 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U505 ( .A(n428), .B(n427), .ZN(n626) );
  NOR2_X1 U506 ( .A1(G902), .A2(n626), .ZN(n429) );
  XNOR2_X1 U507 ( .A(n429), .B(KEYINPUT101), .ZN(n431) );
  INV_X1 U508 ( .A(G478), .ZN(n430) );
  XNOR2_X1 U509 ( .A(n431), .B(n430), .ZN(n472) );
  OR2_X1 U510 ( .A1(n474), .A2(n472), .ZN(n537) );
  INV_X1 U511 ( .A(n432), .ZN(n433) );
  XNOR2_X1 U512 ( .A(n433), .B(KEYINPUT16), .ZN(n437) );
  XNOR2_X1 U513 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U514 ( .A(n437), .B(n436), .ZN(n712) );
  XNOR2_X1 U515 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n439) );
  NAND2_X1 U516 ( .A1(n725), .A2(G224), .ZN(n438) );
  XNOR2_X1 U517 ( .A(n439), .B(n438), .ZN(n441) );
  XNOR2_X1 U518 ( .A(n441), .B(n440), .ZN(n445) );
  XNOR2_X1 U519 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U520 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U521 ( .A(n712), .B(n446), .ZN(n600) );
  NAND2_X1 U522 ( .A1(n447), .A2(G210), .ZN(n449) );
  INV_X1 U523 ( .A(KEYINPUT91), .ZN(n448) );
  XNOR2_X1 U524 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X2 U525 ( .A(n451), .B(n450), .ZN(n484) );
  NOR2_X1 U526 ( .A1(n537), .A2(n484), .ZN(n452) );
  NAND2_X1 U527 ( .A1(n470), .A2(n452), .ZN(n525) );
  XNOR2_X1 U528 ( .A(n525), .B(G143), .ZN(G45) );
  OR2_X2 U529 ( .A1(n484), .A2(n453), .ZN(n499) );
  XNOR2_X1 U530 ( .A(KEYINPUT79), .B(KEYINPUT19), .ZN(n454) );
  XNOR2_X1 U531 ( .A(n454), .B(KEYINPUT67), .ZN(n455) );
  XNOR2_X2 U532 ( .A(n499), .B(n455), .ZN(n506) );
  NOR2_X1 U533 ( .A1(G898), .A2(n456), .ZN(n457) );
  OR2_X1 U534 ( .A1(n458), .A2(n457), .ZN(n459) );
  XNOR2_X1 U535 ( .A(n459), .B(KEYINPUT92), .ZN(n460) );
  NAND2_X1 U536 ( .A1(n506), .A2(n460), .ZN(n461) );
  XNOR2_X1 U537 ( .A(n461), .B(KEYINPUT0), .ZN(n563) );
  NAND2_X1 U538 ( .A1(n474), .A2(n472), .ZN(n680) );
  INV_X1 U539 ( .A(n661), .ZN(n476) );
  OR2_X1 U540 ( .A1(n680), .A2(n476), .ZN(n462) );
  OR2_X2 U541 ( .A1(n563), .A2(n462), .ZN(n465) );
  INV_X1 U542 ( .A(KEYINPUT66), .ZN(n463) );
  XNOR2_X1 U543 ( .A(n463), .B(KEYINPUT22), .ZN(n464) );
  XNOR2_X2 U544 ( .A(n465), .B(n464), .ZN(n567) );
  INV_X1 U545 ( .A(n491), .ZN(n467) );
  INV_X1 U546 ( .A(n543), .ZN(n466) );
  NAND2_X1 U547 ( .A1(n467), .A2(n466), .ZN(n468) );
  XNOR2_X2 U548 ( .A(n493), .B(KEYINPUT1), .ZN(n664) );
  NOR2_X1 U549 ( .A1(n468), .A2(n664), .ZN(n469) );
  NAND2_X1 U550 ( .A1(n567), .A2(n469), .ZN(n550) );
  XNOR2_X1 U551 ( .A(n550), .B(G110), .ZN(G12) );
  XNOR2_X1 U552 ( .A(n484), .B(KEYINPUT38), .ZN(n678) );
  NAND2_X1 U553 ( .A1(n470), .A2(n678), .ZN(n471) );
  INV_X1 U554 ( .A(n472), .ZN(n473) );
  AND2_X1 U555 ( .A1(n474), .A2(n473), .ZN(n644) );
  NAND2_X1 U556 ( .A1(n486), .A2(n644), .ZN(n531) );
  XNOR2_X1 U557 ( .A(n531), .B(G134), .ZN(G36) );
  NOR2_X1 U558 ( .A1(n476), .A2(n475), .ZN(n477) );
  XOR2_X1 U559 ( .A(KEYINPUT72), .B(n477), .Z(n478) );
  NOR2_X1 U560 ( .A1(n478), .A2(n543), .ZN(n490) );
  AND2_X1 U561 ( .A1(n350), .A2(n490), .ZN(n480) );
  XNOR2_X1 U562 ( .A(KEYINPUT103), .B(KEYINPUT6), .ZN(n479) );
  XNOR2_X1 U563 ( .A(n670), .B(n479), .ZN(n569) );
  NAND2_X1 U564 ( .A1(n480), .A2(n569), .ZN(n500) );
  NOR2_X1 U565 ( .A1(n664), .A2(n500), .ZN(n481) );
  NAND2_X1 U566 ( .A1(n677), .A2(n481), .ZN(n482) );
  XNOR2_X1 U567 ( .A(n482), .B(KEYINPUT43), .ZN(n483) );
  NAND2_X1 U568 ( .A1(n484), .A2(n483), .ZN(n530) );
  XNOR2_X1 U569 ( .A(G140), .B(KEYINPUT114), .ZN(n485) );
  XNOR2_X1 U570 ( .A(n530), .B(n485), .ZN(G42) );
  XNOR2_X1 U571 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n487) );
  XNOR2_X2 U572 ( .A(n488), .B(n487), .ZN(n624) );
  NAND2_X1 U573 ( .A1(n678), .A2(n677), .ZN(n682) );
  NOR2_X1 U574 ( .A1(n680), .A2(n682), .ZN(n489) );
  XNOR2_X1 U575 ( .A(n489), .B(KEYINPUT41), .ZN(n697) );
  NAND2_X1 U576 ( .A1(n491), .A2(n490), .ZN(n492) );
  XNOR2_X1 U577 ( .A(n492), .B(KEYINPUT28), .ZN(n495) );
  INV_X1 U578 ( .A(n493), .ZN(n494) );
  OR2_X1 U579 ( .A1(n495), .A2(n494), .ZN(n508) );
  NOR2_X1 U580 ( .A1(n697), .A2(n508), .ZN(n497) );
  XNOR2_X1 U581 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n496) );
  XNOR2_X1 U582 ( .A(n497), .B(n496), .ZN(n730) );
  NAND2_X1 U583 ( .A1(n624), .A2(n730), .ZN(n498) );
  XNOR2_X1 U584 ( .A(n498), .B(KEYINPUT46), .ZN(n527) );
  XNOR2_X1 U585 ( .A(n664), .B(KEYINPUT90), .ZN(n546) );
  NOR2_X1 U586 ( .A1(n500), .A2(n499), .ZN(n502) );
  XNOR2_X1 U587 ( .A(KEYINPUT110), .B(KEYINPUT36), .ZN(n501) );
  XNOR2_X1 U588 ( .A(n502), .B(n501), .ZN(n503) );
  NAND2_X1 U589 ( .A1(n546), .A2(n503), .ZN(n648) );
  NOR2_X1 U590 ( .A1(n644), .A2(n350), .ZN(n504) );
  XNOR2_X1 U591 ( .A(n504), .B(KEYINPUT102), .ZN(n681) );
  INV_X1 U592 ( .A(n681), .ZN(n516) );
  NAND2_X1 U593 ( .A1(n516), .A2(KEYINPUT83), .ZN(n505) );
  NAND2_X1 U594 ( .A1(n648), .A2(n505), .ZN(n510) );
  INV_X1 U595 ( .A(n506), .ZN(n507) );
  OR2_X1 U596 ( .A1(n508), .A2(n507), .ZN(n514) );
  NOR2_X1 U597 ( .A1(n514), .A2(KEYINPUT82), .ZN(n509) );
  OR2_X1 U598 ( .A1(n510), .A2(n509), .ZN(n523) );
  NOR2_X1 U599 ( .A1(n681), .A2(n514), .ZN(n513) );
  NOR2_X1 U600 ( .A1(KEYINPUT83), .A2(KEYINPUT47), .ZN(n511) );
  NAND2_X1 U601 ( .A1(n511), .A2(KEYINPUT82), .ZN(n512) );
  NOR2_X1 U602 ( .A1(n513), .A2(n512), .ZN(n521) );
  INV_X1 U603 ( .A(n514), .ZN(n641) );
  INV_X1 U604 ( .A(KEYINPUT82), .ZN(n515) );
  NOR2_X1 U605 ( .A1(n641), .A2(n515), .ZN(n519) );
  OR2_X1 U606 ( .A1(KEYINPUT83), .A2(n516), .ZN(n517) );
  NAND2_X1 U607 ( .A1(KEYINPUT47), .A2(n517), .ZN(n518) );
  NOR2_X1 U608 ( .A1(n519), .A2(n518), .ZN(n520) );
  NOR2_X1 U609 ( .A1(n521), .A2(n520), .ZN(n522) );
  NOR2_X1 U610 ( .A1(n523), .A2(n522), .ZN(n524) );
  NAND2_X1 U611 ( .A1(n525), .A2(n524), .ZN(n526) );
  NAND2_X1 U612 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X2 U613 ( .A1(n533), .A2(n532), .ZN(n721) );
  NAND2_X1 U614 ( .A1(n562), .A2(n569), .ZN(n534) );
  INV_X1 U615 ( .A(n563), .ZN(n560) );
  INV_X1 U616 ( .A(n537), .ZN(n538) );
  NAND2_X1 U617 ( .A1(n539), .A2(n538), .ZN(n540) );
  INV_X1 U618 ( .A(KEYINPUT69), .ZN(n541) );
  XNOR2_X1 U619 ( .A(n542), .B(n541), .ZN(n553) );
  INV_X1 U620 ( .A(n569), .ZN(n544) );
  XNOR2_X1 U621 ( .A(n543), .B(KEYINPUT104), .ZN(n662) );
  INV_X1 U622 ( .A(n662), .ZN(n568) );
  AND2_X1 U623 ( .A1(n544), .A2(n568), .ZN(n545) );
  AND2_X1 U624 ( .A1(n546), .A2(n545), .ZN(n547) );
  NAND2_X1 U625 ( .A1(n567), .A2(n547), .ZN(n549) );
  XNOR2_X1 U626 ( .A(KEYINPUT80), .B(KEYINPUT32), .ZN(n548) );
  XNOR2_X1 U627 ( .A(n549), .B(n548), .ZN(n607) );
  NAND2_X1 U628 ( .A1(n607), .A2(n550), .ZN(n555) );
  XNOR2_X1 U629 ( .A(n555), .B(n551), .ZN(n552) );
  NAND2_X1 U630 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U631 ( .A(n554), .B(KEYINPUT75), .ZN(n578) );
  INV_X1 U632 ( .A(n623), .ZN(n557) );
  INV_X1 U633 ( .A(n555), .ZN(n556) );
  NAND2_X1 U634 ( .A1(n557), .A2(n556), .ZN(n558) );
  NAND2_X1 U635 ( .A1(n558), .A2(KEYINPUT44), .ZN(n576) );
  NOR2_X1 U636 ( .A1(n559), .A2(n670), .ZN(n561) );
  AND2_X1 U637 ( .A1(n561), .A2(n560), .ZN(n634) );
  NAND2_X1 U638 ( .A1(n562), .A2(n670), .ZN(n672) );
  OR2_X1 U639 ( .A1(n563), .A2(n672), .ZN(n565) );
  XOR2_X1 U640 ( .A(KEYINPUT97), .B(KEYINPUT31), .Z(n564) );
  XNOR2_X1 U641 ( .A(n565), .B(n564), .ZN(n645) );
  NOR2_X1 U642 ( .A1(n634), .A2(n645), .ZN(n566) );
  NOR2_X1 U643 ( .A1(n566), .A2(n681), .ZN(n574) );
  INV_X1 U644 ( .A(n567), .ZN(n573) );
  NOR2_X1 U645 ( .A1(n569), .A2(n568), .ZN(n571) );
  INV_X1 U646 ( .A(n664), .ZN(n570) );
  NAND2_X1 U647 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U648 ( .A1(n573), .A2(n572), .ZN(n630) );
  NOR2_X1 U649 ( .A1(n574), .A2(n630), .ZN(n575) );
  NAND2_X1 U650 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X2 U651 ( .A1(n578), .A2(n577), .ZN(n580) );
  XOR2_X1 U652 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n579) );
  XNOR2_X1 U653 ( .A(n580), .B(n579), .ZN(n656) );
  NAND2_X1 U654 ( .A1(n721), .A2(n656), .ZN(n649) );
  INV_X1 U655 ( .A(KEYINPUT2), .ZN(n581) );
  NAND2_X1 U656 ( .A1(n625), .A2(G217), .ZN(n585) );
  XOR2_X1 U657 ( .A(n586), .B(n585), .Z(n588) );
  INV_X1 U658 ( .A(G952), .ZN(n587) );
  NAND2_X1 U659 ( .A1(n587), .A2(G953), .ZN(n619) );
  INV_X1 U660 ( .A(n619), .ZN(n628) );
  NOR2_X1 U661 ( .A1(n588), .A2(n628), .ZN(G66) );
  NAND2_X1 U662 ( .A1(n625), .A2(G472), .ZN(n592) );
  XNOR2_X1 U663 ( .A(KEYINPUT89), .B(KEYINPUT62), .ZN(n589) );
  XNOR2_X1 U664 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U665 ( .A(n592), .B(n591), .ZN(n593) );
  NAND2_X1 U666 ( .A1(n593), .A2(n619), .ZN(n594) );
  XNOR2_X1 U667 ( .A(n594), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U668 ( .A1(n625), .A2(G210), .ZN(n602) );
  XOR2_X1 U669 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n596) );
  XNOR2_X1 U670 ( .A(KEYINPUT55), .B(KEYINPUT81), .ZN(n595) );
  XNOR2_X1 U671 ( .A(n596), .B(n595), .ZN(n598) );
  XNOR2_X1 U672 ( .A(KEYINPUT119), .B(KEYINPUT54), .ZN(n597) );
  XNOR2_X1 U673 ( .A(n598), .B(n597), .ZN(n599) );
  XNOR2_X1 U674 ( .A(n600), .B(n599), .ZN(n601) );
  XNOR2_X1 U675 ( .A(n602), .B(n601), .ZN(n603) );
  NAND2_X1 U676 ( .A1(n603), .A2(n619), .ZN(n605) );
  INV_X1 U677 ( .A(KEYINPUT56), .ZN(n604) );
  XNOR2_X1 U678 ( .A(n605), .B(n604), .ZN(G51) );
  XNOR2_X1 U679 ( .A(G119), .B(KEYINPUT126), .ZN(n606) );
  XNOR2_X1 U680 ( .A(n607), .B(n606), .ZN(G21) );
  NAND2_X1 U681 ( .A1(n625), .A2(G475), .ZN(n611) );
  XOR2_X1 U682 ( .A(KEYINPUT121), .B(KEYINPUT59), .Z(n608) );
  XNOR2_X1 U683 ( .A(n609), .B(n608), .ZN(n610) );
  XNOR2_X1 U684 ( .A(n611), .B(n610), .ZN(n612) );
  NAND2_X1 U685 ( .A1(n612), .A2(n619), .ZN(n614) );
  XOR2_X1 U686 ( .A(KEYINPUT68), .B(KEYINPUT60), .Z(n613) );
  XNOR2_X1 U687 ( .A(n614), .B(n613), .ZN(G60) );
  NAND2_X1 U688 ( .A1(n625), .A2(G469), .ZN(n618) );
  XNOR2_X1 U689 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n616) );
  XNOR2_X1 U690 ( .A(n615), .B(n616), .ZN(n617) );
  XNOR2_X1 U691 ( .A(n618), .B(n617), .ZN(n620) );
  NAND2_X1 U692 ( .A1(n620), .A2(n619), .ZN(n622) );
  INV_X1 U693 ( .A(KEYINPUT120), .ZN(n621) );
  XNOR2_X1 U694 ( .A(n622), .B(n621), .ZN(G54) );
  XOR2_X1 U695 ( .A(n623), .B(G122), .Z(G24) );
  XNOR2_X1 U696 ( .A(n624), .B(G131), .ZN(G33) );
  NAND2_X1 U697 ( .A1(n625), .A2(G478), .ZN(n627) );
  XNOR2_X1 U698 ( .A(n627), .B(n626), .ZN(n629) );
  NOR2_X1 U699 ( .A1(n629), .A2(n628), .ZN(G63) );
  XNOR2_X1 U700 ( .A(n630), .B(G101), .ZN(n631) );
  XNOR2_X1 U701 ( .A(n631), .B(KEYINPUT111), .ZN(G3) );
  NAND2_X1 U702 ( .A1(n634), .A2(n350), .ZN(n632) );
  XNOR2_X1 U703 ( .A(n632), .B(KEYINPUT112), .ZN(n633) );
  XNOR2_X1 U704 ( .A(G104), .B(n633), .ZN(G6) );
  XOR2_X1 U705 ( .A(KEYINPUT26), .B(KEYINPUT113), .Z(n636) );
  NAND2_X1 U706 ( .A1(n634), .A2(n644), .ZN(n635) );
  XNOR2_X1 U707 ( .A(n636), .B(n635), .ZN(n638) );
  XOR2_X1 U708 ( .A(G107), .B(KEYINPUT27), .Z(n637) );
  XNOR2_X1 U709 ( .A(n638), .B(n637), .ZN(G9) );
  XOR2_X1 U710 ( .A(G128), .B(KEYINPUT29), .Z(n640) );
  NAND2_X1 U711 ( .A1(n641), .A2(n644), .ZN(n639) );
  XNOR2_X1 U712 ( .A(n640), .B(n639), .ZN(G30) );
  NAND2_X1 U713 ( .A1(n641), .A2(n350), .ZN(n642) );
  XNOR2_X1 U714 ( .A(n642), .B(G146), .ZN(G48) );
  NAND2_X1 U715 ( .A1(n645), .A2(n350), .ZN(n643) );
  XNOR2_X1 U716 ( .A(n643), .B(G113), .ZN(G15) );
  NAND2_X1 U717 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U718 ( .A(n646), .B(G116), .ZN(G18) );
  XOR2_X1 U719 ( .A(G125), .B(KEYINPUT37), .Z(n647) );
  XNOR2_X1 U720 ( .A(n648), .B(n647), .ZN(G27) );
  INV_X1 U721 ( .A(n649), .ZN(n650) );
  NAND2_X1 U722 ( .A1(n650), .A2(KEYINPUT2), .ZN(n655) );
  INV_X1 U723 ( .A(n721), .ZN(n651) );
  NAND2_X1 U724 ( .A1(n651), .A2(n581), .ZN(n653) );
  NAND2_X1 U725 ( .A1(n655), .A2(n654), .ZN(n660) );
  INV_X1 U726 ( .A(n656), .ZN(n705) );
  NAND2_X1 U727 ( .A1(n705), .A2(n581), .ZN(n658) );
  XNOR2_X1 U728 ( .A(n658), .B(n657), .ZN(n659) );
  NOR2_X1 U729 ( .A1(n660), .A2(n659), .ZN(n696) );
  NOR2_X1 U730 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U731 ( .A(KEYINPUT49), .B(n663), .ZN(n669) );
  NOR2_X1 U732 ( .A1(n665), .A2(n664), .ZN(n667) );
  XNOR2_X1 U733 ( .A(KEYINPUT115), .B(KEYINPUT50), .ZN(n666) );
  XNOR2_X1 U734 ( .A(n667), .B(n666), .ZN(n668) );
  NAND2_X1 U735 ( .A1(n669), .A2(n668), .ZN(n671) );
  NOR2_X1 U736 ( .A1(n671), .A2(n670), .ZN(n674) );
  INV_X1 U737 ( .A(n672), .ZN(n673) );
  NOR2_X1 U738 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U739 ( .A(KEYINPUT51), .B(n675), .Z(n676) );
  NOR2_X1 U740 ( .A1(n697), .A2(n676), .ZN(n690) );
  NOR2_X1 U741 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U742 ( .A1(n680), .A2(n679), .ZN(n685) );
  NOR2_X1 U743 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U744 ( .A(n683), .B(KEYINPUT116), .ZN(n684) );
  NOR2_X1 U745 ( .A1(n685), .A2(n684), .ZN(n688) );
  INV_X1 U746 ( .A(n698), .ZN(n687) );
  NOR2_X1 U747 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U748 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U749 ( .A(n691), .B(KEYINPUT52), .Z(n692) );
  XNOR2_X1 U750 ( .A(KEYINPUT117), .B(n692), .ZN(n693) );
  NOR2_X1 U751 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U752 ( .A1(n696), .A2(n695), .ZN(n702) );
  INV_X1 U753 ( .A(n697), .ZN(n699) );
  NAND2_X1 U754 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U755 ( .A(n700), .B(KEYINPUT118), .ZN(n701) );
  NAND2_X1 U756 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U757 ( .A(n704), .B(KEYINPUT53), .ZN(G75) );
  NOR2_X1 U758 ( .A1(n705), .A2(G953), .ZN(n711) );
  NAND2_X1 U759 ( .A1(G224), .A2(G953), .ZN(n706) );
  XNOR2_X1 U760 ( .A(n706), .B(KEYINPUT122), .ZN(n707) );
  XNOR2_X1 U761 ( .A(KEYINPUT61), .B(n707), .ZN(n708) );
  NAND2_X1 U762 ( .A1(n708), .A2(G898), .ZN(n709) );
  XNOR2_X1 U763 ( .A(n709), .B(KEYINPUT123), .ZN(n710) );
  NOR2_X1 U764 ( .A1(n711), .A2(n710), .ZN(n716) );
  XOR2_X1 U765 ( .A(KEYINPUT124), .B(n712), .Z(n714) );
  NOR2_X1 U766 ( .A1(n725), .A2(G898), .ZN(n713) );
  NOR2_X1 U767 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U768 ( .A(n716), .B(n715), .Z(G69) );
  XNOR2_X1 U769 ( .A(n718), .B(n717), .ZN(n719) );
  XOR2_X1 U770 ( .A(n720), .B(n719), .Z(n723) );
  XNOR2_X1 U771 ( .A(n721), .B(n723), .ZN(n722) );
  NAND2_X1 U772 ( .A1(n722), .A2(n725), .ZN(n728) );
  XOR2_X1 U773 ( .A(n723), .B(G227), .Z(n724) );
  NOR2_X1 U774 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U775 ( .A1(G900), .A2(n726), .ZN(n727) );
  NAND2_X1 U776 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U777 ( .A(KEYINPUT125), .B(n729), .ZN(G72) );
  XOR2_X1 U778 ( .A(G137), .B(n730), .Z(n731) );
  XNOR2_X1 U779 ( .A(KEYINPUT127), .B(n731), .ZN(G39) );
endmodule

