

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X2 U548 ( .A(n722), .Z(n513) );
  BUF_X1 U549 ( .A(n691), .Z(n722) );
  AND2_X2 U550 ( .A1(n519), .A2(G2104), .ZN(n879) );
  NOR2_X2 U551 ( .A1(G2104), .A2(G2105), .ZN(n516) );
  NOR2_X2 U552 ( .A1(G1384), .A2(G164), .ZN(n743) );
  AND2_X1 U553 ( .A1(n729), .A2(n728), .ZN(n730) );
  INV_X1 U554 ( .A(KEYINPUT17), .ZN(n515) );
  NAND2_X1 U555 ( .A1(n743), .A2(n677), .ZN(n691) );
  XNOR2_X2 U556 ( .A(n730), .B(KEYINPUT32), .ZN(n784) );
  NAND2_X1 U557 ( .A1(n880), .A2(G137), .ZN(n517) );
  AND2_X1 U558 ( .A1(n521), .A2(n520), .ZN(n514) );
  INV_X1 U559 ( .A(KEYINPUT26), .ZN(n692) );
  NOR2_X1 U560 ( .A1(n696), .A2(n974), .ZN(n697) );
  AND2_X1 U561 ( .A1(n733), .A2(n732), .ZN(n736) );
  NOR2_X1 U562 ( .A1(G651), .A2(n623), .ZN(n644) );
  AND2_X1 U563 ( .A1(n522), .A2(n514), .ZN(n523) );
  XNOR2_X2 U564 ( .A(n516), .B(n515), .ZN(n880) );
  XOR2_X1 U565 ( .A(KEYINPUT65), .B(n517), .Z(n524) );
  INV_X1 U566 ( .A(G2105), .ZN(n519) );
  NAND2_X1 U567 ( .A1(G101), .A2(n879), .ZN(n518) );
  XOR2_X1 U568 ( .A(KEYINPUT23), .B(n518), .Z(n522) );
  NOR2_X2 U569 ( .A1(G2104), .A2(n519), .ZN(n875) );
  NAND2_X1 U570 ( .A1(G125), .A2(n875), .ZN(n521) );
  AND2_X1 U571 ( .A1(G2104), .A2(G2105), .ZN(n876) );
  NAND2_X1 U572 ( .A1(G113), .A2(n876), .ZN(n520) );
  AND2_X2 U573 ( .A1(n524), .A2(n523), .ZN(G160) );
  NAND2_X1 U574 ( .A1(n876), .A2(G114), .ZN(n531) );
  NAND2_X1 U575 ( .A1(G126), .A2(n875), .ZN(n526) );
  NAND2_X1 U576 ( .A1(G138), .A2(n880), .ZN(n525) );
  NAND2_X1 U577 ( .A1(n526), .A2(n525), .ZN(n529) );
  NAND2_X1 U578 ( .A1(G102), .A2(n879), .ZN(n527) );
  XNOR2_X1 U579 ( .A(KEYINPUT87), .B(n527), .ZN(n528) );
  NOR2_X1 U580 ( .A1(n529), .A2(n528), .ZN(n530) );
  AND2_X1 U581 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U582 ( .A(KEYINPUT88), .B(n532), .ZN(G164) );
  AND2_X1 U583 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U584 ( .A(G57), .ZN(G237) );
  INV_X1 U585 ( .A(G132), .ZN(G219) );
  NOR2_X1 U586 ( .A1(G651), .A2(G543), .ZN(n640) );
  NAND2_X1 U587 ( .A1(G88), .A2(n640), .ZN(n534) );
  XOR2_X1 U588 ( .A(G543), .B(KEYINPUT0), .Z(n623) );
  INV_X1 U589 ( .A(G651), .ZN(n535) );
  NOR2_X1 U590 ( .A1(n623), .A2(n535), .ZN(n638) );
  NAND2_X1 U591 ( .A1(G75), .A2(n638), .ZN(n533) );
  NAND2_X1 U592 ( .A1(n534), .A2(n533), .ZN(n541) );
  NOR2_X1 U593 ( .A1(G543), .A2(n535), .ZN(n537) );
  XNOR2_X1 U594 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n536) );
  XNOR2_X1 U595 ( .A(n537), .B(n536), .ZN(n641) );
  NAND2_X1 U596 ( .A1(G62), .A2(n641), .ZN(n539) );
  NAND2_X1 U597 ( .A1(G50), .A2(n644), .ZN(n538) );
  NAND2_X1 U598 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U599 ( .A1(n541), .A2(n540), .ZN(G166) );
  XNOR2_X1 U600 ( .A(KEYINPUT7), .B(KEYINPUT78), .ZN(n553) );
  NAND2_X1 U601 ( .A1(n640), .A2(G89), .ZN(n542) );
  XNOR2_X1 U602 ( .A(n542), .B(KEYINPUT4), .ZN(n544) );
  NAND2_X1 U603 ( .A1(G76), .A2(n638), .ZN(n543) );
  NAND2_X1 U604 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U605 ( .A(n545), .B(KEYINPUT5), .ZN(n551) );
  XNOR2_X1 U606 ( .A(KEYINPUT77), .B(KEYINPUT6), .ZN(n549) );
  NAND2_X1 U607 ( .A1(G63), .A2(n641), .ZN(n547) );
  NAND2_X1 U608 ( .A1(G51), .A2(n644), .ZN(n546) );
  NAND2_X1 U609 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U610 ( .A(n549), .B(n548), .ZN(n550) );
  NAND2_X1 U611 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U612 ( .A(n553), .B(n552), .ZN(G168) );
  XOR2_X1 U613 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U614 ( .A1(G7), .A2(G661), .ZN(n554) );
  XNOR2_X1 U615 ( .A(n554), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U616 ( .A(G223), .ZN(n822) );
  NAND2_X1 U617 ( .A1(n822), .A2(G567), .ZN(n555) );
  XNOR2_X1 U618 ( .A(n555), .B(KEYINPUT11), .ZN(n556) );
  XNOR2_X1 U619 ( .A(KEYINPUT71), .B(n556), .ZN(G234) );
  NAND2_X1 U620 ( .A1(G81), .A2(n640), .ZN(n557) );
  XOR2_X1 U621 ( .A(KEYINPUT73), .B(n557), .Z(n558) );
  XNOR2_X1 U622 ( .A(n558), .B(KEYINPUT12), .ZN(n560) );
  NAND2_X1 U623 ( .A1(G68), .A2(n638), .ZN(n559) );
  NAND2_X1 U624 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U625 ( .A(KEYINPUT13), .B(n561), .ZN(n568) );
  XOR2_X1 U626 ( .A(KEYINPUT14), .B(KEYINPUT72), .Z(n563) );
  NAND2_X1 U627 ( .A1(G56), .A2(n641), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(n566) );
  NAND2_X1 U629 ( .A1(G43), .A2(n644), .ZN(n564) );
  XOR2_X1 U630 ( .A(KEYINPUT74), .B(n564), .Z(n565) );
  NOR2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U632 ( .A1(n568), .A2(n567), .ZN(n974) );
  INV_X1 U633 ( .A(G860), .ZN(n615) );
  OR2_X1 U634 ( .A1(n974), .A2(n615), .ZN(G153) );
  NAND2_X1 U635 ( .A1(G90), .A2(n640), .ZN(n570) );
  NAND2_X1 U636 ( .A1(G77), .A2(n638), .ZN(n569) );
  NAND2_X1 U637 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U638 ( .A(KEYINPUT9), .B(n571), .ZN(n575) );
  NAND2_X1 U639 ( .A1(G64), .A2(n641), .ZN(n573) );
  NAND2_X1 U640 ( .A1(G52), .A2(n644), .ZN(n572) );
  AND2_X1 U641 ( .A1(n573), .A2(n572), .ZN(n574) );
  NAND2_X1 U642 ( .A1(n575), .A2(n574), .ZN(G301) );
  NAND2_X1 U643 ( .A1(G868), .A2(G301), .ZN(n586) );
  NAND2_X1 U644 ( .A1(G54), .A2(n644), .ZN(n576) );
  XNOR2_X1 U645 ( .A(n576), .B(KEYINPUT76), .ZN(n583) );
  NAND2_X1 U646 ( .A1(G79), .A2(n638), .ZN(n578) );
  NAND2_X1 U647 ( .A1(G66), .A2(n641), .ZN(n577) );
  NAND2_X1 U648 ( .A1(n578), .A2(n577), .ZN(n581) );
  NAND2_X1 U649 ( .A1(G92), .A2(n640), .ZN(n579) );
  XNOR2_X1 U650 ( .A(KEYINPUT75), .B(n579), .ZN(n580) );
  NOR2_X1 U651 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U652 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U653 ( .A(KEYINPUT15), .B(n584), .ZN(n979) );
  OR2_X1 U654 ( .A1(n979), .A2(G868), .ZN(n585) );
  NAND2_X1 U655 ( .A1(n586), .A2(n585), .ZN(G284) );
  NAND2_X1 U656 ( .A1(G91), .A2(n640), .ZN(n588) );
  NAND2_X1 U657 ( .A1(G78), .A2(n638), .ZN(n587) );
  NAND2_X1 U658 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U659 ( .A1(G53), .A2(n644), .ZN(n589) );
  XNOR2_X1 U660 ( .A(KEYINPUT69), .B(n589), .ZN(n590) );
  NOR2_X1 U661 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U662 ( .A1(n641), .A2(G65), .ZN(n592) );
  NAND2_X1 U663 ( .A1(n593), .A2(n592), .ZN(G299) );
  NAND2_X1 U664 ( .A1(G868), .A2(G286), .ZN(n596) );
  INV_X1 U665 ( .A(G868), .ZN(n594) );
  NAND2_X1 U666 ( .A1(G299), .A2(n594), .ZN(n595) );
  NAND2_X1 U667 ( .A1(n596), .A2(n595), .ZN(G297) );
  NAND2_X1 U668 ( .A1(n615), .A2(G559), .ZN(n597) );
  NAND2_X1 U669 ( .A1(n597), .A2(n979), .ZN(n598) );
  XNOR2_X1 U670 ( .A(n598), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U671 ( .A1(G868), .A2(n974), .ZN(n601) );
  NAND2_X1 U672 ( .A1(G868), .A2(n979), .ZN(n599) );
  NOR2_X1 U673 ( .A1(G559), .A2(n599), .ZN(n600) );
  NOR2_X1 U674 ( .A1(n601), .A2(n600), .ZN(G282) );
  NAND2_X1 U675 ( .A1(G123), .A2(n875), .ZN(n602) );
  XOR2_X1 U676 ( .A(KEYINPUT18), .B(n602), .Z(n603) );
  XNOR2_X1 U677 ( .A(n603), .B(KEYINPUT79), .ZN(n605) );
  NAND2_X1 U678 ( .A1(G111), .A2(n876), .ZN(n604) );
  NAND2_X1 U679 ( .A1(n605), .A2(n604), .ZN(n609) );
  NAND2_X1 U680 ( .A1(G99), .A2(n879), .ZN(n607) );
  NAND2_X1 U681 ( .A1(G135), .A2(n880), .ZN(n606) );
  NAND2_X1 U682 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U683 ( .A1(n609), .A2(n608), .ZN(n610) );
  XOR2_X1 U684 ( .A(KEYINPUT80), .B(n610), .Z(n924) );
  XNOR2_X1 U685 ( .A(n924), .B(G2096), .ZN(n611) );
  XNOR2_X1 U686 ( .A(n611), .B(KEYINPUT81), .ZN(n613) );
  INV_X1 U687 ( .A(G2100), .ZN(n612) );
  NAND2_X1 U688 ( .A1(n613), .A2(n612), .ZN(G156) );
  NAND2_X1 U689 ( .A1(G559), .A2(n979), .ZN(n614) );
  XOR2_X1 U690 ( .A(n974), .B(n614), .Z(n655) );
  NAND2_X1 U691 ( .A1(n615), .A2(n655), .ZN(n622) );
  NAND2_X1 U692 ( .A1(G67), .A2(n641), .ZN(n617) );
  NAND2_X1 U693 ( .A1(G55), .A2(n644), .ZN(n616) );
  NAND2_X1 U694 ( .A1(n617), .A2(n616), .ZN(n621) );
  NAND2_X1 U695 ( .A1(G93), .A2(n640), .ZN(n619) );
  NAND2_X1 U696 ( .A1(G80), .A2(n638), .ZN(n618) );
  NAND2_X1 U697 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U698 ( .A1(n621), .A2(n620), .ZN(n657) );
  XOR2_X1 U699 ( .A(n622), .B(n657), .Z(G145) );
  NAND2_X1 U700 ( .A1(G87), .A2(n623), .ZN(n624) );
  XNOR2_X1 U701 ( .A(n624), .B(KEYINPUT82), .ZN(n629) );
  NAND2_X1 U702 ( .A1(G49), .A2(n644), .ZN(n626) );
  NAND2_X1 U703 ( .A1(G74), .A2(G651), .ZN(n625) );
  NAND2_X1 U704 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U705 ( .A1(n641), .A2(n627), .ZN(n628) );
  NAND2_X1 U706 ( .A1(n629), .A2(n628), .ZN(G288) );
  NAND2_X1 U707 ( .A1(G85), .A2(n640), .ZN(n631) );
  NAND2_X1 U708 ( .A1(G72), .A2(n638), .ZN(n630) );
  NAND2_X1 U709 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U710 ( .A(KEYINPUT66), .B(n632), .Z(n637) );
  NAND2_X1 U711 ( .A1(n644), .A2(G47), .ZN(n634) );
  NAND2_X1 U712 ( .A1(n641), .A2(G60), .ZN(n633) );
  NAND2_X1 U713 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U714 ( .A(KEYINPUT68), .B(n635), .Z(n636) );
  NAND2_X1 U715 ( .A1(n637), .A2(n636), .ZN(G290) );
  NAND2_X1 U716 ( .A1(G73), .A2(n638), .ZN(n639) );
  XNOR2_X1 U717 ( .A(n639), .B(KEYINPUT2), .ZN(n649) );
  NAND2_X1 U718 ( .A1(G86), .A2(n640), .ZN(n643) );
  NAND2_X1 U719 ( .A1(G61), .A2(n641), .ZN(n642) );
  NAND2_X1 U720 ( .A1(n643), .A2(n642), .ZN(n647) );
  NAND2_X1 U721 ( .A1(G48), .A2(n644), .ZN(n645) );
  XNOR2_X1 U722 ( .A(KEYINPUT83), .B(n645), .ZN(n646) );
  NOR2_X1 U723 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U724 ( .A1(n649), .A2(n648), .ZN(G305) );
  XNOR2_X1 U725 ( .A(G166), .B(KEYINPUT19), .ZN(n654) );
  XNOR2_X1 U726 ( .A(n657), .B(G288), .ZN(n652) );
  XNOR2_X1 U727 ( .A(G290), .B(G299), .ZN(n650) );
  XNOR2_X1 U728 ( .A(n650), .B(G305), .ZN(n651) );
  XNOR2_X1 U729 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U730 ( .A(n654), .B(n653), .ZN(n898) );
  XNOR2_X1 U731 ( .A(n655), .B(n898), .ZN(n656) );
  NAND2_X1 U732 ( .A1(n656), .A2(G868), .ZN(n659) );
  OR2_X1 U733 ( .A1(G868), .A2(n657), .ZN(n658) );
  NAND2_X1 U734 ( .A1(n659), .A2(n658), .ZN(G295) );
  NAND2_X1 U735 ( .A1(G2084), .A2(G2078), .ZN(n661) );
  XOR2_X1 U736 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n660) );
  XNOR2_X1 U737 ( .A(n661), .B(n660), .ZN(n662) );
  NAND2_X1 U738 ( .A1(G2090), .A2(n662), .ZN(n663) );
  XNOR2_X1 U739 ( .A(KEYINPUT21), .B(n663), .ZN(n664) );
  NAND2_X1 U740 ( .A1(n664), .A2(G2072), .ZN(G158) );
  XOR2_X1 U741 ( .A(KEYINPUT70), .B(G82), .Z(G220) );
  XNOR2_X1 U742 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U743 ( .A1(G661), .A2(G483), .ZN(n673) );
  NOR2_X1 U744 ( .A1(G220), .A2(G219), .ZN(n666) );
  XNOR2_X1 U745 ( .A(KEYINPUT22), .B(KEYINPUT85), .ZN(n665) );
  XNOR2_X1 U746 ( .A(n666), .B(n665), .ZN(n667) );
  NOR2_X1 U747 ( .A1(n667), .A2(G218), .ZN(n668) );
  NAND2_X1 U748 ( .A1(G96), .A2(n668), .ZN(n826) );
  NAND2_X1 U749 ( .A1(n826), .A2(G2106), .ZN(n672) );
  NAND2_X1 U750 ( .A1(G120), .A2(G69), .ZN(n669) );
  NOR2_X1 U751 ( .A1(G237), .A2(n669), .ZN(n670) );
  NAND2_X1 U752 ( .A1(G108), .A2(n670), .ZN(n827) );
  NAND2_X1 U753 ( .A1(n827), .A2(G567), .ZN(n671) );
  NAND2_X1 U754 ( .A1(n672), .A2(n671), .ZN(n850) );
  NOR2_X1 U755 ( .A1(n673), .A2(n850), .ZN(n674) );
  XNOR2_X1 U756 ( .A(n674), .B(KEYINPUT86), .ZN(n825) );
  NAND2_X1 U757 ( .A1(G36), .A2(n825), .ZN(G176) );
  INV_X1 U758 ( .A(G166), .ZN(G303) );
  INV_X1 U759 ( .A(G301), .ZN(G171) );
  INV_X1 U760 ( .A(KEYINPUT94), .ZN(n676) );
  NAND2_X1 U761 ( .A1(G160), .A2(G40), .ZN(n742) );
  XNOR2_X1 U762 ( .A(n676), .B(n742), .ZN(n677) );
  INV_X1 U763 ( .A(n513), .ZN(n687) );
  OR2_X1 U764 ( .A1(n687), .A2(G1961), .ZN(n679) );
  XNOR2_X1 U765 ( .A(KEYINPUT25), .B(G2078), .ZN(n951) );
  NAND2_X1 U766 ( .A1(n687), .A2(n951), .ZN(n678) );
  NAND2_X1 U767 ( .A1(n679), .A2(n678), .ZN(n713) );
  NOR2_X1 U768 ( .A1(G171), .A2(n713), .ZN(n685) );
  NAND2_X1 U769 ( .A1(G8), .A2(n513), .ZN(n778) );
  NOR2_X1 U770 ( .A1(G1966), .A2(n778), .ZN(n731) );
  NOR2_X1 U771 ( .A1(G2084), .A2(n513), .ZN(n734) );
  NOR2_X1 U772 ( .A1(n731), .A2(n734), .ZN(n680) );
  XOR2_X1 U773 ( .A(KEYINPUT97), .B(n680), .Z(n681) );
  NAND2_X1 U774 ( .A1(G8), .A2(n681), .ZN(n682) );
  XNOR2_X1 U775 ( .A(KEYINPUT30), .B(n682), .ZN(n683) );
  NOR2_X1 U776 ( .A1(n683), .A2(G168), .ZN(n684) );
  NOR2_X1 U777 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U778 ( .A(KEYINPUT31), .B(n686), .ZN(n718) );
  NAND2_X1 U779 ( .A1(n687), .A2(G2072), .ZN(n688) );
  XOR2_X1 U780 ( .A(KEYINPUT27), .B(n688), .Z(n690) );
  NAND2_X1 U781 ( .A1(G1956), .A2(n513), .ZN(n689) );
  NAND2_X1 U782 ( .A1(n690), .A2(n689), .ZN(n708) );
  NOR2_X1 U783 ( .A1(G299), .A2(n708), .ZN(n706) );
  INV_X1 U784 ( .A(G1996), .ZN(n952) );
  NOR2_X1 U785 ( .A1(n691), .A2(n952), .ZN(n693) );
  XNOR2_X1 U786 ( .A(n693), .B(n692), .ZN(n695) );
  NAND2_X1 U787 ( .A1(n722), .A2(G1341), .ZN(n694) );
  NAND2_X1 U788 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U789 ( .A(n697), .B(KEYINPUT64), .ZN(n702) );
  AND2_X1 U790 ( .A1(n702), .A2(n979), .ZN(n701) );
  OR2_X1 U791 ( .A1(G2067), .A2(n513), .ZN(n699) );
  INV_X1 U792 ( .A(G1348), .ZN(n995) );
  NAND2_X1 U793 ( .A1(n995), .A2(n513), .ZN(n698) );
  NAND2_X1 U794 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U795 ( .A1(n701), .A2(n700), .ZN(n704) );
  NOR2_X1 U796 ( .A1(n702), .A2(n979), .ZN(n703) );
  NOR2_X1 U797 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U798 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U799 ( .A(n707), .B(KEYINPUT95), .ZN(n711) );
  NAND2_X1 U800 ( .A1(G299), .A2(n708), .ZN(n709) );
  XNOR2_X1 U801 ( .A(KEYINPUT28), .B(n709), .ZN(n710) );
  NAND2_X1 U802 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U803 ( .A(n712), .B(KEYINPUT29), .ZN(n715) );
  AND2_X1 U804 ( .A1(G171), .A2(n713), .ZN(n714) );
  NOR2_X1 U805 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U806 ( .A(KEYINPUT96), .B(n716), .ZN(n717) );
  NOR2_X1 U807 ( .A1(n718), .A2(n717), .ZN(n720) );
  INV_X1 U808 ( .A(KEYINPUT98), .ZN(n719) );
  XNOR2_X1 U809 ( .A(n720), .B(n719), .ZN(n733) );
  NAND2_X1 U810 ( .A1(n733), .A2(G286), .ZN(n729) );
  INV_X1 U811 ( .A(G8), .ZN(n727) );
  NOR2_X1 U812 ( .A1(G1971), .A2(n778), .ZN(n721) );
  XNOR2_X1 U813 ( .A(KEYINPUT99), .B(n721), .ZN(n725) );
  NOR2_X1 U814 ( .A1(G2090), .A2(n513), .ZN(n723) );
  NOR2_X1 U815 ( .A1(G166), .A2(n723), .ZN(n724) );
  NAND2_X1 U816 ( .A1(n725), .A2(n724), .ZN(n726) );
  OR2_X1 U817 ( .A1(n727), .A2(n726), .ZN(n728) );
  INV_X1 U818 ( .A(n731), .ZN(n732) );
  NAND2_X1 U819 ( .A1(G8), .A2(n734), .ZN(n735) );
  NAND2_X1 U820 ( .A1(n736), .A2(n735), .ZN(n782) );
  INV_X1 U821 ( .A(n778), .ZN(n737) );
  NAND2_X1 U822 ( .A1(G1976), .A2(G288), .ZN(n971) );
  AND2_X1 U823 ( .A1(n737), .A2(n971), .ZN(n738) );
  NOR2_X1 U824 ( .A1(KEYINPUT33), .A2(n738), .ZN(n741) );
  NOR2_X1 U825 ( .A1(G1976), .A2(G288), .ZN(n770) );
  NAND2_X1 U826 ( .A1(n770), .A2(KEYINPUT33), .ZN(n739) );
  NOR2_X1 U827 ( .A1(n778), .A2(n739), .ZN(n740) );
  NOR2_X1 U828 ( .A1(n741), .A2(n740), .ZN(n766) );
  XOR2_X1 U829 ( .A(G1981), .B(G305), .Z(n987) );
  NOR2_X1 U830 ( .A1(n743), .A2(n742), .ZN(n817) );
  NAND2_X1 U831 ( .A1(G107), .A2(n876), .ZN(n750) );
  NAND2_X1 U832 ( .A1(G95), .A2(n879), .ZN(n745) );
  NAND2_X1 U833 ( .A1(G119), .A2(n875), .ZN(n744) );
  NAND2_X1 U834 ( .A1(n745), .A2(n744), .ZN(n748) );
  NAND2_X1 U835 ( .A1(G131), .A2(n880), .ZN(n746) );
  XNOR2_X1 U836 ( .A(KEYINPUT89), .B(n746), .ZN(n747) );
  NOR2_X1 U837 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U838 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U839 ( .A(n751), .B(KEYINPUT90), .ZN(n888) );
  NAND2_X1 U840 ( .A1(G1991), .A2(n888), .ZN(n762) );
  NAND2_X1 U841 ( .A1(G129), .A2(n875), .ZN(n753) );
  NAND2_X1 U842 ( .A1(G117), .A2(n876), .ZN(n752) );
  NAND2_X1 U843 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U844 ( .A(KEYINPUT91), .B(n754), .ZN(n760) );
  NAND2_X1 U845 ( .A1(G105), .A2(n879), .ZN(n755) );
  XOR2_X1 U846 ( .A(KEYINPUT38), .B(n755), .Z(n758) );
  NAND2_X1 U847 ( .A1(n880), .A2(G141), .ZN(n756) );
  XOR2_X1 U848 ( .A(KEYINPUT92), .B(n756), .Z(n757) );
  NOR2_X1 U849 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U850 ( .A1(n760), .A2(n759), .ZN(n890) );
  NAND2_X1 U851 ( .A1(G1996), .A2(n890), .ZN(n761) );
  NAND2_X1 U852 ( .A1(n762), .A2(n761), .ZN(n763) );
  XOR2_X1 U853 ( .A(KEYINPUT93), .B(n763), .Z(n933) );
  NAND2_X1 U854 ( .A1(n817), .A2(n933), .ZN(n806) );
  XNOR2_X1 U855 ( .A(G1986), .B(G290), .ZN(n985) );
  NAND2_X1 U856 ( .A1(n817), .A2(n985), .ZN(n764) );
  AND2_X1 U857 ( .A1(n806), .A2(n764), .ZN(n779) );
  AND2_X1 U858 ( .A1(n987), .A2(n779), .ZN(n765) );
  AND2_X1 U859 ( .A1(n766), .A2(n765), .ZN(n768) );
  AND2_X1 U860 ( .A1(n782), .A2(n768), .ZN(n767) );
  NAND2_X1 U861 ( .A1(n784), .A2(n767), .ZN(n775) );
  INV_X1 U862 ( .A(n768), .ZN(n773) );
  NOR2_X1 U863 ( .A1(G1971), .A2(G303), .ZN(n769) );
  NOR2_X1 U864 ( .A1(n770), .A2(n769), .ZN(n978) );
  INV_X1 U865 ( .A(KEYINPUT33), .ZN(n771) );
  AND2_X1 U866 ( .A1(n978), .A2(n771), .ZN(n772) );
  OR2_X1 U867 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U868 ( .A1(n775), .A2(n774), .ZN(n794) );
  NOR2_X1 U869 ( .A1(G1981), .A2(G305), .ZN(n776) );
  XOR2_X1 U870 ( .A(n776), .B(KEYINPUT24), .Z(n777) );
  NOR2_X1 U871 ( .A1(n778), .A2(n777), .ZN(n786) );
  OR2_X1 U872 ( .A1(n786), .A2(n778), .ZN(n780) );
  NAND2_X1 U873 ( .A1(n780), .A2(n779), .ZN(n790) );
  INV_X1 U874 ( .A(n790), .ZN(n781) );
  AND2_X1 U875 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U876 ( .A1(n784), .A2(n783), .ZN(n792) );
  NOR2_X1 U877 ( .A1(G2090), .A2(G303), .ZN(n785) );
  NAND2_X1 U878 ( .A1(G8), .A2(n785), .ZN(n788) );
  INV_X1 U879 ( .A(n786), .ZN(n787) );
  AND2_X1 U880 ( .A1(n788), .A2(n787), .ZN(n789) );
  OR2_X1 U881 ( .A1(n790), .A2(n789), .ZN(n791) );
  AND2_X1 U882 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U883 ( .A1(n794), .A2(n793), .ZN(n804) );
  NAND2_X1 U884 ( .A1(G104), .A2(n879), .ZN(n796) );
  NAND2_X1 U885 ( .A1(G140), .A2(n880), .ZN(n795) );
  NAND2_X1 U886 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U887 ( .A(KEYINPUT34), .B(n797), .ZN(n802) );
  NAND2_X1 U888 ( .A1(G128), .A2(n875), .ZN(n799) );
  NAND2_X1 U889 ( .A1(G116), .A2(n876), .ZN(n798) );
  NAND2_X1 U890 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U891 ( .A(KEYINPUT35), .B(n800), .Z(n801) );
  NOR2_X1 U892 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U893 ( .A(KEYINPUT36), .B(n803), .ZN(n859) );
  XNOR2_X1 U894 ( .A(G2067), .B(KEYINPUT37), .ZN(n815) );
  NOR2_X1 U895 ( .A1(n859), .A2(n815), .ZN(n930) );
  NAND2_X1 U896 ( .A1(n817), .A2(n930), .ZN(n813) );
  NAND2_X1 U897 ( .A1(n804), .A2(n813), .ZN(n805) );
  XNOR2_X1 U898 ( .A(n805), .B(KEYINPUT100), .ZN(n820) );
  NOR2_X1 U899 ( .A1(G1996), .A2(n890), .ZN(n938) );
  INV_X1 U900 ( .A(n806), .ZN(n809) );
  NOR2_X1 U901 ( .A1(G1991), .A2(n888), .ZN(n927) );
  NOR2_X1 U902 ( .A1(G1986), .A2(G290), .ZN(n807) );
  NOR2_X1 U903 ( .A1(n927), .A2(n807), .ZN(n808) );
  NOR2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U905 ( .A1(n938), .A2(n810), .ZN(n811) );
  XOR2_X1 U906 ( .A(n811), .B(KEYINPUT39), .Z(n812) );
  XNOR2_X1 U907 ( .A(KEYINPUT101), .B(n812), .ZN(n814) );
  NAND2_X1 U908 ( .A1(n814), .A2(n813), .ZN(n816) );
  NAND2_X1 U909 ( .A1(n859), .A2(n815), .ZN(n940) );
  NAND2_X1 U910 ( .A1(n816), .A2(n940), .ZN(n818) );
  NAND2_X1 U911 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U912 ( .A1(n820), .A2(n819), .ZN(n821) );
  XNOR2_X1 U913 ( .A(n821), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U914 ( .A1(G2106), .A2(n822), .ZN(G217) );
  AND2_X1 U915 ( .A1(G15), .A2(G2), .ZN(n823) );
  NAND2_X1 U916 ( .A1(G661), .A2(n823), .ZN(G259) );
  NAND2_X1 U917 ( .A1(G3), .A2(G1), .ZN(n824) );
  NAND2_X1 U918 ( .A1(n825), .A2(n824), .ZN(G188) );
  XOR2_X1 U919 ( .A(G69), .B(KEYINPUT102), .Z(G235) );
  INV_X1 U921 ( .A(G120), .ZN(G236) );
  INV_X1 U922 ( .A(G96), .ZN(G221) );
  NOR2_X1 U923 ( .A1(n827), .A2(n826), .ZN(G325) );
  INV_X1 U924 ( .A(G325), .ZN(G261) );
  XOR2_X1 U925 ( .A(G1976), .B(G1971), .Z(n829) );
  XNOR2_X1 U926 ( .A(G1996), .B(G1991), .ZN(n828) );
  XNOR2_X1 U927 ( .A(n829), .B(n828), .ZN(n839) );
  XOR2_X1 U928 ( .A(KEYINPUT41), .B(KEYINPUT105), .Z(n831) );
  XNOR2_X1 U929 ( .A(G1966), .B(G2474), .ZN(n830) );
  XNOR2_X1 U930 ( .A(n831), .B(n830), .ZN(n835) );
  XOR2_X1 U931 ( .A(G1981), .B(G1956), .Z(n833) );
  XNOR2_X1 U932 ( .A(G1986), .B(G1961), .ZN(n832) );
  XNOR2_X1 U933 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U934 ( .A(n835), .B(n834), .Z(n837) );
  XNOR2_X1 U935 ( .A(KEYINPUT107), .B(KEYINPUT106), .ZN(n836) );
  XNOR2_X1 U936 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U937 ( .A(n839), .B(n838), .Z(G229) );
  XOR2_X1 U938 ( .A(G2100), .B(KEYINPUT104), .Z(n841) );
  XNOR2_X1 U939 ( .A(KEYINPUT103), .B(KEYINPUT43), .ZN(n840) );
  XNOR2_X1 U940 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U941 ( .A(KEYINPUT42), .B(G2090), .Z(n843) );
  XNOR2_X1 U942 ( .A(G2067), .B(G2072), .ZN(n842) );
  XNOR2_X1 U943 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U944 ( .A(n845), .B(n844), .Z(n847) );
  XNOR2_X1 U945 ( .A(G2678), .B(G2096), .ZN(n846) );
  XNOR2_X1 U946 ( .A(n847), .B(n846), .ZN(n849) );
  XOR2_X1 U947 ( .A(G2084), .B(G2078), .Z(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(G227) );
  INV_X1 U949 ( .A(n850), .ZN(G319) );
  NAND2_X1 U950 ( .A1(n875), .A2(G124), .ZN(n851) );
  XNOR2_X1 U951 ( .A(n851), .B(KEYINPUT44), .ZN(n853) );
  NAND2_X1 U952 ( .A1(G136), .A2(n880), .ZN(n852) );
  NAND2_X1 U953 ( .A1(n853), .A2(n852), .ZN(n854) );
  XNOR2_X1 U954 ( .A(KEYINPUT108), .B(n854), .ZN(n858) );
  NAND2_X1 U955 ( .A1(G100), .A2(n879), .ZN(n856) );
  NAND2_X1 U956 ( .A1(G112), .A2(n876), .ZN(n855) );
  NAND2_X1 U957 ( .A1(n856), .A2(n855), .ZN(n857) );
  NOR2_X1 U958 ( .A1(n858), .A2(n857), .ZN(G162) );
  XNOR2_X1 U959 ( .A(n924), .B(G164), .ZN(n860) );
  XNOR2_X1 U960 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U961 ( .A(KEYINPUT46), .B(KEYINPUT112), .Z(n862) );
  XNOR2_X1 U962 ( .A(KEYINPUT113), .B(KEYINPUT48), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U964 ( .A(n864), .B(n863), .Z(n874) );
  NAND2_X1 U965 ( .A1(G103), .A2(n879), .ZN(n866) );
  NAND2_X1 U966 ( .A1(G139), .A2(n880), .ZN(n865) );
  NAND2_X1 U967 ( .A1(n866), .A2(n865), .ZN(n872) );
  NAND2_X1 U968 ( .A1(G127), .A2(n875), .ZN(n868) );
  NAND2_X1 U969 ( .A1(G115), .A2(n876), .ZN(n867) );
  NAND2_X1 U970 ( .A1(n868), .A2(n867), .ZN(n869) );
  XNOR2_X1 U971 ( .A(KEYINPUT111), .B(n869), .ZN(n870) );
  XNOR2_X1 U972 ( .A(KEYINPUT47), .B(n870), .ZN(n871) );
  NOR2_X1 U973 ( .A1(n872), .A2(n871), .ZN(n919) );
  XNOR2_X1 U974 ( .A(G162), .B(n919), .ZN(n873) );
  XNOR2_X1 U975 ( .A(n874), .B(n873), .ZN(n894) );
  NAND2_X1 U976 ( .A1(G130), .A2(n875), .ZN(n878) );
  NAND2_X1 U977 ( .A1(G118), .A2(n876), .ZN(n877) );
  NAND2_X1 U978 ( .A1(n878), .A2(n877), .ZN(n887) );
  XNOR2_X1 U979 ( .A(KEYINPUT45), .B(KEYINPUT110), .ZN(n885) );
  NAND2_X1 U980 ( .A1(n879), .A2(G106), .ZN(n883) );
  NAND2_X1 U981 ( .A1(n880), .A2(G142), .ZN(n881) );
  XOR2_X1 U982 ( .A(KEYINPUT109), .B(n881), .Z(n882) );
  NAND2_X1 U983 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U984 ( .A(n885), .B(n884), .Z(n886) );
  NOR2_X1 U985 ( .A1(n887), .A2(n886), .ZN(n892) );
  XOR2_X1 U986 ( .A(G160), .B(n888), .Z(n889) );
  XNOR2_X1 U987 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U988 ( .A(n892), .B(n891), .Z(n893) );
  XNOR2_X1 U989 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U990 ( .A1(G37), .A2(n895), .ZN(G395) );
  XNOR2_X1 U991 ( .A(n974), .B(KEYINPUT114), .ZN(n897) );
  XNOR2_X1 U992 ( .A(G171), .B(n979), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n897), .B(n896), .ZN(n900) );
  XNOR2_X1 U994 ( .A(G286), .B(n898), .ZN(n899) );
  XNOR2_X1 U995 ( .A(n900), .B(n899), .ZN(n901) );
  NOR2_X1 U996 ( .A1(G37), .A2(n901), .ZN(n902) );
  XOR2_X1 U997 ( .A(KEYINPUT115), .B(n902), .Z(G397) );
  NOR2_X1 U998 ( .A1(G229), .A2(G227), .ZN(n904) );
  XNOR2_X1 U999 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n903) );
  XNOR2_X1 U1000 ( .A(n904), .B(n903), .ZN(n915) );
  XOR2_X1 U1001 ( .A(G2451), .B(G2430), .Z(n906) );
  XNOR2_X1 U1002 ( .A(G2438), .B(G2443), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(n906), .B(n905), .ZN(n912) );
  XOR2_X1 U1004 ( .A(G2435), .B(G2454), .Z(n908) );
  XNOR2_X1 U1005 ( .A(G1348), .B(G1341), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n908), .B(n907), .ZN(n910) );
  XOR2_X1 U1007 ( .A(G2446), .B(G2427), .Z(n909) );
  XNOR2_X1 U1008 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1009 ( .A(n912), .B(n911), .Z(n913) );
  NAND2_X1 U1010 ( .A1(G14), .A2(n913), .ZN(n918) );
  NAND2_X1 U1011 ( .A1(G319), .A2(n918), .ZN(n914) );
  NOR2_X1 U1012 ( .A1(n915), .A2(n914), .ZN(n917) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n916) );
  NAND2_X1 U1014 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(G108), .ZN(G238) );
  INV_X1 U1017 ( .A(n918), .ZN(G401) );
  XOR2_X1 U1018 ( .A(G2072), .B(n919), .Z(n921) );
  XOR2_X1 U1019 ( .A(G164), .B(G2078), .Z(n920) );
  NOR2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(KEYINPUT50), .B(n922), .ZN(n923) );
  XNOR2_X1 U1022 ( .A(n923), .B(KEYINPUT120), .ZN(n936) );
  XNOR2_X1 U1023 ( .A(G160), .B(G2084), .ZN(n925) );
  NAND2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1026 ( .A(n928), .B(KEYINPUT117), .ZN(n929) );
  NOR2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1028 ( .A(KEYINPUT118), .B(n931), .Z(n932) );
  NOR2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1030 ( .A(KEYINPUT119), .B(n934), .Z(n935) );
  NAND2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n943) );
  XOR2_X1 U1032 ( .A(G2090), .B(G162), .Z(n937) );
  NOR2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1034 ( .A(KEYINPUT51), .B(n939), .Z(n941) );
  NAND2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1036 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1037 ( .A(KEYINPUT52), .B(n944), .ZN(n945) );
  XNOR2_X1 U1038 ( .A(KEYINPUT55), .B(KEYINPUT121), .ZN(n947) );
  NAND2_X1 U1039 ( .A1(n945), .A2(n947), .ZN(n946) );
  NAND2_X1 U1040 ( .A1(n946), .A2(G29), .ZN(n1025) );
  XNOR2_X1 U1041 ( .A(G29), .B(KEYINPUT123), .ZN(n968) );
  XNOR2_X1 U1042 ( .A(n947), .B(KEYINPUT122), .ZN(n966) );
  XNOR2_X1 U1043 ( .A(G2090), .B(G35), .ZN(n961) );
  XOR2_X1 U1044 ( .A(G1991), .B(G25), .Z(n948) );
  NAND2_X1 U1045 ( .A1(n948), .A2(G28), .ZN(n958) );
  XNOR2_X1 U1046 ( .A(G2067), .B(G26), .ZN(n950) );
  XNOR2_X1 U1047 ( .A(G33), .B(G2072), .ZN(n949) );
  NOR2_X1 U1048 ( .A1(n950), .A2(n949), .ZN(n956) );
  XOR2_X1 U1049 ( .A(n951), .B(G27), .Z(n954) );
  XOR2_X1 U1050 ( .A(n952), .B(G32), .Z(n953) );
  NOR2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1054 ( .A(KEYINPUT53), .B(n959), .ZN(n960) );
  NOR2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n964) );
  XOR2_X1 U1056 ( .A(G2084), .B(G34), .Z(n962) );
  XNOR2_X1 U1057 ( .A(KEYINPUT54), .B(n962), .ZN(n963) );
  NAND2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1059 ( .A(n966), .B(n965), .ZN(n967) );
  NAND2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1061 ( .A1(n969), .A2(G11), .ZN(n1023) );
  XNOR2_X1 U1062 ( .A(G16), .B(KEYINPUT56), .ZN(n993) );
  NAND2_X1 U1063 ( .A1(G1971), .A2(G303), .ZN(n970) );
  NAND2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n973) );
  XNOR2_X1 U1065 ( .A(G1961), .B(G301), .ZN(n972) );
  NOR2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n983) );
  XNOR2_X1 U1067 ( .A(n974), .B(G1341), .ZN(n976) );
  XNOR2_X1 U1068 ( .A(G299), .B(G1956), .ZN(n975) );
  NOR2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n981) );
  XNOR2_X1 U1071 ( .A(n979), .B(n995), .ZN(n980) );
  NOR2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1073 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1074 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1075 ( .A(KEYINPUT124), .B(n986), .ZN(n991) );
  XNOR2_X1 U1076 ( .A(G1966), .B(G168), .ZN(n988) );
  NAND2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1078 ( .A(KEYINPUT57), .B(n989), .ZN(n990) );
  NAND2_X1 U1079 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1080 ( .A1(n993), .A2(n992), .ZN(n1021) );
  INV_X1 U1081 ( .A(G16), .ZN(n1019) );
  XNOR2_X1 U1082 ( .A(KEYINPUT125), .B(G1966), .ZN(n994) );
  XNOR2_X1 U1083 ( .A(n994), .B(G21), .ZN(n1014) );
  XNOR2_X1 U1084 ( .A(KEYINPUT59), .B(G4), .ZN(n996) );
  XNOR2_X1 U1085 ( .A(n996), .B(n995), .ZN(n998) );
  XNOR2_X1 U1086 ( .A(G20), .B(G1956), .ZN(n997) );
  NOR2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n1002) );
  XNOR2_X1 U1088 ( .A(G1341), .B(G19), .ZN(n1000) );
  XNOR2_X1 U1089 ( .A(G1981), .B(G6), .ZN(n999) );
  NOR2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(n1003), .B(KEYINPUT60), .ZN(n1012) );
  XNOR2_X1 U1093 ( .A(G1971), .B(G22), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(G1976), .B(G23), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1096 ( .A(KEYINPUT126), .B(n1006), .Z(n1008) );
  XNOR2_X1 U1097 ( .A(G1986), .B(G24), .ZN(n1007) );
  NOR2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1099 ( .A(KEYINPUT58), .B(n1009), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(KEYINPUT127), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1016) );
  XNOR2_X1 U1103 ( .A(G5), .B(G1961), .ZN(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1105 ( .A(KEYINPUT61), .B(n1017), .ZN(n1018) );
  NAND2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1109 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1110 ( .A(KEYINPUT62), .B(n1026), .Z(G311) );
  INV_X1 U1111 ( .A(G311), .ZN(G150) );
endmodule

