

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U554 ( .A(n1009), .ZN(n753) );
  NOR2_X1 U555 ( .A1(G2105), .A2(G2104), .ZN(n520) );
  AND2_X1 U556 ( .A1(n799), .A2(n785), .ZN(n519) );
  INV_X1 U557 ( .A(n728), .ZN(n697) );
  INV_X1 U558 ( .A(KEYINPUT28), .ZN(n708) );
  INV_X1 U559 ( .A(KEYINPUT31), .ZN(n723) );
  NAND2_X1 U560 ( .A1(n726), .A2(n725), .ZN(n740) );
  NAND2_X1 U561 ( .A1(n746), .A2(n745), .ZN(n759) );
  OR2_X1 U562 ( .A1(n750), .A2(KEYINPUT33), .ZN(n756) );
  NOR2_X1 U563 ( .A1(G1384), .A2(G164), .ZN(n677) );
  NAND2_X1 U564 ( .A1(n519), .A2(n808), .ZN(n796) );
  NOR2_X1 U565 ( .A1(G651), .A2(n638), .ZN(n642) );
  XOR2_X2 U566 ( .A(KEYINPUT17), .B(n520), .Z(n886) );
  NAND2_X1 U567 ( .A1(G138), .A2(n886), .ZN(n522) );
  INV_X1 U568 ( .A(G2105), .ZN(n523) );
  AND2_X1 U569 ( .A1(n523), .A2(G2104), .ZN(n888) );
  NAND2_X1 U570 ( .A1(G102), .A2(n888), .ZN(n521) );
  NAND2_X1 U571 ( .A1(n522), .A2(n521), .ZN(n527) );
  NOR2_X1 U572 ( .A1(G2104), .A2(n523), .ZN(n881) );
  NAND2_X1 U573 ( .A1(G126), .A2(n881), .ZN(n525) );
  AND2_X1 U574 ( .A1(G2105), .A2(G2104), .ZN(n882) );
  NAND2_X1 U575 ( .A1(G114), .A2(n882), .ZN(n524) );
  NAND2_X1 U576 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X1 U577 ( .A1(n527), .A2(n526), .ZN(G164) );
  INV_X1 U578 ( .A(G651), .ZN(n531) );
  NOR2_X1 U579 ( .A1(G543), .A2(n531), .ZN(n528) );
  XOR2_X1 U580 ( .A(KEYINPUT1), .B(n528), .Z(n529) );
  XNOR2_X1 U581 ( .A(KEYINPUT66), .B(n529), .ZN(n641) );
  NAND2_X1 U582 ( .A1(n641), .A2(G64), .ZN(n530) );
  XNOR2_X1 U583 ( .A(n530), .B(KEYINPUT67), .ZN(n538) );
  NOR2_X1 U584 ( .A1(G651), .A2(G543), .ZN(n643) );
  NAND2_X1 U585 ( .A1(G90), .A2(n643), .ZN(n533) );
  XOR2_X1 U586 ( .A(KEYINPUT0), .B(G543), .Z(n638) );
  NOR2_X1 U587 ( .A1(n638), .A2(n531), .ZN(n648) );
  NAND2_X1 U588 ( .A1(G77), .A2(n648), .ZN(n532) );
  NAND2_X1 U589 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U590 ( .A(n534), .B(KEYINPUT9), .ZN(n536) );
  NAND2_X1 U591 ( .A1(G52), .A2(n642), .ZN(n535) );
  NAND2_X1 U592 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U593 ( .A1(n538), .A2(n537), .ZN(G171) );
  AND2_X1 U594 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U595 ( .A(G860), .ZN(n596) );
  NAND2_X1 U596 ( .A1(G56), .A2(n641), .ZN(n539) );
  XNOR2_X1 U597 ( .A(n539), .B(KEYINPUT14), .ZN(n541) );
  NAND2_X1 U598 ( .A1(G43), .A2(n642), .ZN(n540) );
  NAND2_X1 U599 ( .A1(n541), .A2(n540), .ZN(n548) );
  NAND2_X1 U600 ( .A1(n643), .A2(G81), .ZN(n542) );
  XNOR2_X1 U601 ( .A(n542), .B(KEYINPUT12), .ZN(n544) );
  NAND2_X1 U602 ( .A1(G68), .A2(n648), .ZN(n543) );
  NAND2_X1 U603 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U604 ( .A(KEYINPUT13), .B(n545), .ZN(n546) );
  XNOR2_X1 U605 ( .A(KEYINPUT71), .B(n546), .ZN(n547) );
  NOR2_X1 U606 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U607 ( .A(KEYINPUT72), .B(n549), .Z(n993) );
  OR2_X1 U608 ( .A1(n596), .A2(n993), .ZN(G153) );
  INV_X1 U609 ( .A(G57), .ZN(G237) );
  INV_X1 U610 ( .A(G132), .ZN(G219) );
  NAND2_X1 U611 ( .A1(G88), .A2(n643), .ZN(n551) );
  NAND2_X1 U612 ( .A1(G75), .A2(n648), .ZN(n550) );
  NAND2_X1 U613 ( .A1(n551), .A2(n550), .ZN(n555) );
  NAND2_X1 U614 ( .A1(n642), .A2(G50), .ZN(n553) );
  NAND2_X1 U615 ( .A1(G62), .A2(n641), .ZN(n552) );
  NAND2_X1 U616 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U617 ( .A1(n555), .A2(n554), .ZN(G166) );
  NAND2_X1 U618 ( .A1(n886), .A2(G137), .ZN(n556) );
  XOR2_X1 U619 ( .A(KEYINPUT65), .B(n556), .Z(n559) );
  NAND2_X1 U620 ( .A1(G101), .A2(n888), .ZN(n557) );
  XOR2_X1 U621 ( .A(KEYINPUT23), .B(n557), .Z(n558) );
  NAND2_X1 U622 ( .A1(n559), .A2(n558), .ZN(n681) );
  NAND2_X1 U623 ( .A1(G125), .A2(n881), .ZN(n561) );
  NAND2_X1 U624 ( .A1(G113), .A2(n882), .ZN(n560) );
  NAND2_X1 U625 ( .A1(n561), .A2(n560), .ZN(n678) );
  NOR2_X1 U626 ( .A1(n681), .A2(n678), .ZN(G160) );
  NAND2_X1 U627 ( .A1(n643), .A2(G89), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(KEYINPUT4), .ZN(n564) );
  NAND2_X1 U629 ( .A1(G76), .A2(n648), .ZN(n563) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(KEYINPUT5), .B(n565), .ZN(n572) );
  XNOR2_X1 U632 ( .A(KEYINPUT73), .B(KEYINPUT74), .ZN(n570) );
  NAND2_X1 U633 ( .A1(n642), .A2(G51), .ZN(n567) );
  NAND2_X1 U634 ( .A1(G63), .A2(n641), .ZN(n566) );
  NAND2_X1 U635 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n568), .B(KEYINPUT6), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(n571) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(KEYINPUT7), .B(n573), .ZN(G168) );
  XOR2_X1 U640 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U641 ( .A1(G7), .A2(G661), .ZN(n574) );
  XNOR2_X1 U642 ( .A(n574), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U643 ( .A(KEYINPUT70), .B(KEYINPUT11), .Z(n576) );
  INV_X1 U644 ( .A(G223), .ZN(n816) );
  NAND2_X1 U645 ( .A1(G567), .A2(n816), .ZN(n575) );
  XNOR2_X1 U646 ( .A(n576), .B(n575), .ZN(G234) );
  INV_X1 U647 ( .A(G171), .ZN(G301) );
  NAND2_X1 U648 ( .A1(G868), .A2(G301), .ZN(n585) );
  NAND2_X1 U649 ( .A1(G92), .A2(n643), .ZN(n578) );
  NAND2_X1 U650 ( .A1(G79), .A2(n648), .ZN(n577) );
  NAND2_X1 U651 ( .A1(n578), .A2(n577), .ZN(n582) );
  NAND2_X1 U652 ( .A1(n642), .A2(G54), .ZN(n580) );
  NAND2_X1 U653 ( .A1(G66), .A2(n641), .ZN(n579) );
  NAND2_X1 U654 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U655 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U656 ( .A(n583), .B(KEYINPUT15), .ZN(n1003) );
  INV_X1 U657 ( .A(G868), .ZN(n660) );
  NAND2_X1 U658 ( .A1(n1003), .A2(n660), .ZN(n584) );
  NAND2_X1 U659 ( .A1(n585), .A2(n584), .ZN(G284) );
  NAND2_X1 U660 ( .A1(G91), .A2(n643), .ZN(n587) );
  NAND2_X1 U661 ( .A1(G78), .A2(n648), .ZN(n586) );
  NAND2_X1 U662 ( .A1(n587), .A2(n586), .ZN(n590) );
  NAND2_X1 U663 ( .A1(n641), .A2(G65), .ZN(n588) );
  XOR2_X1 U664 ( .A(KEYINPUT68), .B(n588), .Z(n589) );
  NOR2_X1 U665 ( .A1(n590), .A2(n589), .ZN(n592) );
  NAND2_X1 U666 ( .A1(n642), .A2(G53), .ZN(n591) );
  NAND2_X1 U667 ( .A1(n592), .A2(n591), .ZN(G299) );
  NOR2_X1 U668 ( .A1(G286), .A2(n660), .ZN(n594) );
  NOR2_X1 U669 ( .A1(G868), .A2(G299), .ZN(n593) );
  NOR2_X1 U670 ( .A1(n594), .A2(n593), .ZN(n595) );
  XOR2_X1 U671 ( .A(KEYINPUT75), .B(n595), .Z(G297) );
  NAND2_X1 U672 ( .A1(n596), .A2(G559), .ZN(n597) );
  INV_X1 U673 ( .A(n1003), .ZN(n899) );
  NAND2_X1 U674 ( .A1(n597), .A2(n899), .ZN(n598) );
  XNOR2_X1 U675 ( .A(n598), .B(KEYINPUT16), .ZN(n599) );
  XNOR2_X1 U676 ( .A(KEYINPUT76), .B(n599), .ZN(G148) );
  NOR2_X1 U677 ( .A1(n993), .A2(G868), .ZN(n602) );
  NAND2_X1 U678 ( .A1(G868), .A2(n899), .ZN(n600) );
  NOR2_X1 U679 ( .A1(G559), .A2(n600), .ZN(n601) );
  NOR2_X1 U680 ( .A1(n602), .A2(n601), .ZN(G282) );
  NAND2_X1 U681 ( .A1(G123), .A2(n881), .ZN(n603) );
  XOR2_X1 U682 ( .A(KEYINPUT77), .B(n603), .Z(n604) );
  XNOR2_X1 U683 ( .A(n604), .B(KEYINPUT18), .ZN(n606) );
  NAND2_X1 U684 ( .A1(G135), .A2(n886), .ZN(n605) );
  NAND2_X1 U685 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U686 ( .A(KEYINPUT78), .B(n607), .ZN(n611) );
  NAND2_X1 U687 ( .A1(G99), .A2(n888), .ZN(n609) );
  NAND2_X1 U688 ( .A1(G111), .A2(n882), .ZN(n608) );
  NAND2_X1 U689 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U690 ( .A1(n611), .A2(n610), .ZN(n941) );
  XNOR2_X1 U691 ( .A(n941), .B(G2096), .ZN(n613) );
  INV_X1 U692 ( .A(G2100), .ZN(n612) );
  NAND2_X1 U693 ( .A1(n613), .A2(n612), .ZN(G156) );
  NAND2_X1 U694 ( .A1(G559), .A2(n899), .ZN(n614) );
  XNOR2_X1 U695 ( .A(n614), .B(n993), .ZN(n657) );
  NOR2_X1 U696 ( .A1(G860), .A2(n657), .ZN(n622) );
  NAND2_X1 U697 ( .A1(G93), .A2(n643), .ZN(n616) );
  NAND2_X1 U698 ( .A1(G80), .A2(n648), .ZN(n615) );
  NAND2_X1 U699 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U700 ( .A(KEYINPUT79), .B(n617), .ZN(n621) );
  NAND2_X1 U701 ( .A1(n641), .A2(G67), .ZN(n619) );
  NAND2_X1 U702 ( .A1(n642), .A2(G55), .ZN(n618) );
  AND2_X1 U703 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U704 ( .A1(n621), .A2(n620), .ZN(n659) );
  XOR2_X1 U705 ( .A(n622), .B(n659), .Z(G145) );
  XOR2_X1 U706 ( .A(KEYINPUT83), .B(KEYINPUT2), .Z(n624) );
  NAND2_X1 U707 ( .A1(G73), .A2(n648), .ZN(n623) );
  XNOR2_X1 U708 ( .A(n624), .B(n623), .ZN(n632) );
  NAND2_X1 U709 ( .A1(n643), .A2(G86), .ZN(n626) );
  NAND2_X1 U710 ( .A1(G61), .A2(n641), .ZN(n625) );
  NAND2_X1 U711 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U712 ( .A(KEYINPUT82), .B(n627), .ZN(n630) );
  NAND2_X1 U713 ( .A1(n642), .A2(G48), .ZN(n628) );
  XOR2_X1 U714 ( .A(KEYINPUT84), .B(n628), .Z(n629) );
  NOR2_X1 U715 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U716 ( .A1(n632), .A2(n631), .ZN(G305) );
  NAND2_X1 U717 ( .A1(G49), .A2(n642), .ZN(n634) );
  NAND2_X1 U718 ( .A1(G74), .A2(G651), .ZN(n633) );
  NAND2_X1 U719 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U720 ( .A(KEYINPUT80), .B(n635), .ZN(n636) );
  NOR2_X1 U721 ( .A1(n641), .A2(n636), .ZN(n637) );
  XOR2_X1 U722 ( .A(KEYINPUT81), .B(n637), .Z(n640) );
  NAND2_X1 U723 ( .A1(n638), .A2(G87), .ZN(n639) );
  NAND2_X1 U724 ( .A1(n640), .A2(n639), .ZN(G288) );
  AND2_X1 U725 ( .A1(G60), .A2(n641), .ZN(n647) );
  NAND2_X1 U726 ( .A1(G47), .A2(n642), .ZN(n645) );
  NAND2_X1 U727 ( .A1(G85), .A2(n643), .ZN(n644) );
  NAND2_X1 U728 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U729 ( .A1(n647), .A2(n646), .ZN(n650) );
  NAND2_X1 U730 ( .A1(n648), .A2(G72), .ZN(n649) );
  NAND2_X1 U731 ( .A1(n650), .A2(n649), .ZN(G290) );
  XNOR2_X1 U732 ( .A(G305), .B(G288), .ZN(n656) );
  INV_X1 U733 ( .A(G299), .ZN(n996) );
  XNOR2_X1 U734 ( .A(n659), .B(KEYINPUT19), .ZN(n652) );
  XNOR2_X1 U735 ( .A(G166), .B(KEYINPUT85), .ZN(n651) );
  XNOR2_X1 U736 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U737 ( .A(n996), .B(n653), .ZN(n654) );
  XNOR2_X1 U738 ( .A(n654), .B(G290), .ZN(n655) );
  XNOR2_X1 U739 ( .A(n656), .B(n655), .ZN(n902) );
  XNOR2_X1 U740 ( .A(n902), .B(n657), .ZN(n658) );
  NAND2_X1 U741 ( .A1(n658), .A2(G868), .ZN(n662) );
  NAND2_X1 U742 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U743 ( .A1(n662), .A2(n661), .ZN(G295) );
  NAND2_X1 U744 ( .A1(G2078), .A2(G2084), .ZN(n664) );
  XOR2_X1 U745 ( .A(KEYINPUT20), .B(KEYINPUT86), .Z(n663) );
  XNOR2_X1 U746 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U747 ( .A1(n665), .A2(G2090), .ZN(n666) );
  XOR2_X1 U748 ( .A(KEYINPUT21), .B(n666), .Z(n667) );
  XNOR2_X1 U749 ( .A(KEYINPUT87), .B(n667), .ZN(n668) );
  NAND2_X1 U750 ( .A1(n668), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U751 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U752 ( .A(KEYINPUT69), .B(G82), .ZN(G220) );
  NOR2_X1 U753 ( .A1(G219), .A2(G220), .ZN(n669) );
  XOR2_X1 U754 ( .A(KEYINPUT22), .B(n669), .Z(n670) );
  NOR2_X1 U755 ( .A1(G218), .A2(n670), .ZN(n671) );
  NAND2_X1 U756 ( .A1(G96), .A2(n671), .ZN(n821) );
  NAND2_X1 U757 ( .A1(n821), .A2(G2106), .ZN(n675) );
  NAND2_X1 U758 ( .A1(G69), .A2(G120), .ZN(n672) );
  NOR2_X1 U759 ( .A1(G237), .A2(n672), .ZN(n673) );
  NAND2_X1 U760 ( .A1(G108), .A2(n673), .ZN(n822) );
  NAND2_X1 U761 ( .A1(n822), .A2(G567), .ZN(n674) );
  NAND2_X1 U762 ( .A1(n675), .A2(n674), .ZN(n910) );
  NAND2_X1 U763 ( .A1(G483), .A2(G661), .ZN(n676) );
  NOR2_X1 U764 ( .A1(n910), .A2(n676), .ZN(n818) );
  NAND2_X1 U765 ( .A1(n818), .A2(G36), .ZN(G176) );
  INV_X1 U766 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U767 ( .A(n677), .B(KEYINPUT64), .ZN(n767) );
  INV_X1 U768 ( .A(n767), .ZN(n682) );
  INV_X1 U769 ( .A(G40), .ZN(n679) );
  OR2_X1 U770 ( .A1(n679), .A2(n678), .ZN(n680) );
  OR2_X1 U771 ( .A1(n681), .A2(n680), .ZN(n766) );
  OR2_X1 U772 ( .A1(n682), .A2(n766), .ZN(n728) );
  NAND2_X2 U773 ( .A1(G8), .A2(n728), .ZN(n760) );
  NOR2_X1 U774 ( .A1(G1981), .A2(G305), .ZN(n683) );
  XNOR2_X1 U775 ( .A(n683), .B(KEYINPUT24), .ZN(n684) );
  XNOR2_X1 U776 ( .A(KEYINPUT91), .B(n684), .ZN(n685) );
  NOR2_X1 U777 ( .A1(n760), .A2(n685), .ZN(n765) );
  XOR2_X1 U778 ( .A(G2078), .B(KEYINPUT25), .Z(n686) );
  XNOR2_X1 U779 ( .A(KEYINPUT93), .B(n686), .ZN(n969) );
  NAND2_X1 U780 ( .A1(n697), .A2(n969), .ZN(n687) );
  XNOR2_X1 U781 ( .A(n687), .B(KEYINPUT94), .ZN(n689) );
  XOR2_X1 U782 ( .A(G1961), .B(KEYINPUT92), .Z(n922) );
  NAND2_X1 U783 ( .A1(n922), .A2(n728), .ZN(n688) );
  NAND2_X1 U784 ( .A1(n689), .A2(n688), .ZN(n720) );
  NAND2_X1 U785 ( .A1(n720), .A2(G171), .ZN(n715) );
  XNOR2_X1 U786 ( .A(KEYINPUT29), .B(KEYINPUT95), .ZN(n713) );
  NAND2_X1 U787 ( .A1(n697), .A2(G2072), .ZN(n690) );
  XNOR2_X1 U788 ( .A(n690), .B(KEYINPUT27), .ZN(n692) );
  INV_X1 U789 ( .A(G1956), .ZN(n911) );
  NOR2_X1 U790 ( .A1(n911), .A2(n697), .ZN(n691) );
  NOR2_X1 U791 ( .A1(n692), .A2(n691), .ZN(n707) );
  NAND2_X1 U792 ( .A1(n996), .A2(n707), .ZN(n706) );
  INV_X1 U793 ( .A(G1996), .ZN(n975) );
  NOR2_X1 U794 ( .A1(n728), .A2(n975), .ZN(n693) );
  XOR2_X1 U795 ( .A(n693), .B(KEYINPUT26), .Z(n695) );
  NAND2_X1 U796 ( .A1(n728), .A2(G1341), .ZN(n694) );
  NAND2_X1 U797 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U798 ( .A1(n993), .A2(n696), .ZN(n701) );
  NAND2_X1 U799 ( .A1(G1348), .A2(n728), .ZN(n699) );
  NAND2_X1 U800 ( .A1(G2067), .A2(n697), .ZN(n698) );
  NAND2_X1 U801 ( .A1(n699), .A2(n698), .ZN(n702) );
  NOR2_X1 U802 ( .A1(n1003), .A2(n702), .ZN(n700) );
  OR2_X1 U803 ( .A1(n701), .A2(n700), .ZN(n704) );
  NAND2_X1 U804 ( .A1(n1003), .A2(n702), .ZN(n703) );
  NAND2_X1 U805 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U806 ( .A1(n706), .A2(n705), .ZN(n711) );
  NOR2_X1 U807 ( .A1(n996), .A2(n707), .ZN(n709) );
  XNOR2_X1 U808 ( .A(n709), .B(n708), .ZN(n710) );
  NAND2_X1 U809 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U810 ( .A(n713), .B(n712), .ZN(n714) );
  NAND2_X1 U811 ( .A1(n715), .A2(n714), .ZN(n726) );
  NOR2_X1 U812 ( .A1(G1966), .A2(n760), .ZN(n742) );
  NOR2_X1 U813 ( .A1(G2084), .A2(n728), .ZN(n739) );
  NOR2_X1 U814 ( .A1(n742), .A2(n739), .ZN(n716) );
  XNOR2_X1 U815 ( .A(n716), .B(KEYINPUT96), .ZN(n717) );
  NAND2_X1 U816 ( .A1(n717), .A2(G8), .ZN(n718) );
  XNOR2_X1 U817 ( .A(n718), .B(KEYINPUT30), .ZN(n719) );
  NOR2_X1 U818 ( .A1(n719), .A2(G168), .ZN(n722) );
  NOR2_X1 U819 ( .A1(G171), .A2(n720), .ZN(n721) );
  NOR2_X1 U820 ( .A1(n722), .A2(n721), .ZN(n724) );
  XNOR2_X1 U821 ( .A(n724), .B(n723), .ZN(n725) );
  NAND2_X1 U822 ( .A1(n740), .A2(G286), .ZN(n737) );
  INV_X1 U823 ( .A(G8), .ZN(n735) );
  NOR2_X1 U824 ( .A1(G1971), .A2(n760), .ZN(n727) );
  XOR2_X1 U825 ( .A(KEYINPUT97), .B(n727), .Z(n730) );
  NOR2_X1 U826 ( .A1(G2090), .A2(n728), .ZN(n729) );
  NOR2_X1 U827 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U828 ( .A(KEYINPUT98), .B(n731), .Z(n732) );
  NOR2_X1 U829 ( .A1(G166), .A2(n732), .ZN(n733) );
  XNOR2_X1 U830 ( .A(n733), .B(KEYINPUT99), .ZN(n734) );
  OR2_X1 U831 ( .A1(n735), .A2(n734), .ZN(n736) );
  AND2_X1 U832 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U833 ( .A(n738), .B(KEYINPUT32), .ZN(n746) );
  NAND2_X1 U834 ( .A1(G8), .A2(n739), .ZN(n744) );
  INV_X1 U835 ( .A(n740), .ZN(n741) );
  NOR2_X1 U836 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U837 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n751) );
  NOR2_X1 U839 ( .A1(G1971), .A2(G303), .ZN(n747) );
  NOR2_X1 U840 ( .A1(n751), .A2(n747), .ZN(n1015) );
  NAND2_X1 U841 ( .A1(n759), .A2(n1015), .ZN(n748) );
  NAND2_X1 U842 ( .A1(G1976), .A2(G288), .ZN(n994) );
  NAND2_X1 U843 ( .A1(n748), .A2(n994), .ZN(n749) );
  NOR2_X1 U844 ( .A1(n749), .A2(n760), .ZN(n750) );
  NAND2_X1 U845 ( .A1(n751), .A2(KEYINPUT33), .ZN(n752) );
  NOR2_X1 U846 ( .A1(n760), .A2(n752), .ZN(n754) );
  XOR2_X1 U847 ( .A(G1981), .B(G305), .Z(n1009) );
  NOR2_X1 U848 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U849 ( .A1(n756), .A2(n755), .ZN(n763) );
  NOR2_X1 U850 ( .A1(G2090), .A2(G303), .ZN(n757) );
  NAND2_X1 U851 ( .A1(G8), .A2(n757), .ZN(n758) );
  NAND2_X1 U852 ( .A1(n759), .A2(n758), .ZN(n761) );
  NAND2_X1 U853 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U854 ( .A1(n763), .A2(n762), .ZN(n764) );
  NOR2_X1 U855 ( .A1(n765), .A2(n764), .ZN(n797) );
  NOR2_X1 U856 ( .A1(n767), .A2(n766), .ZN(n811) );
  NAND2_X1 U857 ( .A1(G105), .A2(n888), .ZN(n768) );
  XOR2_X1 U858 ( .A(KEYINPUT89), .B(n768), .Z(n769) );
  XNOR2_X1 U859 ( .A(n769), .B(KEYINPUT38), .ZN(n771) );
  NAND2_X1 U860 ( .A1(G129), .A2(n881), .ZN(n770) );
  NAND2_X1 U861 ( .A1(n771), .A2(n770), .ZN(n775) );
  NAND2_X1 U862 ( .A1(G141), .A2(n886), .ZN(n773) );
  NAND2_X1 U863 ( .A1(G117), .A2(n882), .ZN(n772) );
  NAND2_X1 U864 ( .A1(n773), .A2(n772), .ZN(n774) );
  NOR2_X1 U865 ( .A1(n775), .A2(n774), .ZN(n776) );
  XOR2_X1 U866 ( .A(KEYINPUT90), .B(n776), .Z(n863) );
  NAND2_X1 U867 ( .A1(G1996), .A2(n863), .ZN(n784) );
  NAND2_X1 U868 ( .A1(G131), .A2(n886), .ZN(n778) );
  NAND2_X1 U869 ( .A1(G119), .A2(n881), .ZN(n777) );
  NAND2_X1 U870 ( .A1(n778), .A2(n777), .ZN(n782) );
  NAND2_X1 U871 ( .A1(G95), .A2(n888), .ZN(n780) );
  NAND2_X1 U872 ( .A1(G107), .A2(n882), .ZN(n779) );
  NAND2_X1 U873 ( .A1(n780), .A2(n779), .ZN(n781) );
  OR2_X1 U874 ( .A1(n782), .A2(n781), .ZN(n862) );
  NAND2_X1 U875 ( .A1(G1991), .A2(n862), .ZN(n783) );
  NAND2_X1 U876 ( .A1(n784), .A2(n783), .ZN(n947) );
  NAND2_X1 U877 ( .A1(n811), .A2(n947), .ZN(n799) );
  XNOR2_X1 U878 ( .A(G1986), .B(G290), .ZN(n1000) );
  NAND2_X1 U879 ( .A1(n811), .A2(n1000), .ZN(n785) );
  NAND2_X1 U880 ( .A1(G140), .A2(n886), .ZN(n787) );
  NAND2_X1 U881 ( .A1(G104), .A2(n888), .ZN(n786) );
  NAND2_X1 U882 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U883 ( .A(KEYINPUT34), .B(n788), .ZN(n793) );
  NAND2_X1 U884 ( .A1(G128), .A2(n881), .ZN(n790) );
  NAND2_X1 U885 ( .A1(G116), .A2(n882), .ZN(n789) );
  NAND2_X1 U886 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U887 ( .A(n791), .B(KEYINPUT35), .Z(n792) );
  NOR2_X1 U888 ( .A1(n793), .A2(n792), .ZN(n794) );
  XOR2_X1 U889 ( .A(KEYINPUT36), .B(n794), .Z(n795) );
  XOR2_X1 U890 ( .A(KEYINPUT88), .B(n795), .Z(n897) );
  XNOR2_X1 U891 ( .A(G2067), .B(KEYINPUT37), .ZN(n809) );
  NOR2_X1 U892 ( .A1(n897), .A2(n809), .ZN(n939) );
  NAND2_X1 U893 ( .A1(n811), .A2(n939), .ZN(n808) );
  OR2_X1 U894 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U895 ( .A(n798), .B(KEYINPUT100), .ZN(n814) );
  NOR2_X1 U896 ( .A1(G1996), .A2(n863), .ZN(n956) );
  INV_X1 U897 ( .A(n799), .ZN(n802) );
  NOR2_X1 U898 ( .A1(G1986), .A2(G290), .ZN(n800) );
  NOR2_X1 U899 ( .A1(G1991), .A2(n862), .ZN(n942) );
  NOR2_X1 U900 ( .A1(n800), .A2(n942), .ZN(n801) );
  NOR2_X1 U901 ( .A1(n802), .A2(n801), .ZN(n803) );
  XOR2_X1 U902 ( .A(KEYINPUT101), .B(n803), .Z(n804) );
  NOR2_X1 U903 ( .A1(n956), .A2(n804), .ZN(n805) );
  XOR2_X1 U904 ( .A(KEYINPUT102), .B(n805), .Z(n806) );
  XOR2_X1 U905 ( .A(KEYINPUT39), .B(n806), .Z(n807) );
  NAND2_X1 U906 ( .A1(n808), .A2(n807), .ZN(n810) );
  NAND2_X1 U907 ( .A1(n897), .A2(n809), .ZN(n938) );
  NAND2_X1 U908 ( .A1(n810), .A2(n938), .ZN(n812) );
  NAND2_X1 U909 ( .A1(n812), .A2(n811), .ZN(n813) );
  NAND2_X1 U910 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U911 ( .A(n815), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U912 ( .A1(G2106), .A2(n816), .ZN(G217) );
  AND2_X1 U913 ( .A1(G15), .A2(G2), .ZN(n817) );
  NAND2_X1 U914 ( .A1(G661), .A2(n817), .ZN(G259) );
  NAND2_X1 U915 ( .A1(G3), .A2(G1), .ZN(n819) );
  NAND2_X1 U916 ( .A1(n819), .A2(n818), .ZN(n820) );
  XOR2_X1 U917 ( .A(KEYINPUT105), .B(n820), .Z(G188) );
  INV_X1 U919 ( .A(G120), .ZN(G236) );
  INV_X1 U920 ( .A(G96), .ZN(G221) );
  INV_X1 U921 ( .A(G69), .ZN(G235) );
  NOR2_X1 U922 ( .A1(n822), .A2(n821), .ZN(G325) );
  INV_X1 U923 ( .A(G325), .ZN(G261) );
  XOR2_X1 U924 ( .A(KEYINPUT103), .B(G2451), .Z(n824) );
  XNOR2_X1 U925 ( .A(G2446), .B(G2427), .ZN(n823) );
  XNOR2_X1 U926 ( .A(n824), .B(n823), .ZN(n831) );
  XOR2_X1 U927 ( .A(G2438), .B(G2435), .Z(n826) );
  XNOR2_X1 U928 ( .A(G2443), .B(G2430), .ZN(n825) );
  XNOR2_X1 U929 ( .A(n826), .B(n825), .ZN(n827) );
  XOR2_X1 U930 ( .A(n827), .B(G2454), .Z(n829) );
  XNOR2_X1 U931 ( .A(G1341), .B(G1348), .ZN(n828) );
  XNOR2_X1 U932 ( .A(n829), .B(n828), .ZN(n830) );
  XNOR2_X1 U933 ( .A(n831), .B(n830), .ZN(n832) );
  NAND2_X1 U934 ( .A1(n832), .A2(G14), .ZN(n833) );
  XOR2_X1 U935 ( .A(KEYINPUT104), .B(n833), .Z(G401) );
  XOR2_X1 U936 ( .A(KEYINPUT109), .B(G1981), .Z(n835) );
  XNOR2_X1 U937 ( .A(G1996), .B(G1991), .ZN(n834) );
  XNOR2_X1 U938 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U939 ( .A(n836), .B(KEYINPUT41), .Z(n838) );
  XNOR2_X1 U940 ( .A(G1971), .B(G1976), .ZN(n837) );
  XNOR2_X1 U941 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U942 ( .A(G1961), .B(G1956), .Z(n840) );
  XNOR2_X1 U943 ( .A(G1986), .B(G1966), .ZN(n839) );
  XNOR2_X1 U944 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U945 ( .A(n842), .B(n841), .Z(n844) );
  XNOR2_X1 U946 ( .A(KEYINPUT108), .B(G2474), .ZN(n843) );
  XNOR2_X1 U947 ( .A(n844), .B(n843), .ZN(G229) );
  XOR2_X1 U948 ( .A(KEYINPUT43), .B(KEYINPUT107), .Z(n846) );
  XNOR2_X1 U949 ( .A(KEYINPUT42), .B(G2678), .ZN(n845) );
  XNOR2_X1 U950 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U951 ( .A(KEYINPUT106), .B(G2090), .Z(n848) );
  XNOR2_X1 U952 ( .A(G2067), .B(G2072), .ZN(n847) );
  XNOR2_X1 U953 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U954 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U955 ( .A(G2096), .B(G2100), .ZN(n851) );
  XNOR2_X1 U956 ( .A(n852), .B(n851), .ZN(n854) );
  XOR2_X1 U957 ( .A(G2078), .B(G2084), .Z(n853) );
  XNOR2_X1 U958 ( .A(n854), .B(n853), .ZN(G227) );
  NAND2_X1 U959 ( .A1(n881), .A2(G124), .ZN(n855) );
  XNOR2_X1 U960 ( .A(n855), .B(KEYINPUT44), .ZN(n857) );
  NAND2_X1 U961 ( .A1(G112), .A2(n882), .ZN(n856) );
  NAND2_X1 U962 ( .A1(n857), .A2(n856), .ZN(n861) );
  NAND2_X1 U963 ( .A1(G136), .A2(n886), .ZN(n859) );
  NAND2_X1 U964 ( .A1(G100), .A2(n888), .ZN(n858) );
  NAND2_X1 U965 ( .A1(n859), .A2(n858), .ZN(n860) );
  NOR2_X1 U966 ( .A1(n861), .A2(n860), .ZN(G162) );
  XNOR2_X1 U967 ( .A(n862), .B(G162), .ZN(n865) );
  XNOR2_X1 U968 ( .A(G160), .B(n863), .ZN(n864) );
  XNOR2_X1 U969 ( .A(n865), .B(n864), .ZN(n869) );
  XOR2_X1 U970 ( .A(KEYINPUT48), .B(KEYINPUT114), .Z(n867) );
  XNOR2_X1 U971 ( .A(G164), .B(KEYINPUT46), .ZN(n866) );
  XNOR2_X1 U972 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U973 ( .A(n869), .B(n868), .Z(n880) );
  NAND2_X1 U974 ( .A1(G127), .A2(n881), .ZN(n871) );
  NAND2_X1 U975 ( .A1(G115), .A2(n882), .ZN(n870) );
  NAND2_X1 U976 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U977 ( .A(n872), .B(KEYINPUT47), .ZN(n874) );
  NAND2_X1 U978 ( .A1(G139), .A2(n886), .ZN(n873) );
  NAND2_X1 U979 ( .A1(n874), .A2(n873), .ZN(n877) );
  NAND2_X1 U980 ( .A1(n888), .A2(G103), .ZN(n875) );
  XOR2_X1 U981 ( .A(KEYINPUT112), .B(n875), .Z(n876) );
  NOR2_X1 U982 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U983 ( .A(KEYINPUT113), .B(n878), .Z(n950) );
  XNOR2_X1 U984 ( .A(n950), .B(n941), .ZN(n879) );
  XNOR2_X1 U985 ( .A(n880), .B(n879), .ZN(n895) );
  NAND2_X1 U986 ( .A1(G130), .A2(n881), .ZN(n884) );
  NAND2_X1 U987 ( .A1(G118), .A2(n882), .ZN(n883) );
  NAND2_X1 U988 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U989 ( .A(KEYINPUT110), .B(n885), .ZN(n893) );
  NAND2_X1 U990 ( .A1(n886), .A2(G142), .ZN(n887) );
  XOR2_X1 U991 ( .A(KEYINPUT111), .B(n887), .Z(n890) );
  NAND2_X1 U992 ( .A1(n888), .A2(G106), .ZN(n889) );
  NAND2_X1 U993 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U994 ( .A(n891), .B(KEYINPUT45), .Z(n892) );
  NOR2_X1 U995 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U996 ( .A(n895), .B(n894), .Z(n896) );
  XOR2_X1 U997 ( .A(n897), .B(n896), .Z(n898) );
  NOR2_X1 U998 ( .A1(G37), .A2(n898), .ZN(G395) );
  XOR2_X1 U999 ( .A(G286), .B(G171), .Z(n901) );
  XNOR2_X1 U1000 ( .A(n993), .B(n899), .ZN(n900) );
  XNOR2_X1 U1001 ( .A(n901), .B(n900), .ZN(n903) );
  XNOR2_X1 U1002 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n904), .ZN(G397) );
  OR2_X1 U1004 ( .A1(n910), .A2(G401), .ZN(n907) );
  NOR2_X1 U1005 ( .A1(G229), .A2(G227), .ZN(n905) );
  XNOR2_X1 U1006 ( .A(KEYINPUT49), .B(n905), .ZN(n906) );
  NOR2_X1 U1007 ( .A1(n907), .A2(n906), .ZN(n909) );
  NOR2_X1 U1008 ( .A1(G395), .A2(G397), .ZN(n908) );
  NAND2_X1 U1009 ( .A1(n909), .A2(n908), .ZN(G225) );
  INV_X1 U1010 ( .A(G225), .ZN(G308) );
  INV_X1 U1011 ( .A(n910), .ZN(G319) );
  INV_X1 U1012 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1013 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n921) );
  XOR2_X1 U1014 ( .A(G1341), .B(G19), .Z(n913) );
  XNOR2_X1 U1015 ( .A(n911), .B(G20), .ZN(n912) );
  NAND2_X1 U1016 ( .A1(n913), .A2(n912), .ZN(n915) );
  XNOR2_X1 U1017 ( .A(G6), .B(G1981), .ZN(n914) );
  NOR2_X1 U1018 ( .A1(n915), .A2(n914), .ZN(n919) );
  XOR2_X1 U1019 ( .A(G4), .B(KEYINPUT125), .Z(n917) );
  XNOR2_X1 U1020 ( .A(G1348), .B(KEYINPUT59), .ZN(n916) );
  XNOR2_X1 U1021 ( .A(n917), .B(n916), .ZN(n918) );
  NAND2_X1 U1022 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1023 ( .A(n921), .B(n920), .ZN(n926) );
  XOR2_X1 U1024 ( .A(n922), .B(G5), .Z(n924) );
  XNOR2_X1 U1025 ( .A(G21), .B(G1966), .ZN(n923) );
  NOR2_X1 U1026 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n933) );
  XNOR2_X1 U1028 ( .A(G1986), .B(G24), .ZN(n928) );
  XNOR2_X1 U1029 ( .A(G1971), .B(G22), .ZN(n927) );
  NOR2_X1 U1030 ( .A1(n928), .A2(n927), .ZN(n930) );
  XOR2_X1 U1031 ( .A(G1976), .B(G23), .Z(n929) );
  NAND2_X1 U1032 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1033 ( .A(KEYINPUT58), .B(n931), .ZN(n932) );
  NOR2_X1 U1034 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1035 ( .A(KEYINPUT61), .B(n934), .Z(n935) );
  NOR2_X1 U1036 ( .A1(G16), .A2(n935), .ZN(n936) );
  XNOR2_X1 U1037 ( .A(KEYINPUT127), .B(n936), .ZN(n937) );
  NAND2_X1 U1038 ( .A1(n937), .A2(G11), .ZN(n968) );
  INV_X1 U1039 ( .A(n938), .ZN(n940) );
  NOR2_X1 U1040 ( .A1(n940), .A2(n939), .ZN(n949) );
  NOR2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n945) );
  XOR2_X1 U1042 ( .A(G160), .B(G2084), .Z(n943) );
  XNOR2_X1 U1043 ( .A(KEYINPUT115), .B(n943), .ZN(n944) );
  NAND2_X1 U1044 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1046 ( .A1(n949), .A2(n948), .ZN(n961) );
  XOR2_X1 U1047 ( .A(G2072), .B(n950), .Z(n952) );
  XOR2_X1 U1048 ( .A(G164), .B(G2078), .Z(n951) );
  NOR2_X1 U1049 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1050 ( .A(KEYINPUT50), .B(n953), .ZN(n954) );
  XNOR2_X1 U1051 ( .A(n954), .B(KEYINPUT116), .ZN(n959) );
  XOR2_X1 U1052 ( .A(G2090), .B(G162), .Z(n955) );
  NOR2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1054 ( .A(KEYINPUT51), .B(n957), .Z(n958) );
  NAND2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n960) );
  NOR2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(n962), .B(KEYINPUT52), .ZN(n964) );
  INV_X1 U1058 ( .A(KEYINPUT55), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1060 ( .A1(G29), .A2(n965), .ZN(n966) );
  XNOR2_X1 U1061 ( .A(KEYINPUT117), .B(n966), .ZN(n967) );
  NOR2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n1023) );
  XOR2_X1 U1063 ( .A(G2090), .B(G35), .Z(n985) );
  XOR2_X1 U1064 ( .A(n969), .B(G27), .Z(n974) );
  XNOR2_X1 U1065 ( .A(G2067), .B(G26), .ZN(n971) );
  XNOR2_X1 U1066 ( .A(G2072), .B(G33), .ZN(n970) );
  NOR2_X1 U1067 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1068 ( .A(KEYINPUT119), .B(n972), .ZN(n973) );
  NOR2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n981) );
  XNOR2_X1 U1070 ( .A(G32), .B(n975), .ZN(n976) );
  NAND2_X1 U1071 ( .A1(n976), .A2(G28), .ZN(n979) );
  XNOR2_X1 U1072 ( .A(G25), .B(G1991), .ZN(n977) );
  XNOR2_X1 U1073 ( .A(KEYINPUT118), .B(n977), .ZN(n978) );
  NOR2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1076 ( .A(n982), .B(KEYINPUT120), .ZN(n983) );
  XNOR2_X1 U1077 ( .A(n983), .B(KEYINPUT53), .ZN(n984) );
  NAND2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n988) );
  XNOR2_X1 U1079 ( .A(G34), .B(G2084), .ZN(n986) );
  XNOR2_X1 U1080 ( .A(KEYINPUT54), .B(n986), .ZN(n987) );
  NOR2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1082 ( .A(KEYINPUT55), .B(n989), .Z(n990) );
  NOR2_X1 U1083 ( .A1(G29), .A2(n990), .ZN(n991) );
  XOR2_X1 U1084 ( .A(KEYINPUT121), .B(n991), .Z(n1021) );
  XOR2_X1 U1085 ( .A(G16), .B(KEYINPUT56), .Z(n992) );
  XNOR2_X1 U1086 ( .A(KEYINPUT122), .B(n992), .ZN(n1019) );
  XOR2_X1 U1087 ( .A(n993), .B(G1341), .Z(n995) );
  NAND2_X1 U1088 ( .A1(n995), .A2(n994), .ZN(n1017) );
  XNOR2_X1 U1089 ( .A(G171), .B(G1961), .ZN(n1007) );
  XNOR2_X1 U1090 ( .A(G1956), .B(n996), .ZN(n997) );
  XNOR2_X1 U1091 ( .A(n997), .B(KEYINPUT124), .ZN(n1002) );
  INV_X1 U1092 ( .A(G1971), .ZN(n998) );
  NOR2_X1 U1093 ( .A1(G166), .A2(n998), .ZN(n999) );
  NOR2_X1 U1094 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1095 ( .A1(n1002), .A2(n1001), .ZN(n1005) );
  XNOR2_X1 U1096 ( .A(G1348), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1097 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1013) );
  XOR2_X1 U1099 ( .A(G1966), .B(G168), .Z(n1008) );
  XNOR2_X1 U1100 ( .A(KEYINPUT123), .B(n1008), .ZN(n1010) );
  NAND2_X1 U1101 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1102 ( .A(KEYINPUT57), .B(n1011), .Z(n1012) );
  NOR2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1024), .Z(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

