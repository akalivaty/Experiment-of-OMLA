//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 0 0 0 0 1 0 1 1 0 0 0 1 0 1 1 0 1 0 0 0 0 1 1 0 0 1 1 0 0 0 0 1 0 0 1 1 0 0 1 0 1 0 1 1 1 1 1 1 0 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n565, new_n566, new_n567, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n587, new_n588, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n625, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1206;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT66), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT67), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n465), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT70), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n470), .B1(new_n462), .B2(KEYINPUT3), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n468), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G137), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n464), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G125), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n465), .A2(G2104), .ZN(new_n477));
  OAI21_X1  g052(.A(KEYINPUT68), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n465), .A2(G2104), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n479), .A2(new_n467), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n475), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(G113), .A2(G2104), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g059(.A(G2105), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT69), .ZN(new_n486));
  AND3_X1   g061(.A1(new_n479), .A2(new_n467), .A3(new_n480), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n480), .B1(new_n479), .B2(new_n467), .ZN(new_n488));
  OAI21_X1  g063(.A(G125), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(new_n483), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n490), .A2(new_n491), .A3(G2105), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n474), .B1(new_n486), .B2(new_n492), .ZN(G160));
  OR2_X1    g068(.A1(G100), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n495));
  INV_X1    g070(.A(G124), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n471), .A2(new_n466), .A3(G2105), .A4(new_n467), .ZN(new_n497));
  INV_X1    g072(.A(G136), .ZN(new_n498));
  OAI221_X1 g073(.A(new_n495), .B1(new_n496), .B2(new_n497), .C1(new_n472), .C2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G162));
  OAI21_X1  g075(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n502), .B1(G114), .B2(new_n469), .ZN(new_n503));
  INV_X1    g078(.A(G126), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n497), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G138), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n506), .A2(G2105), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n471), .A2(new_n466), .A3(new_n507), .A4(new_n467), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT4), .ZN(new_n509));
  NOR3_X1   g084(.A1(new_n506), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n510), .B1(new_n487), .B2(new_n488), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n505), .B1(new_n509), .B2(new_n511), .ZN(G164));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n513), .B1(new_n514), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n516), .A2(KEYINPUT71), .A3(KEYINPUT5), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n514), .A2(G543), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT6), .B(G651), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n520), .A2(G88), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(G543), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G50), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT72), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT72), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n522), .A2(new_n528), .A3(new_n525), .ZN(new_n529));
  NAND2_X1  g104(.A1(G75), .A2(G543), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n518), .A2(new_n519), .ZN(new_n531));
  INV_X1    g106(.A(G62), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n527), .A2(new_n529), .B1(G651), .B2(new_n533), .ZN(G166));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT75), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n520), .A2(new_n521), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G89), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n524), .A2(G51), .ZN(new_n540));
  AND2_X1   g115(.A1(G63), .A2(G651), .ZN(new_n541));
  AOI21_X1  g116(.A(KEYINPUT73), .B1(new_n520), .B2(new_n541), .ZN(new_n542));
  AND4_X1   g117(.A1(KEYINPUT73), .A2(new_n518), .A3(new_n519), .A4(new_n541), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n540), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT74), .ZN(new_n545));
  OAI211_X1 g120(.A(new_n537), .B(new_n539), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n544), .A2(new_n545), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n546), .A2(new_n547), .ZN(G168));
  AOI22_X1  g123(.A1(new_n520), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G651), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n524), .A2(G52), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n520), .A2(new_n521), .ZN(new_n553));
  XNOR2_X1  g128(.A(KEYINPUT76), .B(G90), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n551), .A2(new_n555), .ZN(G171));
  AOI22_X1  g131(.A1(new_n520), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n557), .A2(new_n550), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n524), .A2(G43), .ZN(new_n559));
  INV_X1    g134(.A(G81), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n553), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT77), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  AND2_X1   g144(.A1(KEYINPUT78), .A2(KEYINPUT9), .ZN(new_n570));
  OR3_X1    g145(.A1(new_n523), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NOR2_X1   g146(.A1(KEYINPUT78), .A2(KEYINPUT9), .ZN(new_n572));
  OAI22_X1  g147(.A1(new_n523), .A2(new_n569), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT79), .ZN(new_n575));
  NAND2_X1  g150(.A1(G78), .A2(G543), .ZN(new_n576));
  XOR2_X1   g151(.A(new_n576), .B(KEYINPUT80), .Z(new_n577));
  INV_X1    g152(.A(G65), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n531), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G651), .ZN(new_n580));
  INV_X1    g155(.A(G91), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n581), .B2(new_n553), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n575), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G299));
  INV_X1    g159(.A(G171), .ZN(G301));
  INV_X1    g160(.A(G168), .ZN(G286));
  NAND2_X1  g161(.A1(new_n527), .A2(new_n529), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n533), .A2(G651), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(G303));
  NAND2_X1  g164(.A1(new_n538), .A2(G87), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n524), .A2(G49), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(G288));
  NAND3_X1  g168(.A1(new_n518), .A2(G61), .A3(new_n519), .ZN(new_n594));
  NAND2_X1  g169(.A1(G73), .A2(G543), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n550), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  NAND4_X1  g172(.A1(new_n518), .A2(G86), .A3(new_n519), .A4(new_n521), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n521), .A2(G48), .A3(G543), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n597), .A2(new_n601), .ZN(G305));
  AOI22_X1  g177(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n603), .A2(new_n550), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n524), .A2(G47), .ZN(new_n605));
  INV_X1    g180(.A(G85), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n553), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(G301), .A2(G868), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT81), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n538), .A2(new_n611), .A3(G92), .ZN(new_n612));
  INV_X1    g187(.A(G92), .ZN(new_n613));
  OAI21_X1  g188(.A(KEYINPUT81), .B1(new_n553), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g189(.A(KEYINPUT10), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n524), .A2(G54), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n520), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(new_n550), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n612), .A2(KEYINPUT10), .A3(new_n614), .ZN(new_n620));
  AND2_X1   g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n610), .B1(new_n621), .B2(G868), .ZN(G284));
  XNOR2_X1  g197(.A(G284), .B(KEYINPUT82), .ZN(G321));
  INV_X1    g198(.A(G868), .ZN(new_n624));
  NAND2_X1  g199(.A1(G299), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(new_n624), .B2(G168), .ZN(G297));
  OAI21_X1  g201(.A(new_n625), .B1(new_n624), .B2(G168), .ZN(G280));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n621), .B1(new_n628), .B2(G860), .ZN(G148));
  INV_X1    g204(.A(new_n562), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(new_n624), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n619), .A2(new_n620), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n632), .A2(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n631), .B1(new_n633), .B2(new_n624), .ZN(G323));
  XOR2_X1   g209(.A(KEYINPUT83), .B(KEYINPUT11), .Z(new_n635));
  XNOR2_X1  g210(.A(G323), .B(new_n635), .ZN(G282));
  NAND2_X1  g211(.A1(new_n478), .A2(new_n481), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(new_n463), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT12), .Z(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT13), .Z(new_n640));
  XOR2_X1   g215(.A(KEYINPUT84), .B(G2100), .Z(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  INV_X1    g218(.A(G123), .ZN(new_n644));
  INV_X1    g219(.A(KEYINPUT85), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(new_n469), .B2(G111), .ZN(new_n646));
  OR2_X1    g221(.A1(G99), .A2(G2105), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(G2104), .A3(new_n647), .ZN(new_n648));
  NOR3_X1   g223(.A1(new_n645), .A2(new_n469), .A3(G111), .ZN(new_n649));
  OAI22_X1  g224(.A1(new_n497), .A2(new_n644), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(new_n472), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n650), .B1(new_n651), .B2(G135), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2096), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n642), .A2(new_n643), .A3(new_n653), .ZN(G156));
  INV_X1    g229(.A(KEYINPUT14), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2427), .B(G2438), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2430), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT15), .B(G2435), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n659), .B1(new_n658), .B2(new_n657), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2451), .B(G2454), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT16), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1341), .B(G1348), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n660), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2443), .B(G2446), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  AND3_X1   g243(.A1(new_n667), .A2(G14), .A3(new_n668), .ZN(G401));
  INV_X1    g244(.A(KEYINPUT18), .ZN(new_n670));
  XOR2_X1   g245(.A(G2084), .B(G2090), .Z(new_n671));
  XNOR2_X1  g246(.A(G2067), .B(G2678), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(KEYINPUT17), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n671), .A2(new_n672), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n670), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G2100), .ZN(new_n677));
  XOR2_X1   g252(.A(G2072), .B(G2078), .Z(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(new_n673), .B2(KEYINPUT18), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(G2096), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n677), .B(new_n680), .ZN(G227));
  XNOR2_X1  g256(.A(G1971), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT86), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1956), .B(G2474), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1961), .B(G1966), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n683), .B1(new_n684), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(new_n684), .B2(new_n689), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT20), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n686), .A2(new_n688), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n694), .A2(new_n689), .A3(new_n683), .ZN(new_n695));
  OAI211_X1 g270(.A(new_n692), .B(new_n695), .C1(new_n683), .C2(new_n694), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1991), .B(G1996), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(G229));
  NOR2_X1   g277(.A1(G4), .A2(G16), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n621), .B2(G16), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT89), .B(G1348), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT24), .ZN(new_n707));
  INV_X1    g282(.A(G34), .ZN(new_n708));
  AOI21_X1  g283(.A(G29), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(new_n707), .B2(new_n708), .ZN(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(G160), .B2(new_n711), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n712), .A2(G2084), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n711), .A2(G27), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G164), .B2(new_n711), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT95), .Z(new_n716));
  OR2_X1    g291(.A1(new_n716), .A2(G2078), .ZN(new_n717));
  INV_X1    g292(.A(G16), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G20), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT97), .Z(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT23), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G299), .B2(G16), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G1956), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n706), .A2(new_n713), .A3(new_n717), .A4(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n718), .A2(G21), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G168), .B2(new_n718), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G1966), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT93), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n711), .A2(G35), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G162), .B2(new_n711), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT29), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n731), .A2(G2090), .ZN(new_n732));
  INV_X1    g307(.A(new_n726), .ZN(new_n733));
  INV_X1    g308(.A(G1966), .ZN(new_n734));
  AOI22_X1  g309(.A1(KEYINPUT96), .A2(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n728), .B(new_n735), .C1(KEYINPUT96), .C2(new_n732), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n651), .A2(G141), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT92), .ZN(new_n738));
  INV_X1    g313(.A(new_n497), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G129), .ZN(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT26), .Z(new_n742));
  NAND2_X1  g317(.A1(new_n463), .A2(G105), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n738), .A2(new_n740), .A3(new_n742), .A4(new_n743), .ZN(new_n744));
  MUX2_X1   g319(.A(G32), .B(new_n744), .S(G29), .Z(new_n745));
  XOR2_X1   g320(.A(KEYINPUT27), .B(G1996), .Z(new_n746));
  XOR2_X1   g321(.A(new_n745), .B(new_n746), .Z(new_n747));
  NOR2_X1   g322(.A1(G29), .A2(G33), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT25), .Z(new_n750));
  INV_X1    g325(.A(G139), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n750), .B1(new_n472), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n637), .A2(G127), .ZN(new_n753));
  INV_X1    g328(.A(G115), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n753), .B1(new_n754), .B2(new_n462), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n752), .B1(new_n755), .B2(G2105), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n748), .B1(new_n756), .B2(G29), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n757), .A2(G2072), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n759), .A2(KEYINPUT91), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n711), .A2(G26), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT28), .ZN(new_n762));
  INV_X1    g337(.A(G128), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n469), .A2(G116), .ZN(new_n764));
  OAI21_X1  g339(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n765));
  OAI22_X1  g340(.A1(new_n497), .A2(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n651), .B2(G140), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n762), .B1(new_n767), .B2(new_n711), .ZN(new_n768));
  INV_X1    g343(.A(G2067), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n759), .A2(KEYINPUT91), .ZN(new_n771));
  AND3_X1   g346(.A1(new_n760), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(G171), .A2(G16), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G5), .B2(G16), .ZN(new_n774));
  INV_X1    g349(.A(G1961), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n774), .A2(new_n775), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n757), .A2(G2072), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n652), .A2(G29), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT30), .B(G28), .ZN(new_n780));
  OR2_X1    g355(.A1(KEYINPUT31), .A2(G11), .ZN(new_n781));
  NAND2_X1  g356(.A1(KEYINPUT31), .A2(G11), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n780), .A2(new_n711), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(KEYINPUT94), .B1(new_n779), .B2(new_n783), .ZN(new_n784));
  NOR4_X1   g359(.A1(new_n776), .A2(new_n777), .A3(new_n778), .A4(new_n784), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n747), .A2(new_n772), .A3(new_n785), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n716), .A2(G2078), .B1(G2084), .B2(new_n712), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n731), .A2(G2090), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n718), .A2(G19), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n562), .B2(new_n718), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT90), .B(G1341), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n779), .A2(KEYINPUT94), .A3(new_n783), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n787), .A2(new_n788), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  NOR4_X1   g369(.A1(new_n724), .A2(new_n736), .A3(new_n786), .A4(new_n794), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT98), .Z(new_n796));
  NAND2_X1  g371(.A1(new_n718), .A2(G24), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n608), .B2(new_n718), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(G1986), .Z(new_n799));
  NAND2_X1  g374(.A1(new_n711), .A2(G25), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT87), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n651), .A2(G131), .ZN(new_n802));
  INV_X1    g377(.A(G119), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n469), .A2(G107), .ZN(new_n804));
  OAI21_X1  g379(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n805));
  OAI22_X1  g380(.A1(new_n497), .A2(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n802), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n801), .B1(new_n807), .B2(new_n711), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT35), .B(G1991), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n808), .B(new_n809), .Z(new_n810));
  NAND2_X1  g385(.A1(G166), .A2(G16), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G16), .B2(G22), .ZN(new_n812));
  INV_X1    g387(.A(G1971), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n812), .A2(new_n813), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n718), .A2(G23), .ZN(new_n816));
  INV_X1    g391(.A(G288), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(new_n718), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT33), .B(G1976), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT88), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n818), .B(new_n820), .ZN(new_n821));
  MUX2_X1   g396(.A(G6), .B(G305), .S(G16), .Z(new_n822));
  XOR2_X1   g397(.A(KEYINPUT32), .B(G1981), .Z(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n814), .A2(new_n815), .A3(new_n821), .A4(new_n824), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n799), .B(new_n810), .C1(new_n825), .C2(KEYINPUT34), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(KEYINPUT34), .B2(new_n825), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT36), .Z(new_n828));
  NAND2_X1  g403(.A1(new_n796), .A2(new_n828), .ZN(G150));
  INV_X1    g404(.A(G150), .ZN(G311));
  NAND2_X1  g405(.A1(G80), .A2(G543), .ZN(new_n831));
  INV_X1    g406(.A(G67), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n831), .B1(new_n531), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(G651), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n834), .A2(KEYINPUT99), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(KEYINPUT99), .ZN(new_n836));
  AOI22_X1  g411(.A1(new_n538), .A2(G93), .B1(G55), .B2(new_n524), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(KEYINPUT100), .B2(new_n562), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(KEYINPUT100), .B2(new_n562), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT100), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n838), .A2(new_n630), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT38), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n621), .A2(G559), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT39), .ZN(new_n847));
  AOI21_X1  g422(.A(G860), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n847), .B2(new_n846), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n838), .A2(G860), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT102), .ZN(new_n851));
  XNOR2_X1  g426(.A(KEYINPUT101), .B(KEYINPUT37), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n849), .A2(new_n853), .ZN(G145));
  INV_X1    g429(.A(KEYINPUT103), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n756), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n744), .B(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n739), .A2(G130), .ZN(new_n858));
  INV_X1    g433(.A(G142), .ZN(new_n859));
  NOR3_X1   g434(.A1(new_n469), .A2(KEYINPUT104), .A3(G118), .ZN(new_n860));
  OAI21_X1  g435(.A(KEYINPUT104), .B1(new_n469), .B2(G118), .ZN(new_n861));
  OR2_X1    g436(.A1(G106), .A2(G2105), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n861), .A2(G2104), .A3(new_n862), .ZN(new_n863));
  OAI221_X1 g438(.A(new_n858), .B1(new_n472), .B2(new_n859), .C1(new_n860), .C2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n639), .B(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n857), .B(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n767), .B(G164), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n807), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n866), .B(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n652), .B(new_n499), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(G160), .ZN(new_n871));
  AOI21_X1  g446(.A(G37), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n872), .B1(new_n871), .B2(new_n869), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g449(.A(G166), .B(G290), .ZN(new_n875));
  XOR2_X1   g450(.A(G288), .B(G305), .Z(new_n876));
  XNOR2_X1  g451(.A(new_n875), .B(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT107), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n877), .B1(new_n878), .B2(KEYINPUT42), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT108), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT105), .ZN(new_n882));
  NAND2_X1  g457(.A1(G299), .A2(new_n632), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(G299), .A2(new_n632), .ZN(new_n885));
  OAI21_X1  g460(.A(KEYINPUT41), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n621), .A2(new_n583), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT41), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n887), .A2(new_n888), .A3(new_n883), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n882), .B1(new_n886), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n887), .A2(new_n883), .ZN(new_n891));
  AOI21_X1  g466(.A(KEYINPUT105), .B1(new_n891), .B2(KEYINPUT41), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n633), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n843), .B(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n891), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT106), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  NOR3_X1   g475(.A1(new_n893), .A2(KEYINPUT106), .A3(new_n895), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n881), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OR3_X1    g477(.A1(new_n893), .A2(KEYINPUT106), .A3(new_n895), .ZN(new_n903));
  OAI211_X1 g478(.A(new_n903), .B(new_n880), .C1(new_n896), .C2(new_n899), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n878), .A2(KEYINPUT42), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n902), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n905), .B1(new_n902), .B2(new_n904), .ZN(new_n907));
  OAI21_X1  g482(.A(G868), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n838), .A2(new_n624), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(G295));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n909), .ZN(G331));
  XNOR2_X1  g486(.A(G168), .B(G171), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n843), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(G168), .B(G301), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n914), .A2(new_n842), .A3(new_n840), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(new_n890), .B2(new_n892), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n913), .A2(new_n915), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(new_n897), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n917), .A2(new_n877), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT109), .ZN(new_n921));
  AOI21_X1  g496(.A(G37), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n917), .A2(new_n919), .ZN(new_n923));
  INV_X1    g498(.A(new_n877), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n917), .A2(new_n919), .A3(KEYINPUT109), .A4(new_n877), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n922), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n918), .B1(new_n886), .B2(new_n889), .ZN(new_n930));
  INV_X1    g505(.A(new_n919), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n924), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AND4_X1   g507(.A1(KEYINPUT43), .A2(new_n922), .A3(new_n926), .A4(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT44), .B1(new_n929), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n927), .A2(KEYINPUT43), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n922), .A2(new_n928), .A3(new_n926), .A4(new_n932), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n934), .A2(new_n939), .ZN(G397));
  INV_X1    g515(.A(KEYINPUT127), .ZN(new_n941));
  INV_X1    g516(.A(new_n474), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n491), .B1(new_n490), .B2(G2105), .ZN(new_n943));
  AOI211_X1 g518(.A(KEYINPUT69), .B(new_n469), .C1(new_n489), .C2(new_n483), .ZN(new_n944));
  OAI211_X1 g519(.A(G40), .B(new_n942), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT45), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n946), .B1(G164), .B2(G1384), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n744), .B(G1996), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n767), .B(new_n769), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n807), .B(new_n809), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n608), .B(G1986), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n949), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(G8), .ZN(new_n958));
  INV_X1    g533(.A(G1384), .ZN(new_n959));
  AOI22_X1  g534(.A1(new_n637), .A2(new_n510), .B1(KEYINPUT4), .B2(new_n508), .ZN(new_n960));
  OAI211_X1 g535(.A(KEYINPUT45), .B(new_n959), .C1(new_n960), .C2(new_n505), .ZN(new_n961));
  NAND4_X1  g536(.A1(G160), .A2(G40), .A3(new_n947), .A4(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n813), .ZN(new_n963));
  INV_X1    g538(.A(G40), .ZN(new_n964));
  AOI211_X1 g539(.A(new_n964), .B(new_n474), .C1(new_n486), .C2(new_n492), .ZN(new_n965));
  INV_X1    g540(.A(G2090), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT110), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n967), .B1(G164), .B2(G1384), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT50), .ZN(new_n969));
  OAI211_X1 g544(.A(KEYINPUT110), .B(new_n959), .C1(new_n960), .C2(new_n505), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n965), .A2(new_n966), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n958), .B1(new_n963), .B2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT55), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n976), .B1(G166), .B2(new_n958), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n974), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT111), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n974), .A2(new_n981), .A3(new_n978), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n590), .A2(G1976), .A3(new_n591), .A4(new_n592), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n968), .A2(new_n970), .ZN(new_n985));
  OAI211_X1 g560(.A(G8), .B(new_n984), .C1(new_n945), .C2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT52), .ZN(new_n987));
  INV_X1    g562(.A(G1981), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n597), .A2(new_n601), .A3(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(G1981), .B1(new_n596), .B2(new_n600), .ZN(new_n990));
  AND3_X1   g565(.A1(new_n989), .A2(KEYINPUT49), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT49), .B1(new_n989), .B2(new_n990), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND4_X1  g568(.A1(G160), .A2(G40), .A3(new_n968), .A4(new_n970), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n993), .A2(new_n994), .A3(G8), .ZN(new_n995));
  INV_X1    g570(.A(G1976), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT52), .B1(G288), .B2(new_n996), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n994), .A2(G8), .A3(new_n984), .A4(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n987), .A2(new_n995), .A3(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n983), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n945), .A2(new_n985), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n995), .A2(new_n996), .A3(new_n817), .ZN(new_n1002));
  AOI211_X1 g577(.A(new_n958), .B(new_n1001), .C1(new_n1002), .C2(new_n989), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1004));
  AND3_X1   g579(.A1(new_n987), .A2(new_n995), .A3(new_n998), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n963), .A2(new_n973), .ZN(new_n1006));
  AND4_X1   g581(.A1(new_n981), .A2(new_n1006), .A3(new_n978), .A4(G8), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n981), .B1(new_n974), .B2(new_n978), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1005), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n970), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n511), .A2(new_n509), .ZN(new_n1011));
  INV_X1    g586(.A(new_n505), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT110), .B1(new_n1013), .B2(new_n959), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT50), .B1(new_n1010), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1015), .A2(KEYINPUT112), .A3(new_n965), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT112), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n969), .B1(new_n968), .B2(new_n970), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1017), .B1(new_n1018), .B2(new_n945), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1013), .A2(new_n969), .A3(new_n959), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1016), .A2(new_n1019), .A3(new_n966), .A4(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n963), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n978), .B1(new_n1022), .B2(G8), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1009), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n961), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n945), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n985), .A2(new_n946), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT113), .B1(new_n1028), .B2(new_n734), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n486), .A2(new_n492), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1030), .A2(G40), .A3(new_n942), .A4(new_n961), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT45), .B1(new_n968), .B2(new_n970), .ZN(new_n1032));
  OAI211_X1 g607(.A(KEYINPUT113), .B(new_n734), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G2084), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n965), .A2(new_n1034), .A3(new_n971), .A4(new_n972), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  OAI211_X1 g611(.A(G8), .B(G168), .C1(new_n1029), .C2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT114), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n734), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1042), .A2(new_n1035), .A3(new_n1033), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1043), .A2(KEYINPUT114), .A3(G8), .A4(G168), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1039), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT63), .B1(new_n1024), .B2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1005), .B(KEYINPUT115), .C1(new_n978), .C2(new_n974), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT115), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n978), .B1(new_n1006), .B2(G8), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1048), .B1(new_n1049), .B2(new_n999), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1047), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT63), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(new_n980), .B2(new_n982), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1045), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1004), .B1(new_n1046), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(G8), .B1(new_n1029), .B2(new_n1036), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n1057));
  OAI21_X1  g632(.A(KEYINPUT119), .B1(G168), .B2(new_n958), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT119), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1059), .B(G8), .C1(new_n546), .C2(new_n547), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1056), .A2(new_n1057), .A3(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1061), .B1(new_n1029), .B2(new_n1036), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT51), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1061), .B1(new_n1043), .B2(G8), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1063), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT62), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1056), .A2(new_n1062), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1057), .B1(new_n1043), .B2(new_n1061), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1072), .A2(KEYINPUT62), .A3(new_n1063), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1074), .B1(new_n962), .B2(G2078), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1030), .A2(new_n972), .A3(G40), .A4(new_n942), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1076), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n965), .A2(KEYINPUT117), .A3(new_n971), .A4(new_n972), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1079), .A2(new_n775), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT120), .ZN(new_n1082));
  INV_X1    g657(.A(G2078), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1026), .A2(new_n1027), .A3(new_n1082), .A4(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT53), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1082), .B1(new_n1086), .B2(new_n1083), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1075), .B(new_n1081), .C1(new_n1085), .C2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(G171), .ZN(new_n1089));
  NOR3_X1   g664(.A1(new_n1009), .A2(new_n1089), .A3(new_n1023), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1069), .A2(new_n1073), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1055), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n582), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT57), .B1(new_n571), .B2(new_n573), .ZN(new_n1095));
  AOI22_X1  g670(.A1(G299), .A2(KEYINPUT57), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT45), .B1(new_n1013), .B2(new_n959), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n945), .A2(new_n1097), .A3(new_n1025), .ZN(new_n1098));
  XNOR2_X1  g673(.A(KEYINPUT56), .B(G2072), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1096), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1016), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT116), .ZN(new_n1103));
  INV_X1    g678(.A(G1956), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1102), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1103), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1101), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT116), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1102), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1096), .B1(new_n1111), .B2(new_n1100), .ZN(new_n1112));
  INV_X1    g687(.A(G1348), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1079), .A2(new_n1113), .A3(new_n1080), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1001), .A2(new_n769), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n621), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1107), .B1(new_n1112), .B2(new_n1118), .ZN(new_n1119));
  OR2_X1    g694(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n1120));
  NAND2_X1  g695(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n1121));
  INV_X1    g696(.A(G1996), .ZN(new_n1122));
  XOR2_X1   g697(.A(KEYINPUT58), .B(G1341), .Z(new_n1123));
  AOI22_X1  g698(.A1(new_n1098), .A2(new_n1122), .B1(new_n994), .B2(new_n1123), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1120), .B(new_n1121), .C1(new_n1124), .C2(new_n630), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n632), .A2(KEYINPUT60), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1114), .A2(new_n1115), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1123), .ZN(new_n1128));
  OAI22_X1  g703(.A1(new_n1001), .A2(new_n1128), .B1(new_n962), .B2(G1996), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1129), .A2(KEYINPUT118), .A3(KEYINPUT59), .A4(new_n562), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1125), .A2(new_n1127), .A3(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1114), .A2(new_n632), .A3(new_n1115), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1117), .A2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1131), .B1(new_n1133), .B2(KEYINPUT60), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1107), .A2(KEYINPUT61), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1134), .B1(new_n1112), .B2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1100), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1096), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(KEYINPUT61), .B1(new_n1139), .B2(new_n1107), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1119), .B1(new_n1136), .B2(new_n1140), .ZN(new_n1141));
  OR2_X1    g716(.A1(new_n1088), .A2(G171), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(KEYINPUT54), .ZN(new_n1143));
  XNOR2_X1  g718(.A(KEYINPUT121), .B(G2078), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n942), .A2(KEYINPUT53), .A3(G40), .A4(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1145), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1146), .A2(new_n485), .A3(new_n947), .A4(new_n961), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1081), .A2(new_n1075), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT123), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1081), .A2(KEYINPUT123), .A3(new_n1075), .A4(new_n1147), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1150), .A2(G171), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(KEYINPUT124), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT124), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1150), .A2(new_n1154), .A3(G171), .A4(new_n1151), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1143), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n999), .B1(new_n980), .B2(new_n982), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1022), .A2(G8), .ZN(new_n1159));
  INV_X1    g734(.A(new_n978), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1072), .A2(new_n1158), .A3(new_n1161), .A4(new_n1063), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1081), .A2(G301), .A3(new_n1075), .A4(new_n1147), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1164), .B1(G171), .B2(new_n1088), .ZN(new_n1165));
  OAI21_X1  g740(.A(KEYINPUT122), .B1(new_n1165), .B2(KEYINPUT54), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1089), .A2(new_n1163), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT122), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT54), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1162), .B1(new_n1166), .B2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1141), .A2(new_n1157), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n957), .B1(new_n1093), .B2(new_n1172), .ZN(new_n1173));
  OR3_X1    g748(.A1(new_n949), .A2(G1986), .A3(G290), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT48), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  OR2_X1    g751(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1177));
  OAI211_X1 g752(.A(new_n1176), .B(new_n1177), .C1(new_n955), .C2(new_n949), .ZN(new_n1178));
  NOR3_X1   g753(.A1(new_n802), .A2(new_n809), .A3(new_n806), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1179), .B1(new_n952), .B2(new_n949), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n767), .A2(new_n769), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1180), .A2(KEYINPUT125), .A3(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(new_n948), .ZN(new_n1183));
  AOI21_X1  g758(.A(KEYINPUT125), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1178), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n948), .A2(new_n1122), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1186), .B(KEYINPUT46), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n948), .B1(new_n744), .B2(new_n951), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  XNOR2_X1  g764(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1189), .B(new_n1190), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n1185), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(new_n1192), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n941), .B1(new_n1173), .B2(new_n1193), .ZN(new_n1194));
  OAI211_X1 g769(.A(new_n1091), .B(new_n1004), .C1(new_n1046), .C2(new_n1054), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n983), .A2(new_n1161), .A3(new_n1005), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1196), .A2(new_n1067), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1168), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1198));
  AOI211_X1 g773(.A(KEYINPUT122), .B(KEYINPUT54), .C1(new_n1089), .C2(new_n1163), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1197), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NOR2_X1   g775(.A1(new_n1200), .A2(new_n1156), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1195), .B1(new_n1141), .B2(new_n1201), .ZN(new_n1202));
  OAI211_X1 g777(.A(KEYINPUT127), .B(new_n1192), .C1(new_n1202), .C2(new_n957), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1194), .A2(new_n1203), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g779(.A1(G229), .A2(new_n460), .A3(G401), .A4(G227), .ZN(new_n1206));
  NAND3_X1  g780(.A1(new_n937), .A2(new_n873), .A3(new_n1206), .ZN(G225));
  INV_X1    g781(.A(G225), .ZN(G308));
endmodule


