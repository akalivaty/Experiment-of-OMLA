//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 1 1 1 1 1 1 1 1 1 1 0 0 1 1 0 0 0 1 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1 0 0 1 1 1 0 1 0 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1259, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT64), .Z(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(KEYINPUT65), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n216));
  NAND3_X1  g0016(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n213), .A2(KEYINPUT65), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n207), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  OR2_X1    g0019(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(new_n201), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n223), .A2(G50), .A3(new_n224), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n210), .A2(new_n220), .A3(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n219), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XOR2_X1   g0036(.A(G107), .B(G116), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  OR2_X1    g0042(.A1(KEYINPUT3), .A2(G33), .ZN(new_n243));
  NAND2_X1  g0043(.A1(KEYINPUT3), .A2(G33), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(G1698), .ZN(new_n246));
  NAND3_X1  g0046(.A1(new_n245), .A2(G222), .A3(new_n246), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n245), .A2(G223), .A3(G1698), .ZN(new_n248));
  INV_X1    g0048(.A(G77), .ZN(new_n249));
  OAI211_X1 g0049(.A(new_n247), .B(new_n248), .C1(new_n249), .C2(new_n245), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G1), .A3(G13), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G274), .ZN(new_n255));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n256), .B1(G41), .B2(G45), .ZN(new_n257));
  NOR3_X1   g0057(.A1(new_n253), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT66), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G41), .A2(G45), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n259), .B1(new_n260), .B2(G1), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n256), .B(KEYINPUT66), .C1(G41), .C2(G45), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n261), .A2(new_n252), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n258), .B1(new_n264), .B2(G226), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n254), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G179), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(new_n221), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G58), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT8), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT8), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G58), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n222), .A2(G33), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G20), .A2(G33), .ZN(new_n279));
  AOI22_X1  g0079(.A1(new_n276), .A2(new_n278), .B1(G150), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n203), .A2(G20), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n271), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(KEYINPUT67), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(KEYINPUT67), .ZN(new_n285));
  INV_X1    g0085(.A(G13), .ZN(new_n286));
  NOR3_X1   g0086(.A1(new_n286), .A2(new_n222), .A3(G1), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(new_n270), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n202), .B1(new_n256), .B2(G20), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n288), .A2(new_n289), .B1(new_n202), .B2(new_n287), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n284), .A2(new_n285), .A3(new_n290), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n268), .B(new_n291), .C1(G169), .C2(new_n266), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n286), .A2(G1), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G20), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT68), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT68), .ZN(new_n296));
  AND4_X1   g0096(.A1(new_n296), .A2(new_n256), .A3(G13), .A4(G20), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n270), .B1(new_n295), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n256), .A2(G20), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n299), .A2(G77), .A3(new_n300), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n273), .A2(new_n275), .ZN(new_n302));
  INV_X1    g0102(.A(new_n279), .ZN(new_n303));
  OAI22_X1  g0103(.A1(new_n302), .A2(new_n303), .B1(new_n222), .B2(new_n249), .ZN(new_n304));
  XNOR2_X1  g0104(.A(KEYINPUT15), .B(G87), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n305), .A2(new_n277), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n270), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n296), .B1(new_n293), .B2(G20), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n308), .A2(new_n297), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n249), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n301), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n245), .A2(G232), .A3(new_n246), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n245), .A2(G238), .A3(G1698), .ZN(new_n313));
  INV_X1    g0113(.A(G107), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n312), .B(new_n313), .C1(new_n314), .C2(new_n245), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n253), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n258), .B1(new_n264), .B2(G244), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n311), .B1(new_n319), .B2(G190), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(G200), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n307), .A2(new_n310), .ZN(new_n322));
  INV_X1    g0122(.A(G169), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n301), .A2(new_n322), .B1(new_n318), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n319), .A2(new_n267), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n320), .A2(new_n321), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n285), .A2(new_n290), .ZN(new_n327));
  OAI21_X1  g0127(.A(KEYINPUT9), .B1(new_n327), .B2(new_n283), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT9), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n284), .A2(new_n329), .A3(new_n285), .A4(new_n290), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT10), .ZN(new_n332));
  INV_X1    g0132(.A(G200), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n333), .B1(new_n254), .B2(new_n265), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n334), .B1(G190), .B2(new_n266), .ZN(new_n335));
  AND3_X1   g0135(.A1(new_n331), .A2(new_n332), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n332), .B1(new_n331), .B2(new_n335), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n292), .B(new_n326), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  AND2_X1   g0138(.A1(G1), .A2(G13), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n257), .A2(new_n259), .B1(new_n339), .B2(new_n251), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n340), .A2(G232), .A3(new_n262), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n255), .B1(new_n339), .B2(new_n251), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n342), .B(new_n256), .C1(G41), .C2(G45), .ZN(new_n343));
  MUX2_X1   g0143(.A(G223), .B(G226), .S(G1698), .Z(new_n344));
  AOI22_X1  g0144(.A1(new_n344), .A2(new_n245), .B1(G33), .B2(G87), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n341), .B(new_n343), .C1(new_n345), .C2(new_n252), .ZN(new_n346));
  INV_X1    g0146(.A(G190), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n348), .B1(G200), .B2(new_n346), .ZN(new_n349));
  INV_X1    g0149(.A(G68), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n272), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(G20), .B1(new_n351), .B2(new_n201), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n279), .A2(G159), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  AND2_X1   g0155(.A1(KEYINPUT3), .A2(G33), .ZN(new_n356));
  NOR2_X1   g0156(.A1(KEYINPUT3), .A2(G33), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(KEYINPUT7), .B1(new_n358), .B2(new_n222), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT7), .ZN(new_n360));
  NOR4_X1   g0160(.A1(new_n356), .A2(new_n357), .A3(new_n360), .A4(G20), .ZN(new_n361));
  NOR3_X1   g0161(.A1(new_n359), .A2(new_n361), .A3(KEYINPUT72), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n360), .B1(new_n245), .B2(G20), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT72), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n364), .A2(KEYINPUT7), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(G68), .B1(new_n363), .B2(new_n366), .ZN(new_n367));
  OAI211_X1 g0167(.A(KEYINPUT16), .B(new_n355), .C1(new_n362), .C2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT16), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n358), .A2(KEYINPUT7), .A3(new_n222), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n350), .B1(new_n363), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n369), .B1(new_n371), .B2(new_n354), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n368), .A2(new_n270), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n271), .A2(new_n294), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n276), .A2(new_n300), .ZN(new_n375));
  OAI22_X1  g0175(.A1(new_n374), .A2(new_n375), .B1(new_n294), .B2(new_n276), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n349), .A2(new_n373), .A3(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT17), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n350), .B1(new_n359), .B2(new_n365), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n363), .A2(new_n364), .A3(new_n370), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n354), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n271), .B1(new_n383), .B2(KEYINPUT16), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n376), .B1(new_n384), .B2(new_n372), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n346), .A2(G169), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(new_n267), .B2(new_n346), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(KEYINPUT18), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n373), .A2(new_n377), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT18), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(new_n391), .A3(new_n387), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n385), .A2(KEYINPUT17), .A3(new_n349), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n380), .A2(new_n389), .A3(new_n392), .A4(new_n393), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n338), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT12), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n396), .B1(new_n309), .B2(new_n350), .ZN(new_n397));
  XNOR2_X1  g0197(.A(new_n397), .B(KEYINPUT71), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n293), .A2(new_n396), .A3(G20), .A4(new_n350), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n303), .A2(new_n202), .ZN(new_n401));
  OAI22_X1  g0201(.A1(new_n277), .A2(new_n249), .B1(new_n222), .B2(G68), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n270), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  XNOR2_X1  g0203(.A(new_n403), .B(KEYINPUT11), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n299), .A2(G68), .A3(new_n300), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n400), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  OR2_X1    g0206(.A1(new_n246), .A2(G232), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n245), .B(new_n407), .C1(G226), .C2(G1698), .ZN(new_n408));
  INV_X1    g0208(.A(G33), .ZN(new_n409));
  INV_X1    g0209(.A(G97), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n252), .B1(new_n408), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT70), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT69), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n261), .A2(new_n416), .A3(new_n252), .A4(new_n262), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(G238), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n416), .B1(new_n340), .B2(new_n262), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n415), .B(new_n343), .C1(new_n418), .C2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n263), .A2(KEYINPUT69), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n422), .A2(G238), .A3(new_n417), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n415), .B1(new_n423), .B2(new_n343), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n414), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT13), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n343), .B1(new_n418), .B2(new_n419), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT70), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n420), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT13), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n429), .A2(new_n430), .A3(new_n414), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n426), .A2(G179), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n430), .B1(new_n429), .B2(new_n414), .ZN(new_n433));
  AOI211_X1 g0233(.A(KEYINPUT13), .B(new_n413), .C1(new_n428), .C2(new_n420), .ZN(new_n434));
  OAI21_X1  g0234(.A(G169), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n432), .B1(new_n435), .B2(KEYINPUT14), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT14), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n426), .A2(new_n431), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n437), .B1(new_n438), .B2(G169), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n406), .B1(new_n436), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(G200), .B1(new_n433), .B2(new_n434), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n426), .A2(G190), .A3(new_n431), .ZN(new_n442));
  INV_X1    g0242(.A(new_n406), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n395), .A2(new_n440), .A3(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n288), .B1(G1), .B2(new_n409), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n305), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n222), .ZN(new_n451));
  INV_X1    g0251(.A(G87), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n452), .A2(new_n410), .A3(new_n314), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n222), .B(G68), .C1(new_n356), .C2(new_n357), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT19), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n456), .B1(new_n277), .B2(new_n410), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n454), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n270), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n309), .A2(new_n305), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n459), .A2(new_n460), .A3(KEYINPUT80), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT80), .B1(new_n459), .B2(new_n460), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n449), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT81), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT81), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n465), .B(new_n449), .C1(new_n461), .C2(new_n462), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT78), .ZN(new_n468));
  OAI211_X1 g0268(.A(G244), .B(G1698), .C1(new_n356), .C2(new_n357), .ZN(new_n469));
  OAI211_X1 g0269(.A(G238), .B(new_n246), .C1(new_n356), .C2(new_n357), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G33), .A2(G116), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n253), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n256), .A2(G45), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n252), .A2(G250), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(G45), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(G1), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n252), .A2(G274), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n473), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n323), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n473), .A2(new_n267), .A3(new_n480), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n468), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n479), .B1(new_n253), .B2(new_n472), .ZN(new_n485));
  AOI21_X1  g0285(.A(KEYINPUT78), .B1(new_n485), .B2(new_n267), .ZN(new_n486));
  OAI21_X1  g0286(.A(KEYINPUT79), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n483), .B1(G169), .B2(new_n485), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n486), .B1(new_n488), .B2(KEYINPUT78), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT79), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n467), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n485), .A2(G190), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT82), .ZN(new_n494));
  XNOR2_X1  g0294(.A(new_n493), .B(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n459), .A2(new_n460), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT80), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n459), .A2(new_n460), .A3(KEYINPUT80), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n447), .A2(G87), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n481), .A2(G200), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  OR2_X1    g0303(.A1(new_n495), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n492), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(G107), .B1(new_n359), .B2(new_n361), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n410), .A2(new_n314), .A3(KEYINPUT6), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT6), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G97), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n314), .A2(KEYINPUT73), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT73), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G107), .ZN(new_n512));
  AND4_X1   g0312(.A1(new_n507), .A2(new_n509), .A3(new_n510), .A4(new_n512), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n507), .A2(new_n509), .B1(new_n510), .B2(new_n512), .ZN(new_n514));
  OAI21_X1  g0314(.A(G20), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n279), .A2(G77), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n506), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n270), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n294), .A2(G97), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n520), .B1(new_n446), .B2(new_n410), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT77), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n521), .B1(new_n517), .B2(new_n270), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(KEYINPUT77), .ZN(new_n527));
  OAI211_X1 g0327(.A(G244), .B(new_n246), .C1(new_n356), .C2(new_n357), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT74), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT4), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n530), .B1(new_n528), .B2(new_n529), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(G250), .B(G1698), .C1(new_n356), .C2(new_n357), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT75), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT75), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n245), .A2(new_n537), .A3(G250), .A4(G1698), .ZN(new_n538));
  NAND2_X1  g0338(.A1(G33), .A2(G283), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n252), .B1(new_n534), .B2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(G41), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n542), .A2(KEYINPUT76), .A3(KEYINPUT5), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT5), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT76), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n544), .B1(new_n545), .B2(G41), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n342), .A2(new_n477), .A3(new_n543), .A4(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n546), .A2(new_n477), .A3(new_n543), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n252), .ZN(new_n549));
  INV_X1    g0349(.A(G257), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n547), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(G169), .B1(new_n541), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n528), .A2(new_n529), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT4), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n535), .A2(KEYINPUT75), .B1(G33), .B2(G283), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n554), .A2(new_n538), .A3(new_n555), .A4(new_n531), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n551), .B1(new_n556), .B2(new_n253), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G179), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n525), .A2(new_n527), .B1(new_n552), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n526), .B1(new_n557), .B2(new_n333), .ZN(new_n560));
  NOR3_X1   g0360(.A1(new_n541), .A2(new_n347), .A3(new_n551), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(G264), .B(G1698), .C1(new_n356), .C2(new_n357), .ZN(new_n564));
  OAI211_X1 g0364(.A(G257), .B(new_n246), .C1(new_n356), .C2(new_n357), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n243), .A2(G303), .A3(new_n244), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n253), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n548), .A2(G270), .A3(new_n252), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n568), .A2(new_n547), .A3(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(G116), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n295), .A2(new_n298), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n571), .B1(new_n256), .B2(G33), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n271), .B(new_n573), .C1(new_n308), .C2(new_n297), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n269), .A2(new_n221), .B1(G20), .B2(new_n571), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n539), .B(new_n222), .C1(G33), .C2(new_n410), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n575), .A2(KEYINPUT20), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(KEYINPUT20), .B1(new_n575), .B2(new_n576), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n572), .B(new_n574), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n570), .A2(new_n579), .A3(G169), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT21), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n570), .A2(new_n579), .A3(KEYINPUT21), .A4(G169), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n569), .A2(new_n547), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n579), .A2(new_n584), .A3(G179), .A4(new_n568), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n547), .ZN(new_n587));
  OAI211_X1 g0387(.A(G257), .B(G1698), .C1(new_n356), .C2(new_n357), .ZN(new_n588));
  OAI211_X1 g0388(.A(G250), .B(new_n246), .C1(new_n356), .C2(new_n357), .ZN(new_n589));
  INV_X1    g0389(.A(G294), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n588), .B(new_n589), .C1(new_n409), .C2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(G264), .ZN(new_n592));
  OAI21_X1  g0392(.A(KEYINPUT84), .B1(new_n549), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT84), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n548), .A2(new_n594), .A3(G264), .A4(new_n252), .ZN(new_n595));
  AOI221_X4 g0395(.A(new_n587), .B1(new_n591), .B2(new_n253), .C1(new_n593), .C2(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n222), .B(G87), .C1(new_n356), .C2(new_n357), .ZN(new_n597));
  AND2_X1   g0397(.A1(KEYINPUT83), .A2(KEYINPUT22), .ZN(new_n598));
  NOR2_X1   g0398(.A1(KEYINPUT83), .A2(KEYINPUT22), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n245), .A2(new_n222), .A3(G87), .A4(new_n598), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n471), .A2(G20), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT23), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n604), .B1(new_n222), .B2(G107), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n314), .A2(KEYINPUT23), .A3(G20), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n603), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n601), .A2(new_n602), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(KEYINPUT24), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT24), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n601), .A2(new_n602), .A3(new_n610), .A4(new_n607), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n271), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(KEYINPUT25), .B1(new_n287), .B2(new_n314), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n287), .A2(KEYINPUT25), .A3(new_n314), .ZN(new_n614));
  OAI22_X1  g0414(.A1(new_n446), .A2(new_n314), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI22_X1  g0415(.A1(new_n596), .A2(G169), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n593), .A2(new_n595), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n591), .A2(new_n253), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n617), .A2(new_n547), .A3(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n619), .A2(G179), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n582), .B(new_n586), .C1(new_n616), .C2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n609), .A2(new_n611), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n615), .B1(new_n623), .B2(new_n270), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n619), .A2(G200), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n593), .A2(new_n595), .B1(new_n253), .B2(new_n591), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n626), .A2(G190), .A3(new_n547), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n624), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n579), .B1(new_n570), .B2(G200), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(new_n347), .B2(new_n570), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n563), .A2(new_n622), .A3(new_n631), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n445), .A2(new_n505), .A3(new_n632), .ZN(G372));
  OR2_X1    g0433(.A1(new_n336), .A2(new_n337), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n380), .A2(new_n393), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n324), .A2(new_n325), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n444), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n635), .B1(new_n440), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n389), .A2(new_n392), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n634), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n640), .A2(new_n292), .ZN(new_n641));
  INV_X1    g0441(.A(new_n445), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT26), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n495), .A2(new_n503), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n466), .A2(new_n464), .B1(new_n489), .B2(new_n490), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n644), .B1(new_n645), .B2(new_n487), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n643), .B1(new_n646), .B2(new_n559), .ZN(new_n647));
  INV_X1    g0447(.A(new_n488), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n465), .B1(new_n500), .B2(new_n449), .ZN(new_n649));
  INV_X1    g0449(.A(new_n466), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n500), .A2(new_n501), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n502), .A2(new_n493), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n526), .B1(new_n552), .B2(new_n558), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n651), .A2(new_n643), .A3(new_n654), .A4(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n526), .A2(KEYINPUT77), .ZN(new_n657));
  AOI211_X1 g0457(.A(new_n524), .B(new_n521), .C1(new_n270), .C2(new_n517), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n557), .A2(new_n323), .ZN(new_n659));
  AOI211_X1 g0459(.A(new_n267), .B(new_n551), .C1(new_n556), .C2(new_n253), .ZN(new_n660));
  OAI22_X1  g0460(.A1(new_n657), .A2(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n557), .A2(G190), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n662), .B(new_n526), .C1(new_n333), .C2(new_n557), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n621), .A2(new_n661), .A3(new_n663), .A4(new_n628), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n651), .A2(new_n654), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n651), .B(new_n656), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n642), .B1(new_n647), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n641), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n668), .B(KEYINPUT85), .ZN(G369));
  NAND2_X1  g0469(.A1(new_n586), .A2(new_n582), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n293), .A2(new_n222), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(G213), .A3(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(G343), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n579), .ZN(new_n677));
  XOR2_X1   g0477(.A(new_n670), .B(new_n677), .Z(new_n678));
  NAND3_X1  g0478(.A1(new_n678), .A2(G330), .A3(new_n630), .ZN(new_n679));
  INV_X1    g0479(.A(new_n676), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n628), .B1(new_n624), .B2(new_n680), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n616), .A2(new_n620), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n616), .A2(new_n620), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n680), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n679), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n670), .A2(new_n680), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  AOI22_X1  g0490(.A1(new_n683), .A2(new_n690), .B1(new_n684), .B2(new_n680), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n688), .A2(new_n691), .ZN(G399));
  INV_X1    g0492(.A(new_n208), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(G41), .ZN(new_n694));
  OR4_X1    g0494(.A1(new_n256), .A2(new_n694), .A3(G116), .A4(new_n453), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n224), .A2(G50), .ZN(new_n696));
  INV_X1    g0496(.A(new_n694), .ZN(new_n697));
  OAI211_X1 g0497(.A(new_n695), .B(KEYINPUT86), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(KEYINPUT86), .B2(new_n695), .ZN(new_n699));
  XOR2_X1   g0499(.A(new_n699), .B(KEYINPUT28), .Z(new_n700));
  INV_X1    g0500(.A(G330), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n570), .A2(new_n481), .A3(new_n267), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n702), .A2(new_n626), .A3(new_n557), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT87), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(KEYINPUT30), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n557), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n485), .A2(G179), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n707), .A2(new_n570), .A3(new_n619), .A4(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n705), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n702), .A2(new_n626), .A3(new_n557), .A4(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n706), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n712), .A2(KEYINPUT31), .A3(new_n676), .ZN(new_n713));
  AOI21_X1  g0513(.A(KEYINPUT31), .B1(new_n712), .B2(new_n676), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AND4_X1   g0515(.A1(new_n661), .A2(new_n663), .A3(new_n630), .A4(new_n628), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n716), .A2(new_n646), .A3(new_n622), .A4(new_n680), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n701), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(KEYINPUT88), .B1(new_n664), .B2(new_n665), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n624), .A2(new_n625), .A3(new_n627), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n559), .A2(new_n562), .A3(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT88), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n488), .B1(new_n464), .B2(new_n466), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n652), .A2(new_n653), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n721), .A2(new_n722), .A3(new_n621), .A4(new_n725), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n719), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n651), .A2(new_n654), .A3(new_n655), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(KEYINPUT26), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n492), .A2(new_n643), .A3(new_n504), .A4(new_n559), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n729), .A2(new_n651), .A3(new_n730), .ZN(new_n731));
  OAI211_X1 g0531(.A(KEYINPUT29), .B(new_n680), .C1(new_n727), .C2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n680), .B1(new_n666), .B2(new_n647), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT29), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n718), .B1(new_n732), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n700), .B1(new_n736), .B2(G1), .ZN(G364));
  NOR2_X1   g0537(.A1(G13), .A2(G33), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(G20), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n221), .B1(G20), .B2(new_n323), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n693), .A2(new_n245), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(G45), .B2(new_n696), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n744), .B1(G45), .B2(new_n241), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n208), .A2(G355), .A3(new_n245), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(G116), .B2(new_n208), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n742), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n286), .A2(G20), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G45), .ZN(new_n750));
  OR2_X1    g0550(.A1(new_n750), .A2(KEYINPUT89), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n256), .B1(new_n750), .B2(KEYINPUT89), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n694), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n748), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n222), .A2(new_n267), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G190), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G200), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(G322), .ZN(new_n760));
  NOR4_X1   g0560(.A1(new_n222), .A2(new_n267), .A3(new_n333), .A4(G190), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  XOR2_X1   g0562(.A(KEYINPUT33), .B(G317), .Z(new_n763));
  OAI22_X1  g0563(.A1(new_n759), .A2(new_n760), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT95), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n757), .A2(new_n333), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G179), .A2(G200), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n222), .B1(new_n767), .B2(G190), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n766), .A2(G326), .B1(G294), .B2(new_n769), .ZN(new_n770));
  XOR2_X1   g0570(.A(new_n770), .B(KEYINPUT94), .Z(new_n771));
  NAND3_X1  g0571(.A1(new_n756), .A2(new_n347), .A3(new_n333), .ZN(new_n772));
  INV_X1    g0572(.A(G311), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n358), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n333), .A2(G179), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n775), .A2(G20), .A3(G190), .ZN(new_n776));
  OR2_X1    g0576(.A1(new_n776), .A2(KEYINPUT92), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(KEYINPUT92), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n774), .B1(new_n780), .B2(G303), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT90), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n782), .B1(new_n222), .B2(G190), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n347), .A2(KEYINPUT90), .A3(G20), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n783), .A2(new_n784), .A3(new_n775), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n783), .A2(new_n784), .A3(new_n767), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI22_X1  g0588(.A1(G283), .A2(new_n786), .B1(new_n788), .B2(G329), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n765), .A2(new_n771), .A3(new_n781), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n780), .A2(G87), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n791), .B(new_n245), .C1(new_n314), .C2(new_n785), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n792), .B(KEYINPUT93), .Z(new_n793));
  XOR2_X1   g0593(.A(KEYINPUT91), .B(G159), .Z(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n788), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT32), .ZN(new_n797));
  INV_X1    g0597(.A(new_n772), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n798), .A2(G77), .B1(new_n761), .B2(G68), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(new_n272), .B2(new_n759), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n769), .A2(G97), .ZN(new_n801));
  INV_X1    g0601(.A(new_n766), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n801), .B1(new_n802), .B2(new_n202), .ZN(new_n803));
  OR3_X1    g0603(.A1(new_n797), .A2(new_n800), .A3(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n790), .B1(new_n793), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n755), .B1(new_n805), .B2(new_n741), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n678), .A2(new_n630), .ZN(new_n807));
  INV_X1    g0607(.A(new_n740), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT96), .ZN(new_n810));
  INV_X1    g0610(.A(new_n679), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(new_n754), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(G330), .B2(new_n807), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n810), .A2(new_n813), .ZN(G396));
  INV_X1    g0614(.A(new_n311), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n321), .B(new_n815), .C1(new_n347), .C2(new_n318), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n311), .A2(new_n676), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n816), .A2(new_n817), .B1(new_n325), .B2(new_n324), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n324), .A2(new_n325), .A3(new_n680), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(KEYINPUT99), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT99), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n320), .A2(new_n321), .B1(new_n311), .B2(new_n676), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n822), .B(new_n819), .C1(new_n823), .C2(new_n636), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n733), .A2(new_n825), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n821), .A2(new_n824), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n680), .B(new_n827), .C1(new_n666), .C2(new_n647), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NOR3_X1   g0629(.A1(new_n632), .A2(new_n505), .A3(new_n676), .ZN(new_n830));
  INV_X1    g0630(.A(new_n714), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n712), .A2(KEYINPUT31), .A3(new_n676), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(G330), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n754), .B1(new_n829), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n834), .B2(new_n829), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n741), .A2(new_n738), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n754), .B1(G77), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(G303), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n801), .B1(new_n759), .B2(new_n590), .C1(new_n840), .C2(new_n802), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n779), .A2(new_n314), .B1(new_n773), .B2(new_n787), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n785), .A2(new_n452), .ZN(new_n843));
  INV_X1    g0643(.A(G283), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n358), .B1(new_n571), .B2(new_n772), .C1(new_n762), .C2(new_n844), .ZN(new_n845));
  OR4_X1    g0645(.A1(new_n841), .A2(new_n842), .A3(new_n843), .A4(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT97), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n786), .A2(G68), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n779), .B2(new_n202), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n798), .A2(new_n795), .B1(new_n761), .B2(G150), .ZN(new_n851));
  INV_X1    g0651(.A(G143), .ZN(new_n852));
  INV_X1    g0652(.A(G137), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n851), .B1(new_n759), .B2(new_n852), .C1(new_n853), .C2(new_n802), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT34), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n847), .A2(new_n850), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n855), .B2(new_n854), .ZN(new_n857));
  INV_X1    g0657(.A(G132), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n245), .B1(new_n787), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT98), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n859), .A2(new_n860), .B1(G58), .B2(new_n769), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n861), .B1(new_n860), .B2(new_n859), .C1(new_n850), .C2(new_n847), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n846), .B1(new_n857), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n839), .B1(new_n863), .B2(new_n741), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n827), .B2(new_n739), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n836), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(G384));
  NOR2_X1   g0667(.A1(new_n749), .A2(new_n256), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n732), .A2(new_n642), .A3(new_n735), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n641), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT102), .ZN(new_n871));
  OR2_X1    g0671(.A1(new_n383), .A2(KEYINPUT16), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n376), .B1(new_n872), .B2(new_n384), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n378), .B1(new_n873), .B2(new_n674), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n873), .A2(new_n388), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT37), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n390), .A2(new_n387), .ZN(new_n877));
  INV_X1    g0677(.A(new_n674), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n390), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT37), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n877), .A2(new_n879), .A3(new_n880), .A4(new_n378), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n876), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n873), .A2(new_n674), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n394), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT38), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n882), .A2(new_n884), .A3(KEYINPUT38), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n828), .A2(new_n819), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n406), .A2(new_n676), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n440), .A2(new_n444), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n435), .A2(KEYINPUT14), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n438), .A2(new_n437), .A3(G169), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n894), .A2(new_n895), .A3(new_n432), .ZN(new_n896));
  INV_X1    g0696(.A(new_n444), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n406), .B(new_n676), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n891), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n890), .B1(new_n900), .B2(KEYINPUT101), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n828), .A2(new_n819), .B1(new_n893), .B2(new_n898), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT101), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n639), .A2(new_n674), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT39), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n882), .A2(new_n884), .A3(KEYINPUT38), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n877), .A2(new_n879), .A3(new_n378), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT37), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n881), .ZN(new_n911));
  INV_X1    g0711(.A(new_n879), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n394), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT38), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n907), .B1(new_n908), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n887), .A2(KEYINPUT39), .A3(new_n888), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n896), .A2(new_n406), .A3(new_n680), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n905), .A2(new_n906), .A3(new_n921), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n871), .B(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT103), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n825), .B1(new_n715), .B2(new_n717), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n899), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(KEYINPUT40), .B1(new_n908), .B2(new_n914), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n924), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT40), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n911), .A2(new_n913), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n886), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n929), .B1(new_n931), .B2(new_n888), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n932), .A2(KEYINPUT103), .A3(new_n899), .A4(new_n925), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n889), .A2(new_n899), .A3(new_n925), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n928), .A2(new_n933), .B1(new_n929), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n445), .B1(new_n717), .B2(new_n715), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n701), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n935), .B2(new_n936), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n868), .B1(new_n923), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n923), .B2(new_n938), .ZN(new_n940));
  OAI21_X1  g0740(.A(KEYINPUT35), .B1(new_n513), .B2(new_n514), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n941), .A2(G116), .A3(new_n223), .ZN(new_n942));
  NOR3_X1   g0742(.A1(new_n513), .A2(new_n514), .A3(KEYINPUT35), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n944), .B(KEYINPUT36), .Z(new_n945));
  OR3_X1    g0745(.A1(new_n696), .A2(new_n249), .A3(new_n351), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n350), .A2(G50), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT100), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n949), .A2(G1), .A3(new_n286), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n940), .A2(new_n945), .A3(new_n950), .ZN(G367));
  NOR3_X1   g0751(.A1(new_n693), .A2(new_n234), .A3(new_n245), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n742), .B1(new_n208), .B2(new_n305), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n754), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n780), .A2(KEYINPUT46), .A3(G116), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT46), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n779), .B2(new_n571), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n955), .B(new_n957), .C1(new_n590), .C2(new_n762), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT110), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n759), .A2(new_n840), .B1(new_n802), .B2(new_n773), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n358), .B1(new_n768), .B2(new_n314), .C1(new_n772), .C2(new_n844), .ZN(new_n961));
  INV_X1    g0761(.A(G317), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n787), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n785), .A2(new_n410), .ZN(new_n964));
  NOR4_X1   g0764(.A1(new_n960), .A2(new_n961), .A3(new_n963), .A4(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n786), .A2(G77), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n853), .B2(new_n787), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(new_n780), .B2(G58), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n762), .A2(new_n794), .B1(new_n772), .B2(new_n202), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT111), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n768), .A2(new_n350), .ZN(new_n971));
  INV_X1    g0771(.A(G150), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n759), .A2(new_n972), .B1(new_n802), .B2(new_n852), .ZN(new_n973));
  NOR4_X1   g0773(.A1(new_n970), .A2(new_n358), .A3(new_n971), .A4(new_n973), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n959), .A2(new_n965), .B1(new_n968), .B2(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT47), .Z(new_n976));
  AOI21_X1  g0776(.A(new_n954), .B1(new_n976), .B2(new_n741), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT104), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n680), .B1(new_n500), .B2(new_n501), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n723), .A2(new_n979), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n978), .B(new_n980), .C1(new_n665), .C2(new_n979), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n723), .A2(KEYINPUT104), .A3(new_n979), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n977), .B1(new_n808), .B2(new_n984), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n683), .A2(new_n685), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n690), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n686), .A2(new_n689), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n811), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n987), .A2(new_n679), .A3(new_n988), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n719), .A2(new_n726), .ZN(new_n993));
  AND3_X1   g0793(.A1(new_n729), .A2(new_n651), .A3(new_n730), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n734), .B(new_n676), .C1(new_n993), .C2(new_n994), .ZN(new_n995));
  AND2_X1   g0795(.A1(new_n733), .A2(new_n734), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n992), .B(new_n834), .C1(new_n995), .C2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT106), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT107), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n736), .A2(KEYINPUT106), .A3(new_n992), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT45), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n563), .B1(new_n526), .B2(new_n680), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n655), .A2(new_n676), .ZN(new_n1005));
  AND2_X1   g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n691), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1003), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1009), .A2(KEYINPUT45), .A3(new_n691), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1006), .A2(KEYINPUT44), .A3(new_n1007), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT44), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n1009), .B2(new_n691), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n688), .B1(new_n1011), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT108), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1011), .A2(new_n1015), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1017), .B1(new_n1018), .B2(new_n687), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1011), .A2(new_n1015), .A3(KEYINPUT108), .A4(new_n688), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1016), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1002), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1000), .B1(new_n999), .B2(new_n1001), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n736), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n694), .B(KEYINPUT41), .Z(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(KEYINPUT109), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT109), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1024), .A2(new_n1029), .A3(new_n1026), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n753), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n687), .A2(new_n1009), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT105), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1033), .B(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1006), .A2(new_n987), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n1038), .A2(KEYINPUT42), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT42), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n559), .B1(new_n1009), .B2(new_n684), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n1037), .A2(new_n1040), .B1(new_n1041), .B2(new_n676), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1036), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1035), .B(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n985), .B1(new_n1031), .B2(new_n1045), .ZN(G387));
  NAND2_X1  g0846(.A1(new_n992), .A2(new_n753), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n780), .A2(G294), .B1(G283), .B2(new_n769), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n798), .A2(G303), .B1(new_n761), .B2(G311), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(new_n759), .B2(new_n962), .C1(new_n760), .C2(new_n802), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT48), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1048), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT112), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT49), .Z(new_n1056));
  AOI21_X1  g0856(.A(new_n245), .B1(new_n788), .B2(G326), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n571), .B2(new_n785), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n769), .A2(new_n448), .ZN(new_n1060));
  INV_X1    g0860(.A(G159), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1060), .B1(new_n759), .B2(new_n202), .C1(new_n1061), .C2(new_n802), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n779), .A2(new_n249), .B1(new_n972), .B2(new_n787), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n245), .B1(new_n350), .B2(new_n772), .C1(new_n762), .C2(new_n302), .ZN(new_n1064));
  NOR4_X1   g0864(.A1(new_n1062), .A2(new_n1063), .A3(new_n964), .A4(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n741), .B1(new_n1059), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n754), .ZN(new_n1067));
  NOR3_X1   g0867(.A1(new_n231), .A2(new_n476), .A3(new_n245), .ZN(new_n1068));
  OR3_X1    g0868(.A1(new_n302), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1069));
  OAI21_X1  g0869(.A(KEYINPUT50), .B1(new_n302), .B2(G50), .ZN(new_n1070));
  AOI21_X1  g0870(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  AOI211_X1 g0872(.A(G116), .B(new_n453), .C1(new_n1072), .C2(new_n358), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n208), .B1(new_n1068), .B2(new_n1073), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n740), .B(new_n741), .C1(new_n693), .C2(G107), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1067), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1066), .B(new_n1076), .C1(new_n986), .C2(new_n808), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n999), .A2(new_n1001), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n694), .B1(new_n736), .B2(new_n992), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1047), .B(new_n1077), .C1(new_n1079), .C2(new_n1080), .ZN(G393));
  XNOR2_X1  g0881(.A(new_n1016), .B(KEYINPUT113), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n697), .B1(new_n1084), .B2(new_n1078), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1078), .A2(KEYINPUT107), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1086), .A2(new_n1002), .A3(new_n1021), .ZN(new_n1087));
  AND2_X1   g0887(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n743), .A2(new_n238), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n742), .B1(new_n208), .B2(new_n410), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n754), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n358), .B1(new_n590), .B2(new_n772), .C1(new_n762), .C2(new_n840), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(G116), .B2(new_n769), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n780), .A2(G283), .B1(G107), .B2(new_n786), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1093), .B(new_n1094), .C1(new_n760), .C2(new_n787), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(G311), .A2(new_n758), .B1(new_n766), .B2(G317), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT52), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n798), .A2(new_n276), .B1(new_n761), .B2(G50), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT114), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n780), .A2(G68), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1098), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n1101), .A2(KEYINPUT114), .B1(new_n788), .B2(G143), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n358), .B(new_n843), .C1(G77), .C2(new_n769), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1100), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(G150), .A2(new_n766), .B1(new_n758), .B2(G159), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT51), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n1095), .A2(new_n1097), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1091), .B1(new_n1107), .B2(new_n741), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n1009), .B2(new_n808), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n753), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1109), .B1(new_n1084), .B2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1088), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(G390));
  AND2_X1   g0913(.A1(new_n893), .A2(new_n898), .ZN(new_n1114));
  OAI211_X1 g0914(.A(G330), .B(new_n827), .C1(new_n830), .C2(new_n833), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n920), .B1(new_n931), .B2(new_n888), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n680), .B(new_n827), .C1(new_n727), .C2(new_n731), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n819), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1118), .B1(new_n1120), .B2(new_n899), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n900), .A2(new_n919), .B1(new_n915), .B2(new_n916), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1116), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n676), .B1(new_n993), .B2(new_n994), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n820), .B1(new_n1124), .B2(new_n827), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1117), .B1(new_n1125), .B2(new_n1114), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n917), .B1(new_n902), .B2(new_n920), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT115), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n701), .B(new_n825), .C1(new_n715), .C2(new_n717), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1130), .A2(KEYINPUT115), .A3(new_n899), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1126), .A2(new_n1127), .A3(new_n1129), .A4(new_n1131), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1123), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n753), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1067), .B1(new_n302), .B2(new_n837), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n741), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n358), .B1(new_n768), .B2(new_n249), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n791), .B(new_n848), .C1(new_n590), .C2(new_n787), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n1137), .B(new_n1138), .C1(G116), .C2(new_n758), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n798), .A2(G97), .B1(new_n761), .B2(G107), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n844), .B2(new_n802), .ZN(new_n1141));
  XOR2_X1   g0941(.A(new_n1141), .B(KEYINPUT118), .Z(new_n1142));
  NOR2_X1   g0942(.A1(new_n779), .A2(new_n972), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT53), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n766), .A2(G128), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n1145), .B1(new_n1061), .B2(new_n768), .C1(new_n759), .C2(new_n858), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(KEYINPUT54), .B(G143), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n245), .B1(new_n772), .B2(new_n1147), .C1(new_n762), .C2(new_n853), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n788), .A2(G125), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n785), .A2(new_n202), .ZN(new_n1150));
  NOR4_X1   g0950(.A1(new_n1146), .A2(new_n1148), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1139), .A2(new_n1142), .B1(new_n1144), .B2(new_n1151), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1135), .B1(new_n1136), .B2(new_n1152), .C1(new_n918), .C2(new_n739), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1129), .A2(new_n1125), .A3(new_n1131), .A4(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1130), .A2(new_n899), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n891), .B1(new_n1116), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(KEYINPUT116), .B1(new_n834), .B2(new_n445), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT116), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n642), .A2(new_n1160), .A3(new_n718), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  AND3_X1   g0962(.A1(new_n1162), .A2(new_n641), .A3(new_n869), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1123), .A2(new_n1132), .A3(new_n1158), .A4(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n694), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT117), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1162), .A2(new_n641), .A3(new_n869), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(new_n1157), .B2(new_n1155), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n1165), .A2(new_n1166), .B1(new_n1133), .B2(new_n1170), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1134), .B(new_n1153), .C1(new_n1168), .C2(new_n1171), .ZN(G378));
  NAND2_X1  g0972(.A1(new_n634), .A2(new_n292), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n291), .A2(new_n878), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n1174), .B(KEYINPUT121), .Z(new_n1175));
  XNOR2_X1  g0975(.A(new_n1173), .B(new_n1175), .ZN(new_n1176));
  XOR2_X1   g0976(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1176), .B(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n738), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n754), .B1(G50), .B2(new_n838), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n802), .A2(new_n571), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n971), .B(new_n1183), .C1(G107), .C2(new_n758), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n245), .A2(G41), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1185), .B1(new_n305), .B2(new_n772), .C1(new_n762), .C2(new_n410), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(G77), .B2(new_n780), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1184), .B(new_n1187), .C1(new_n844), .C2(new_n787), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n786), .A2(G58), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1189), .B(KEYINPUT119), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT120), .ZN(new_n1192));
  OR2_X1    g0992(.A1(new_n1192), .A2(KEYINPUT58), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(KEYINPUT58), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(G33), .A2(G41), .ZN(new_n1195));
  NOR3_X1   g0995(.A1(new_n1185), .A2(G50), .A3(new_n1195), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n762), .A2(new_n858), .B1(new_n772), .B2(new_n853), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G150), .B2(new_n769), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(G125), .A2(new_n766), .B1(new_n758), .B2(G128), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1198), .B(new_n1199), .C1(new_n779), .C2(new_n1147), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1200), .A2(KEYINPUT59), .ZN(new_n1201));
  INV_X1    g1001(.A(G124), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1195), .B1(new_n787), .B2(new_n1202), .C1(new_n785), .C2(new_n794), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n1200), .B2(KEYINPUT59), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1196), .B1(new_n1201), .B2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1193), .A2(new_n1194), .A3(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1182), .B1(new_n1206), .B2(new_n741), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1181), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n928), .A2(new_n933), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n701), .B1(new_n934), .B2(new_n929), .ZN(new_n1211));
  AND3_X1   g1011(.A1(new_n1210), .A2(new_n1211), .A3(new_n1179), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1179), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n922), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n1180), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n906), .B1(new_n917), .B2(new_n919), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n901), .B2(new_n904), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1210), .A2(new_n1211), .A3(new_n1179), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1216), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1214), .A2(new_n1220), .A3(KEYINPUT122), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(KEYINPUT122), .B1(new_n1214), .B2(new_n1220), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1209), .B1(new_n1224), .B2(new_n753), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1164), .A2(new_n1163), .ZN(new_n1226));
  AOI21_X1  g1026(.A(KEYINPUT57), .B1(new_n1224), .B2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT57), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(new_n1164), .B2(new_n1163), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1214), .A2(new_n1220), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n694), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1225), .B1(new_n1227), .B2(new_n1232), .ZN(G375));
  NAND2_X1  g1033(.A1(new_n1114), .A2(new_n738), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n754), .B1(G68), .B2(new_n838), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n358), .B1(new_n314), .B2(new_n772), .C1(new_n762), .C2(new_n571), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(G77), .B2(new_n786), .ZN(new_n1237));
  OAI221_X1 g1037(.A(new_n1237), .B1(new_n410), .B2(new_n779), .C1(new_n840), .C2(new_n787), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1060), .B1(new_n759), .B2(new_n844), .C1(new_n590), .C2(new_n802), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n245), .B1(new_n772), .B2(new_n972), .C1(new_n762), .C2(new_n1147), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(G128), .B2(new_n788), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n802), .A2(new_n858), .B1(new_n768), .B2(new_n202), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(G137), .B2(new_n758), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1241), .B(new_n1243), .C1(new_n1061), .C2(new_n779), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n1238), .A2(new_n1239), .B1(new_n1244), .B2(new_n1190), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1235), .B1(new_n1245), .B2(new_n741), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n1158), .A2(new_n753), .B1(new_n1234), .B2(new_n1246), .ZN(new_n1247));
  OR2_X1    g1047(.A1(new_n1170), .A2(new_n1025), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1158), .A2(new_n1163), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1247), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1250), .B(KEYINPUT123), .ZN(G381));
  OR2_X1    g1051(.A1(G393), .A2(G396), .ZN(new_n1252));
  NOR4_X1   g1052(.A1(G381), .A2(G390), .A3(G384), .A4(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1134), .A2(new_n1153), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1171), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1254), .B1(new_n1255), .B2(new_n1167), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1253), .A2(new_n1256), .ZN(new_n1257));
  OR3_X1    g1057(.A1(new_n1257), .A2(G387), .A3(G375), .ZN(G407));
  NAND2_X1  g1058(.A1(new_n1256), .A2(new_n675), .ZN(new_n1259));
  OAI211_X1 g1059(.A(G407), .B(G213), .C1(G375), .C2(new_n1259), .ZN(G409));
  XOR2_X1   g1060(.A(G393), .B(G396), .Z(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n1024), .A2(new_n1029), .A3(new_n1026), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1029), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1110), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1044), .ZN(new_n1266));
  AOI21_X1  g1066(.A(G390), .B1(new_n1266), .B2(new_n985), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n985), .ZN(new_n1268));
  AOI211_X1 g1068(.A(new_n1268), .B(new_n1112), .C1(new_n1265), .C2(new_n1044), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1262), .B1(new_n1267), .B2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(G387), .A2(new_n1112), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1266), .A2(new_n985), .A3(G390), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1271), .A2(new_n1261), .A3(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1270), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT60), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1275), .B1(new_n1158), .B2(new_n1163), .ZN(new_n1276));
  OAI21_X1  g1076(.A(KEYINPUT124), .B1(new_n1276), .B2(new_n1249), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT124), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1169), .A2(new_n1157), .A3(new_n1155), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n1278), .B(new_n1279), .C1(new_n1170), .C2(new_n1275), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n697), .B1(new_n1249), .B2(KEYINPUT60), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1277), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1247), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n866), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1282), .A2(G384), .A3(new_n1247), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(G213), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1288), .A2(G343), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT122), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(new_n922), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1218), .B1(new_n1216), .B2(new_n1219), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1291), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1294), .A2(new_n1226), .A3(new_n1221), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1232), .B1(new_n1228), .B2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1294), .A2(new_n753), .A3(new_n1221), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1208), .ZN(new_n1298));
  NOR3_X1   g1098(.A1(new_n1296), .A2(new_n1256), .A3(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1224), .A2(new_n1026), .A3(new_n1226), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1209), .B1(new_n1230), .B2(new_n753), .ZN(new_n1301));
  AOI21_X1  g1101(.A(G378), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  OAI211_X1 g1102(.A(new_n1287), .B(new_n1290), .C1(new_n1299), .C2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(KEYINPUT125), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1256), .ZN(new_n1306));
  OAI211_X1 g1106(.A(G378), .B(new_n1225), .C1(new_n1227), .C2(new_n1232), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT125), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1308), .A2(new_n1309), .A3(new_n1287), .A4(new_n1290), .ZN(new_n1310));
  AOI21_X1  g1110(.A(KEYINPUT62), .B1(new_n1304), .B2(new_n1310), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1290), .B1(new_n1299), .B2(new_n1302), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT126), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1289), .A2(G2897), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  AND3_X1   g1115(.A1(new_n1282), .A2(G384), .A3(new_n1247), .ZN(new_n1316));
  AOI21_X1  g1116(.A(G384), .B1(new_n1282), .B2(new_n1247), .ZN(new_n1317));
  OAI211_X1 g1117(.A(new_n1313), .B(new_n1315), .C1(new_n1316), .C2(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1284), .A2(KEYINPUT126), .A3(new_n1285), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1315), .B1(new_n1286), .B2(new_n1313), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(KEYINPUT61), .B1(new_n1312), .B2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1303), .A2(KEYINPUT62), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1274), .B1(new_n1311), .B2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT63), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1304), .A2(new_n1310), .A3(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1274), .ZN(new_n1329));
  OR2_X1    g1129(.A1(new_n1303), .A2(new_n1327), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1328), .A2(new_n1323), .A3(new_n1329), .A4(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1326), .A2(new_n1331), .ZN(G405));
  NAND2_X1  g1132(.A1(new_n1286), .A2(KEYINPUT127), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1270), .A2(new_n1273), .A3(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1333), .B1(new_n1270), .B2(new_n1273), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(G375), .A2(new_n1256), .ZN(new_n1337));
  OR2_X1    g1137(.A1(new_n1286), .A2(KEYINPUT127), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1337), .A2(new_n1307), .A3(new_n1338), .ZN(new_n1339));
  NOR3_X1   g1139(.A1(new_n1335), .A2(new_n1336), .A3(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1339), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1333), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1274), .A2(new_n1342), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1341), .B1(new_n1343), .B2(new_n1334), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1340), .A2(new_n1344), .ZN(G402));
endmodule


