//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 0 1 0 1 1 0 0 1 1 0 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G140), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G227), .ZN(new_n191));
  XOR2_X1   g005(.A(new_n189), .B(new_n191), .Z(new_n192));
  INV_X1    g006(.A(KEYINPUT11), .ZN(new_n193));
  INV_X1    g007(.A(G134), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(G137), .ZN(new_n195));
  INV_X1    g009(.A(G137), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(KEYINPUT11), .A3(G134), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(G137), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n195), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G131), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n195), .A2(new_n197), .A3(new_n201), .A4(new_n198), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT80), .B(G104), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT3), .B1(new_n204), .B2(G107), .ZN(new_n205));
  AOI21_X1  g019(.A(G101), .B1(new_n204), .B2(G107), .ZN(new_n206));
  INV_X1    g020(.A(G104), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(KEYINPUT3), .ZN(new_n208));
  INV_X1    g022(.A(G107), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT81), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT81), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G107), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n208), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT82), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT81), .B(G107), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(KEYINPUT82), .A3(new_n208), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n205), .A2(new_n206), .A3(new_n215), .A4(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n204), .A2(G107), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n216), .A2(G104), .ZN(new_n220));
  OAI21_X1  g034(.A(G101), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G146), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT64), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT64), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G146), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n223), .A2(new_n225), .A3(G143), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n222), .A2(G143), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G128), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n226), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(KEYINPUT64), .B(G146), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n227), .B1(new_n232), .B2(G143), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n222), .A2(G143), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n229), .B1(new_n234), .B2(KEYINPUT1), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n231), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n218), .A2(new_n221), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n229), .B1(new_n226), .B2(KEYINPUT1), .ZN(new_n239));
  INV_X1    g053(.A(new_n234), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n223), .A2(new_n225), .ZN(new_n241));
  INV_X1    g055(.A(G143), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n240), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n231), .B1(new_n239), .B2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n244), .B1(new_n218), .B2(new_n221), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n203), .B1(new_n238), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT12), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT12), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n248), .B(new_n203), .C1(new_n238), .C2(new_n245), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n218), .A2(new_n221), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT10), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n234), .B1(new_n232), .B2(G143), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT1), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n254), .B1(new_n232), .B2(G143), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n253), .B1(new_n255), .B2(new_n229), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n252), .B1(new_n256), .B2(new_n231), .ZN(new_n257));
  AOI22_X1  g071(.A1(new_n251), .A2(new_n257), .B1(new_n237), .B2(new_n252), .ZN(new_n258));
  INV_X1    g072(.A(new_n203), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n204), .A2(G107), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n205), .A2(new_n215), .A3(new_n260), .A4(new_n217), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G101), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n262), .A2(KEYINPUT4), .A3(new_n218), .ZN(new_n263));
  AND2_X1   g077(.A1(KEYINPUT0), .A2(G128), .ZN(new_n264));
  NOR2_X1   g078(.A1(KEYINPUT0), .A2(G128), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n253), .A2(new_n266), .B1(new_n233), .B2(new_n264), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G101), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n269), .A2(KEYINPUT4), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n261), .A2(KEYINPUT83), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(KEYINPUT83), .B1(new_n261), .B2(new_n270), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n258), .B(new_n259), .C1(new_n268), .C2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT84), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n263), .B(new_n267), .C1(new_n272), .C2(new_n271), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT84), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n276), .A2(new_n277), .A3(new_n259), .A4(new_n258), .ZN(new_n278));
  AOI211_X1 g092(.A(new_n192), .B(new_n250), .C1(new_n275), .C2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n192), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n275), .A2(new_n278), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n259), .B1(new_n276), .B2(new_n258), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n280), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n187), .B(new_n188), .C1(new_n279), .C2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(G469), .A2(G902), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n282), .B1(new_n275), .B2(new_n278), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n280), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n250), .B1(new_n275), .B2(new_n278), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n288), .B(G469), .C1(new_n280), .C2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n285), .A2(new_n286), .A3(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(G214), .B1(G237), .B2(G902), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n218), .A2(new_n221), .ZN(new_n294));
  XOR2_X1   g108(.A(KEYINPUT2), .B(G113), .Z(new_n295));
  XNOR2_X1  g109(.A(G116), .B(G119), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n295), .A2(KEYINPUT66), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(KEYINPUT66), .B1(new_n295), .B2(new_n296), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G119), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G116), .ZN(new_n302));
  OAI21_X1  g116(.A(G113), .B1(new_n302), .B2(KEYINPUT5), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n303), .B1(KEYINPUT5), .B2(new_n296), .ZN(new_n304));
  OR3_X1    g118(.A1(new_n294), .A2(new_n300), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n295), .A2(new_n296), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT66), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT65), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n296), .B1(new_n295), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT2), .B(G113), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT65), .ZN(new_n312));
  AOI22_X1  g126(.A1(new_n308), .A2(new_n297), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n263), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n305), .B1(new_n315), .B2(new_n273), .ZN(new_n316));
  XNOR2_X1  g130(.A(G110), .B(G122), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n305), .B(new_n317), .C1(new_n315), .C2(new_n273), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(KEYINPUT6), .A3(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT6), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n316), .A2(new_n322), .A3(new_n318), .ZN(new_n323));
  INV_X1    g137(.A(G125), .ZN(new_n324));
  OR2_X1    g138(.A1(new_n267), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n256), .A2(new_n324), .A3(new_n231), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n190), .A2(G224), .ZN(new_n328));
  XOR2_X1   g142(.A(new_n327), .B(new_n328), .Z(new_n329));
  NAND3_X1  g143(.A1(new_n321), .A2(new_n323), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(KEYINPUT7), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n325), .A2(new_n326), .A3(KEYINPUT7), .A4(new_n328), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  XOR2_X1   g148(.A(new_n317), .B(KEYINPUT8), .Z(new_n335));
  OAI21_X1  g149(.A(new_n294), .B1(new_n300), .B2(new_n304), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n335), .B1(new_n305), .B2(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(G902), .B1(new_n338), .B2(new_n320), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n330), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(G210), .B1(G237), .B2(G902), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n330), .A2(new_n339), .A3(new_n341), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n293), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT9), .B(G234), .ZN(new_n346));
  OAI21_X1  g160(.A(G221), .B1(new_n346), .B2(G902), .ZN(new_n347));
  INV_X1    g161(.A(G475), .ZN(new_n348));
  INV_X1    g162(.A(G140), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G125), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n324), .A2(G140), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n351), .A3(KEYINPUT73), .ZN(new_n352));
  OR3_X1    g166(.A1(new_n324), .A2(KEYINPUT73), .A3(G140), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n352), .A2(new_n353), .A3(KEYINPUT16), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT16), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n350), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G146), .ZN(new_n358));
  INV_X1    g172(.A(G237), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n359), .A2(new_n190), .A3(G214), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n242), .ZN(new_n361));
  NOR2_X1   g175(.A1(G237), .A2(G953), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(G143), .A3(G214), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G131), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT17), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n361), .A2(new_n201), .A3(new_n363), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n354), .A2(new_n222), .A3(new_n356), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n364), .A2(KEYINPUT17), .A3(G131), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n358), .A2(new_n368), .A3(new_n369), .A4(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT85), .ZN(new_n372));
  AND4_X1   g186(.A1(G143), .A2(new_n359), .A3(new_n190), .A4(G214), .ZN(new_n373));
  AOI21_X1  g187(.A(G143), .B1(new_n362), .B2(G214), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(KEYINPUT18), .A2(G131), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n361), .A2(KEYINPUT85), .A3(new_n363), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n375), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n352), .A2(new_n353), .A3(G146), .ZN(new_n380));
  XNOR2_X1  g194(.A(G125), .B(G140), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n232), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n373), .A2(new_n374), .ZN(new_n384));
  AOI21_X1  g198(.A(KEYINPUT86), .B1(new_n384), .B2(new_n376), .ZN(new_n385));
  AND4_X1   g199(.A1(KEYINPUT86), .A2(new_n361), .A3(new_n376), .A4(new_n363), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n379), .B(new_n383), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n371), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(G113), .B(G122), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n389), .B(new_n207), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n371), .A2(new_n390), .A3(new_n387), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n348), .B1(new_n394), .B2(new_n188), .ZN(new_n395));
  INV_X1    g209(.A(G122), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G116), .ZN(new_n397));
  INV_X1    g211(.A(G116), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G122), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n210), .A2(new_n212), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(G116), .B(G122), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n216), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(G128), .B(G143), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n402), .A2(new_n404), .B1(new_n194), .B2(new_n405), .ZN(new_n406));
  OR2_X1    g220(.A1(KEYINPUT88), .A2(KEYINPUT13), .ZN(new_n407));
  NAND2_X1  g221(.A1(KEYINPUT88), .A2(KEYINPUT13), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(new_n405), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n229), .A2(G143), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(new_n407), .A3(new_n408), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n410), .A2(G134), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n406), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n405), .A2(new_n194), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n242), .A2(G128), .ZN(new_n416));
  OAI21_X1  g230(.A(G134), .B1(new_n411), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n398), .A2(KEYINPUT14), .A3(G122), .ZN(new_n419));
  OAI211_X1 g233(.A(G107), .B(new_n419), .C1(new_n400), .C2(KEYINPUT14), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n418), .A2(new_n420), .A3(new_n404), .ZN(new_n421));
  XOR2_X1   g235(.A(KEYINPUT72), .B(G217), .Z(new_n422));
  NOR3_X1   g236(.A1(new_n422), .A2(G953), .A3(new_n346), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n414), .A2(KEYINPUT89), .A3(new_n421), .A4(new_n423), .ZN(new_n424));
  AOI22_X1  g238(.A1(new_n415), .A2(new_n417), .B1(new_n216), .B2(new_n403), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n406), .A2(new_n413), .B1(new_n425), .B2(new_n420), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n424), .B1(new_n426), .B2(new_n423), .ZN(new_n427));
  AOI21_X1  g241(.A(KEYINPUT89), .B1(new_n426), .B2(new_n423), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n188), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G478), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(KEYINPUT15), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  OAI221_X1 g246(.A(new_n188), .B1(KEYINPUT15), .B2(new_n430), .C1(new_n427), .C2(new_n428), .ZN(new_n433));
  INV_X1    g247(.A(G952), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n434), .A2(G953), .ZN(new_n435));
  NAND2_X1  g249(.A1(G234), .A2(G237), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  XOR2_X1   g251(.A(new_n437), .B(KEYINPUT90), .Z(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(G898), .ZN(new_n440));
  XOR2_X1   g254(.A(new_n440), .B(KEYINPUT91), .Z(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n436), .A2(G902), .A3(G953), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n439), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n432), .A2(new_n433), .A3(new_n446), .ZN(new_n447));
  NOR2_X1   g261(.A1(G475), .A2(G902), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT19), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n449), .B1(new_n352), .B2(new_n353), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n381), .A2(KEYINPUT19), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n232), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n365), .A2(new_n367), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n358), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n387), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT87), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(new_n456), .A3(new_n391), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n393), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n456), .B1(new_n455), .B2(new_n391), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n448), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT20), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n455), .A2(new_n391), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT87), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n463), .A2(new_n393), .A3(new_n457), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT20), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n464), .A2(new_n465), .A3(new_n448), .ZN(new_n466));
  AOI211_X1 g280(.A(new_n395), .B(new_n447), .C1(new_n461), .C2(new_n466), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n291), .A2(new_n345), .A3(new_n347), .A4(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT79), .ZN(new_n469));
  NOR2_X1   g283(.A1(G472), .A2(G902), .ZN(new_n470));
  INV_X1    g284(.A(new_n198), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n194), .A2(G137), .ZN(new_n472));
  OAI21_X1  g286(.A(G131), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n202), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n244), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT30), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n253), .A2(new_n266), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n233), .A2(new_n264), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n203), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n476), .A2(new_n477), .A3(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n477), .B1(new_n476), .B2(new_n480), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n314), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n476), .A2(new_n480), .A3(new_n313), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n362), .A2(G210), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(KEYINPUT27), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT26), .B(G101), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n487), .B(new_n488), .ZN(new_n489));
  XOR2_X1   g303(.A(KEYINPUT67), .B(KEYINPUT31), .Z(new_n490));
  NAND4_X1  g304(.A1(new_n484), .A2(new_n485), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n480), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n474), .B1(new_n256), .B2(new_n231), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT30), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n313), .B1(new_n494), .B2(new_n481), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n476), .A2(new_n480), .A3(new_n313), .ZN(new_n496));
  INV_X1    g310(.A(new_n489), .ZN(new_n497));
  NOR3_X1   g311(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT67), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n499), .A2(KEYINPUT31), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n491), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT28), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n314), .B1(new_n492), .B2(new_n493), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n502), .B1(new_n503), .B2(new_n485), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n485), .A2(new_n502), .ZN(new_n505));
  OAI21_X1  g319(.A(KEYINPUT68), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n313), .B1(new_n476), .B2(new_n480), .ZN(new_n507));
  OAI21_X1  g321(.A(KEYINPUT28), .B1(new_n496), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT68), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n489), .B1(new_n506), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n470), .B1(new_n501), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT32), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n485), .A2(new_n502), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n509), .B1(new_n508), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n503), .A2(new_n485), .ZN(new_n516));
  AOI21_X1  g330(.A(KEYINPUT68), .B1(new_n516), .B2(KEYINPUT28), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n497), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n484), .A2(new_n485), .A3(new_n489), .ZN(new_n519));
  INV_X1    g333(.A(new_n500), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n518), .A2(new_n491), .A3(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT32), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n522), .A2(new_n523), .A3(new_n470), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n506), .A2(new_n510), .A3(new_n489), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n494), .A2(new_n481), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n496), .B1(new_n526), .B2(new_n314), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT69), .B1(new_n527), .B2(new_n489), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT29), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT69), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n530), .B(new_n497), .C1(new_n495), .C2(new_n496), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n525), .A2(new_n528), .A3(new_n529), .A4(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n505), .B1(new_n516), .B2(KEYINPUT28), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n497), .A2(new_n529), .ZN(new_n534));
  AOI21_X1  g348(.A(KEYINPUT70), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n508), .A2(KEYINPUT70), .A3(new_n514), .A4(new_n534), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n188), .ZN(new_n537));
  OAI21_X1  g351(.A(KEYINPUT71), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n508), .A2(new_n514), .A3(new_n534), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT70), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT71), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n541), .A2(new_n542), .A3(new_n188), .A4(new_n536), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n532), .A2(new_n538), .A3(new_n543), .ZN(new_n544));
  AOI22_X1  g358(.A1(new_n513), .A2(new_n524), .B1(new_n544), .B2(G472), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n546), .B(KEYINPUT74), .ZN(new_n547));
  XNOR2_X1  g361(.A(KEYINPUT22), .B(G137), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n547), .B(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT23), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n551), .B1(new_n301), .B2(G128), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n229), .A2(KEYINPUT23), .A3(G119), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n552), .B(new_n553), .C1(G119), .C2(new_n229), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(G110), .ZN(new_n555));
  XOR2_X1   g369(.A(KEYINPUT24), .B(G110), .Z(new_n556));
  XNOR2_X1  g370(.A(G119), .B(G128), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n559), .B1(new_n358), .B2(new_n369), .ZN(new_n560));
  OAI22_X1  g374(.A1(new_n554), .A2(G110), .B1(new_n557), .B2(new_n556), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n382), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n222), .B1(new_n354), .B2(new_n356), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n550), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n369), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n558), .B(new_n555), .C1(new_n566), .C2(new_n563), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n358), .A2(new_n382), .A3(new_n561), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n549), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n188), .B1(new_n565), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n570), .A2(KEYINPUT75), .A3(KEYINPUT25), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT25), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n550), .B1(new_n560), .B2(new_n564), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n567), .A2(new_n568), .A3(new_n549), .ZN(new_n574));
  AOI21_X1  g388(.A(G902), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT75), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n572), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n422), .B1(G234), .B2(new_n188), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n571), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n573), .A2(new_n574), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n578), .A2(G902), .ZN(new_n581));
  XOR2_X1   g395(.A(KEYINPUT76), .B(KEYINPUT77), .Z(new_n582));
  XNOR2_X1  g396(.A(new_n581), .B(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT78), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT78), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n579), .A2(new_n587), .A3(new_n584), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n469), .B1(new_n545), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n513), .A2(new_n524), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n544), .A2(G472), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n589), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(KEYINPUT79), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n468), .B1(new_n590), .B2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(new_n269), .ZN(G3));
  INV_X1    g411(.A(G472), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n598), .B1(new_n522), .B2(new_n188), .ZN(new_n599));
  INV_X1    g413(.A(new_n512), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n594), .A2(new_n291), .A3(new_n347), .A4(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n330), .A2(new_n339), .A3(new_n341), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n341), .B1(new_n330), .B2(new_n339), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n292), .B(new_n446), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n395), .B1(new_n461), .B2(new_n466), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  OR2_X1    g422(.A1(new_n427), .A2(new_n428), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT33), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n426), .A2(new_n423), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n426), .A2(new_n423), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n612), .A2(new_n610), .ZN(new_n613));
  AOI22_X1  g427(.A1(new_n609), .A2(new_n610), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n430), .A2(G902), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n614), .A2(new_n615), .B1(new_n430), .B2(new_n429), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n608), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n606), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n603), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(G104), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT92), .B(KEYINPUT34), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G6));
  NAND3_X1  g437(.A1(new_n461), .A2(KEYINPUT93), .A3(new_n466), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT93), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n460), .A2(new_n625), .A3(KEYINPUT20), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n395), .B1(new_n432), .B2(new_n433), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n624), .A2(new_n626), .A3(new_n446), .A4(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT94), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n292), .B1(new_n604), .B2(new_n605), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n628), .A2(new_n629), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n603), .A2(new_n630), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT95), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT35), .B(G107), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G9));
  OAI211_X1 g451(.A(new_n467), .B(new_n292), .C1(new_n604), .C2(new_n605), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n567), .A2(new_n568), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n549), .A2(KEYINPUT36), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n583), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n579), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n599), .A2(new_n600), .A3(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n639), .A2(new_n347), .A3(new_n291), .A4(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT37), .B(G110), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G12));
  NAND2_X1  g463(.A1(new_n593), .A2(new_n644), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n291), .A2(new_n347), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n624), .A2(new_n626), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n653), .A2(new_n627), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT96), .ZN(new_n655));
  OR2_X1    g469(.A1(new_n655), .A2(G900), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(G900), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n444), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n438), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n660), .A2(new_n631), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n652), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G128), .ZN(G30));
  INV_X1    g477(.A(new_n651), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n659), .B(KEYINPUT39), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(KEYINPUT99), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT99), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n664), .A2(new_n668), .A3(new_n665), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  OR2_X1    g484(.A1(new_n670), .A2(KEYINPUT40), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n343), .A2(new_n344), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(KEYINPUT38), .ZN(new_n673));
  INV_X1    g487(.A(new_n527), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n489), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n188), .B1(new_n516), .B2(new_n489), .ZN(new_n677));
  OAI21_X1  g491(.A(G472), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT97), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n591), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n432), .A2(new_n433), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n292), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n607), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n673), .A2(new_n645), .A3(new_n680), .A4(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT98), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n670), .A2(KEYINPUT40), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n671), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G143), .ZN(G45));
  NOR2_X1   g502(.A1(new_n545), .A2(new_n645), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT100), .ZN(new_n690));
  INV_X1    g504(.A(new_n659), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n607), .A2(new_n616), .A3(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n345), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n692), .ZN(new_n694));
  OAI21_X1  g508(.A(KEYINPUT100), .B1(new_n631), .B2(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n664), .A2(new_n689), .A3(new_n693), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G146), .ZN(G48));
  OAI21_X1  g511(.A(new_n188), .B1(new_n279), .B2(new_n284), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(G469), .ZN(new_n699));
  AND3_X1   g513(.A1(new_n699), .A2(new_n347), .A3(new_n285), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n589), .B1(new_n591), .B2(new_n592), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n700), .A2(new_n619), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT41), .B(G113), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G15));
  NAND4_X1  g518(.A1(new_n700), .A2(new_n633), .A3(new_n701), .A4(new_n630), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G116), .ZN(G18));
  NAND3_X1  g520(.A1(new_n593), .A2(new_n467), .A3(new_n644), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n345), .A2(new_n347), .A3(new_n285), .A4(new_n699), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(new_n301), .ZN(G21));
  OAI211_X1 g524(.A(new_n683), .B(new_n446), .C1(new_n604), .C2(new_n605), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n285), .ZN(new_n713));
  INV_X1    g527(.A(new_n250), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n281), .A2(new_n280), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n715), .B1(new_n287), .B2(new_n280), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n187), .B1(new_n716), .B2(new_n188), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n712), .A2(new_n718), .A3(new_n347), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT101), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n188), .B1(new_n501), .B2(new_n511), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n497), .B1(new_n504), .B2(new_n505), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n491), .B(new_n722), .C1(new_n498), .C2(new_n500), .ZN(new_n723));
  AOI22_X1  g537(.A1(new_n721), .A2(G472), .B1(new_n470), .B2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n585), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n720), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n723), .A2(new_n470), .ZN(new_n727));
  NOR4_X1   g541(.A1(new_n599), .A2(new_n727), .A3(KEYINPUT101), .A4(new_n585), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  OR2_X1    g543(.A1(new_n719), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G122), .ZN(G24));
  NOR3_X1   g545(.A1(new_n599), .A2(new_n645), .A3(new_n727), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n692), .ZN(new_n733));
  OAI21_X1  g547(.A(KEYINPUT102), .B1(new_n708), .B2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT102), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n724), .A2(new_n644), .A3(new_n692), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n700), .A2(new_n735), .A3(new_n736), .A4(new_n345), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G125), .ZN(G27));
  NOR2_X1   g553(.A1(new_n694), .A2(KEYINPUT42), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n347), .A2(new_n292), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n604), .A2(new_n605), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n280), .B1(new_n281), .B2(new_n714), .ZN(new_n743));
  AOI211_X1 g557(.A(new_n192), .B(new_n282), .C1(new_n275), .C2(new_n278), .ZN(new_n744));
  OAI21_X1  g558(.A(KEYINPUT103), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT103), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n288), .A2(new_n746), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n745), .A2(G469), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n285), .A2(new_n286), .ZN(new_n749));
  OAI211_X1 g563(.A(KEYINPUT104), .B(new_n742), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n745), .A2(G469), .A3(new_n747), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n285), .A3(new_n286), .ZN(new_n753));
  AOI21_X1  g567(.A(KEYINPUT104), .B1(new_n753), .B2(new_n742), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n701), .B(new_n740), .C1(new_n751), .C2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n593), .A2(new_n725), .A3(new_n692), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n742), .B1(new_n748), .B2(new_n749), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT104), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n756), .B1(new_n759), .B2(new_n750), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT42), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n755), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  XOR2_X1   g576(.A(KEYINPUT105), .B(G131), .Z(new_n763));
  XNOR2_X1  g577(.A(new_n762), .B(new_n763), .ZN(G33));
  INV_X1    g578(.A(new_n660), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n701), .B(new_n765), .C1(new_n751), .C2(new_n754), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G134), .ZN(G36));
  OR2_X1    g581(.A1(new_n607), .A2(KEYINPUT108), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n607), .A2(KEYINPUT108), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(new_n617), .A3(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT43), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n617), .A2(new_n607), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT107), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n770), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n772), .A2(KEYINPUT107), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n771), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  OAI211_X1 g592(.A(new_n778), .B(new_n644), .C1(new_n600), .C2(new_n599), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT44), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n779), .A2(new_n780), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n672), .A2(new_n293), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n781), .A2(new_n782), .A3(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n347), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n745), .A2(KEYINPUT45), .A3(new_n747), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT45), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n788), .B1(new_n743), .B2(new_n744), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT106), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(new_n790), .A3(G469), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n790), .B1(new_n789), .B2(G469), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n286), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT46), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n713), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI211_X1 g610(.A(KEYINPUT46), .B(new_n286), .C1(new_n792), .C2(new_n793), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n786), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n798), .A2(new_n665), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n785), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G137), .ZN(G39));
  NAND4_X1  g615(.A1(new_n783), .A2(new_n545), .A3(new_n589), .A4(new_n692), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(KEYINPUT109), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n798), .A2(KEYINPUT47), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT47), .ZN(new_n806));
  AOI211_X1 g620(.A(new_n806), .B(new_n786), .C1(new_n796), .C2(new_n797), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n804), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G140), .ZN(G42));
  XNOR2_X1  g623(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n738), .A2(new_n662), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT111), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  AOI22_X1  g628(.A1(new_n737), .A2(new_n734), .B1(new_n652), .B2(new_n661), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT111), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n672), .A2(new_n683), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT112), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n347), .B1(new_n691), .B2(new_n818), .ZN(new_n819));
  AOI211_X1 g633(.A(new_n819), .B(new_n644), .C1(new_n818), .C2(new_n691), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n680), .A2(new_n817), .A3(new_n753), .A4(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n696), .A2(KEYINPUT52), .A3(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n814), .A2(new_n816), .A3(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT52), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n696), .A2(new_n821), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n825), .B1(new_n812), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n604), .A2(new_n605), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n681), .A2(new_n395), .A3(new_n691), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n829), .A2(new_n292), .A3(new_n653), .A4(new_n830), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n650), .A2(new_n831), .A3(new_n651), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n759), .A2(new_n750), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n832), .B1(new_n833), .B2(new_n736), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n705), .A2(new_n702), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n607), .A2(new_n681), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n618), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n345), .A3(new_n446), .ZN(new_n838));
  OAI22_X1  g652(.A1(new_n707), .A2(new_n708), .B1(new_n602), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n835), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n647), .B1(new_n719), .B2(new_n729), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n596), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n834), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n755), .B(new_n766), .C1(new_n760), .C2(new_n761), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n811), .B1(new_n828), .B2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n815), .A2(KEYINPUT52), .A3(new_n696), .A4(new_n821), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n827), .A2(new_n847), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n845), .A2(new_n811), .A3(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n810), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT114), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n845), .A2(new_n848), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(KEYINPUT53), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n828), .A2(new_n811), .A3(new_n845), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n853), .A2(new_n854), .A3(KEYINPUT54), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT114), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n856), .B(new_n810), .C1(new_n846), .C2(new_n849), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n700), .A2(new_n783), .ZN(new_n858));
  NOR4_X1   g672(.A1(new_n858), .A2(new_n589), .A3(new_n438), .A4(new_n680), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n859), .A2(new_n608), .A3(new_n617), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n775), .A2(new_n439), .A3(new_n777), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n861), .A2(new_n729), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n860), .B(new_n435), .C1(new_n708), .C2(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n861), .A2(new_n858), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n593), .A2(new_n725), .ZN(new_n867));
  OR3_X1    g681(.A1(new_n866), .A2(KEYINPUT48), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT48), .B1(new_n866), .B2(new_n867), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n864), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n862), .A2(new_n783), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n805), .A2(new_n807), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n699), .A2(new_n285), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n347), .B1(new_n873), .B2(KEYINPUT115), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n874), .B1(KEYINPUT115), .B2(new_n873), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n871), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT50), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n673), .B1(KEYINPUT118), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n700), .A2(new_n293), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(KEYINPUT117), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n877), .A2(KEYINPUT118), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  OR2_X1    g697(.A1(new_n879), .A2(KEYINPUT117), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n881), .A2(new_n883), .A3(new_n862), .A4(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n884), .A2(new_n878), .A3(new_n880), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n882), .B1(new_n886), .B2(new_n863), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n608), .A2(new_n617), .ZN(new_n888));
  AOI22_X1  g702(.A1(new_n859), .A2(new_n888), .B1(new_n865), .B2(new_n732), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n885), .A2(new_n887), .A3(KEYINPUT51), .A4(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n870), .B1(new_n876), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n796), .A2(new_n797), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n347), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n806), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n798), .A2(KEYINPUT47), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n875), .B(KEYINPUT116), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(new_n871), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n885), .A2(new_n887), .A3(new_n889), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT51), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n891), .A2(new_n901), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n851), .A2(new_n855), .A3(new_n857), .A4(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n434), .A2(new_n190), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n585), .A2(new_n741), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(KEYINPUT110), .Z(new_n907));
  OR3_X1    g721(.A1(new_n907), .A2(new_n680), .A3(new_n770), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n873), .B(KEYINPUT49), .ZN(new_n909));
  OR3_X1    g723(.A1(new_n908), .A2(new_n673), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n905), .A2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT119), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n905), .A2(KEYINPUT119), .A3(new_n910), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(G75));
  NOR2_X1   g729(.A1(new_n190), .A2(G952), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT120), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT56), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n846), .A2(new_n849), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(G902), .ZN(new_n921));
  INV_X1    g735(.A(G210), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n919), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n321), .A2(new_n323), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(new_n329), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT55), .Z(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  OR2_X1    g741(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n923), .A2(new_n927), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n918), .B1(new_n928), .B2(new_n929), .ZN(G51));
  INV_X1    g744(.A(new_n920), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n931), .A2(new_n810), .ZN(new_n932));
  INV_X1    g746(.A(new_n850), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n286), .B(KEYINPUT57), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n716), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OR3_X1    g750(.A1(new_n921), .A2(new_n793), .A3(new_n792), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n916), .B1(new_n936), .B2(new_n937), .ZN(G54));
  INV_X1    g752(.A(new_n464), .ZN(new_n939));
  NAND2_X1  g753(.A1(KEYINPUT58), .A2(G475), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n939), .B1(new_n921), .B2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n916), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n921), .A2(new_n939), .A3(new_n940), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n943), .A2(new_n944), .ZN(G60));
  INV_X1    g759(.A(new_n614), .ZN(new_n946));
  NAND2_X1  g760(.A1(G478), .A2(G902), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT59), .Z(new_n948));
  NOR3_X1   g762(.A1(new_n934), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n851), .A2(new_n855), .A3(new_n857), .ZN(new_n950));
  INV_X1    g764(.A(new_n948), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n614), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n949), .A2(new_n918), .A3(new_n952), .ZN(G63));
  NAND2_X1  g767(.A1(G217), .A2(G902), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT60), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n920), .A2(new_n642), .A3(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n931), .A2(new_n955), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n917), .B(new_n957), .C1(new_n958), .C2(new_n580), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT61), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n959), .B(new_n960), .ZN(G66));
  AND2_X1   g775(.A1(new_n840), .A2(new_n842), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n190), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT121), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n190), .B1(new_n441), .B2(G224), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n924), .B1(G898), .B2(new_n190), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT122), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n967), .B(new_n969), .ZN(G69));
  NOR2_X1   g784(.A1(new_n450), .A2(new_n451), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT123), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n526), .B(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  OAI211_X1 g788(.A(G900), .B(G953), .C1(new_n974), .C2(G227), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n975), .B1(G227), .B2(new_n974), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n814), .A2(new_n816), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n977), .A2(new_n696), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT124), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT62), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n978), .A2(new_n979), .A3(new_n980), .A4(new_n687), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n687), .A2(new_n977), .A3(new_n696), .ZN(new_n982));
  OAI21_X1  g796(.A(KEYINPUT124), .B1(new_n982), .B2(KEYINPUT62), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n982), .A2(KEYINPUT62), .ZN(new_n985));
  INV_X1    g799(.A(new_n670), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n590), .A2(new_n595), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n986), .A2(new_n987), .A3(new_n783), .A4(new_n837), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n800), .A2(new_n808), .A3(new_n988), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n984), .A2(new_n985), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n973), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n799), .A2(new_n593), .A3(new_n725), .A4(new_n817), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(KEYINPUT125), .ZN(new_n993));
  INV_X1    g807(.A(new_n844), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n978), .A2(new_n800), .A3(new_n808), .A4(new_n994), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(G953), .B1(new_n996), .B2(new_n974), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n976), .B1(new_n991), .B2(new_n997), .ZN(G72));
  NOR3_X1   g812(.A1(new_n993), .A2(new_n995), .A3(new_n963), .ZN(new_n999));
  NAND2_X1  g813(.A1(G472), .A2(G902), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT63), .Z(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT126), .Z(new_n1002));
  OAI211_X1 g816(.A(new_n497), .B(new_n527), .C1(new_n999), .C2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n853), .A2(new_n854), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n528), .A2(new_n519), .A3(new_n531), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n1001), .ZN(new_n1006));
  OAI211_X1 g820(.A(new_n1003), .B(new_n942), .C1(new_n1004), .C2(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT127), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n984), .A2(new_n962), .A3(new_n989), .A4(new_n985), .ZN(new_n1009));
  INV_X1    g823(.A(new_n1002), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1008), .B1(new_n1011), .B2(new_n676), .ZN(new_n1012));
  AOI211_X1 g826(.A(KEYINPUT127), .B(new_n675), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1013));
  NOR3_X1   g827(.A1(new_n1007), .A2(new_n1012), .A3(new_n1013), .ZN(G57));
endmodule


