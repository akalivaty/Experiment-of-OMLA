//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 0 1 1 1 1 0 1 1 1 1 1 1 1 1 0 1 1 1 0 1 0 0 1 0 1 0 0 1 0 1 1 1 0 1 1 1 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976;
  XNOR2_X1  g000(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT93), .ZN(new_n203));
  XOR2_X1   g002(.A(G127gat), .B(G155gat), .Z(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(G15gat), .B(G22gat), .Z(new_n207));
  INV_X1    g006(.A(G1gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G15gat), .B(G22gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT16), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n210), .B1(new_n211), .B2(G1gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G8gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n213), .B(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G71gat), .A2(G78gat), .ZN(new_n216));
  INV_X1    g015(.A(G71gat), .ZN(new_n217));
  INV_X1    g016(.A(G78gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n217), .A2(new_n218), .A3(KEYINPUT9), .ZN(new_n219));
  INV_X1    g018(.A(G64gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G57gat), .ZN(new_n221));
  INV_X1    g020(.A(G57gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G64gat), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n216), .A2(new_n219), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n222), .A2(G64gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n220), .A2(G57gat), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT92), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT92), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n221), .A2(new_n223), .A3(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(KEYINPUT9), .A3(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n217), .A2(new_n218), .A3(KEYINPUT91), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT91), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(G71gat), .B2(G78gat), .ZN(new_n233));
  AOI22_X1  g032(.A1(new_n231), .A2(new_n233), .B1(G71gat), .B2(G78gat), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n224), .B1(new_n230), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT21), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n215), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT94), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n235), .A2(KEYINPUT21), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  OR2_X1    g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G183gat), .B(G211gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(G231gat), .A2(G233gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n239), .A2(new_n241), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n242), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n246), .B1(new_n242), .B2(new_n247), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n206), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n250), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n252), .A2(new_n248), .A3(new_n205), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  XOR2_X1   g053(.A(G43gat), .B(G50gat), .Z(new_n255));
  INV_X1    g054(.A(KEYINPUT15), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OR3_X1    g056(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n258));
  OAI21_X1  g057(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n259));
  AOI22_X1  g058(.A1(new_n258), .A2(new_n259), .B1(G29gat), .B2(G36gat), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT87), .ZN(new_n261));
  XNOR2_X1  g060(.A(G43gat), .B(G50gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT15), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n257), .A2(new_n260), .A3(new_n261), .A4(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n257), .A2(new_n260), .A3(new_n263), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(KEYINPUT87), .B1(new_n260), .B2(new_n263), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n264), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  AND2_X1   g068(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n270));
  NOR2_X1   g069(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n271));
  INV_X1    g070(.A(G85gat), .ZN(new_n272));
  INV_X1    g071(.A(G92gat), .ZN(new_n273));
  OAI22_X1  g072(.A1(new_n270), .A2(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT96), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT7), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AND2_X1   g076(.A1(G85gat), .A2(G92gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G99gat), .A2(G106gat), .ZN(new_n281));
  AOI22_X1  g080(.A1(KEYINPUT8), .A2(new_n281), .B1(new_n272), .B2(new_n273), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n274), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  OR2_X1    g082(.A1(G99gat), .A2(G106gat), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(new_n281), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n281), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n274), .A2(new_n280), .A3(new_n286), .A4(new_n282), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT98), .ZN(new_n290));
  XOR2_X1   g089(.A(G190gat), .B(G218gat), .Z(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(KEYINPUT97), .ZN(new_n292));
  AOI22_X1  g091(.A1(new_n269), .A2(new_n289), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n268), .A2(KEYINPUT17), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n265), .B(KEYINPUT87), .C1(new_n260), .C2(new_n263), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT17), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n295), .A2(new_n296), .A3(new_n264), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n294), .A2(new_n297), .A3(new_n288), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT41), .ZN(new_n299));
  NAND2_X1  g098(.A1(G232gat), .A2(G233gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n300), .B(KEYINPUT95), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n293), .B(new_n298), .C1(new_n299), .C2(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n292), .A2(new_n290), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n301), .A2(new_n299), .ZN(new_n305));
  XNOR2_X1  g104(.A(G134gat), .B(G162gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n305), .B(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n304), .B(new_n307), .ZN(new_n308));
  AND2_X1   g107(.A1(new_n254), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(G183gat), .A2(G190gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(G183gat), .A2(G190gat), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n310), .B1(new_n312), .B2(KEYINPUT24), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT24), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT66), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT66), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n311), .A2(new_n317), .A3(new_n314), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n313), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(G169gat), .ZN(new_n320));
  INV_X1    g119(.A(G176gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(KEYINPUT64), .B(KEYINPUT23), .ZN(new_n323));
  NOR2_X1   g122(.A1(G169gat), .A2(G176gat), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n322), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n324), .A2(KEYINPUT65), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT65), .ZN(new_n328));
  NOR3_X1   g127(.A1(new_n328), .A2(G169gat), .A3(G176gat), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT23), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n319), .A2(new_n326), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT25), .ZN(new_n332));
  INV_X1    g131(.A(G190gat), .ZN(new_n333));
  AND2_X1   g132(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n334));
  NOR2_X1   g133(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT28), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n336), .B(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT26), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n339), .B1(new_n327), .B2(new_n329), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n322), .B1(KEYINPUT26), .B2(new_n325), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n312), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n323), .A2(new_n325), .ZN(new_n344));
  INV_X1    g143(.A(new_n322), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n324), .A2(KEYINPUT23), .ZN(new_n346));
  AND3_X1   g145(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT25), .B1(new_n313), .B2(new_n315), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n332), .A2(new_n343), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(G120gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(G113gat), .ZN(new_n352));
  INV_X1    g151(.A(G113gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(G120gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT1), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(G127gat), .A2(G134gat), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(G127gat), .A2(G134gat), .ZN(new_n360));
  AOI22_X1  g159(.A1(new_n359), .A2(new_n360), .B1(KEYINPUT67), .B2(new_n356), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n360), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n363), .A2(new_n358), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n356), .B(new_n355), .C1(new_n364), .C2(KEYINPUT67), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(G227gat), .A2(G233gat), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n342), .A2(new_n338), .B1(new_n347), .B2(new_n348), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT1), .B1(new_n352), .B2(new_n354), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n361), .B(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n370), .A2(new_n372), .A3(new_n332), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n367), .A2(new_n369), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT32), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT33), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G15gat), .B(G43gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(G71gat), .B(G99gat), .ZN(new_n379));
  XOR2_X1   g178(.A(new_n378), .B(new_n379), .Z(new_n380));
  NAND3_X1  g179(.A1(new_n375), .A2(new_n377), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n380), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n374), .B(KEYINPUT32), .C1(new_n376), .C2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT69), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n369), .B1(new_n367), .B2(new_n373), .ZN(new_n386));
  XOR2_X1   g185(.A(KEYINPUT68), .B(KEYINPUT34), .Z(new_n387));
  NOR2_X1   g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT68), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT34), .ZN(new_n390));
  AOI211_X1 g189(.A(new_n369), .B(new_n390), .C1(new_n367), .C2(new_n373), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n385), .B1(new_n388), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT70), .ZN(new_n393));
  INV_X1    g192(.A(new_n390), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n386), .A2(new_n394), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n395), .B(KEYINPUT69), .C1(new_n386), .C2(new_n387), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n384), .A2(new_n392), .A3(new_n393), .A4(new_n396), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n384), .A2(new_n392), .A3(new_n396), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n395), .B1(new_n386), .B2(new_n387), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n399), .A2(new_n381), .A3(new_n383), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT70), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n397), .B1(new_n398), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT36), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT71), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n384), .B(new_n399), .ZN(new_n405));
  OR2_X1    g204(.A1(new_n405), .A2(KEYINPUT36), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT71), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n402), .A2(new_n407), .A3(KEYINPUT36), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n404), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(G228gat), .A2(G233gat), .ZN(new_n412));
  INV_X1    g211(.A(G141gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(G148gat), .ZN(new_n414));
  INV_X1    g213(.A(G148gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(G141gat), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT76), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n414), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(G155gat), .ZN(new_n419));
  INV_X1    g218(.A(G162gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(G155gat), .A2(G162gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(KEYINPUT2), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n415), .A2(KEYINPUT76), .A3(G141gat), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n418), .A2(new_n423), .A3(new_n424), .A4(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(G141gat), .B(G148gat), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n422), .B(new_n421), .C1(new_n427), .C2(KEYINPUT2), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT3), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n426), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT29), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OR2_X1    g231(.A1(G197gat), .A2(G204gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(G197gat), .A2(G204gat), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT22), .ZN(new_n435));
  NAND2_X1  g234(.A1(G211gat), .A2(G218gat), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n433), .A2(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G211gat), .B(G218gat), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(G197gat), .B(G204gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n436), .A2(new_n435), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n438), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT72), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT72), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n437), .A2(new_n445), .A3(new_n438), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n439), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT84), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n449), .B1(new_n437), .B2(new_n438), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n442), .A2(KEYINPUT84), .A3(new_n443), .ZN(new_n451));
  INV_X1    g250(.A(new_n446), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n445), .B1(new_n437), .B2(new_n438), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n450), .B(new_n451), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT3), .B1(new_n454), .B2(new_n431), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n426), .A2(new_n428), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n412), .B(new_n448), .C1(new_n455), .C2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n446), .ZN(new_n460));
  INV_X1    g259(.A(new_n439), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT73), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT73), .ZN(new_n463));
  AOI211_X1 g262(.A(new_n463), .B(new_n439), .C1(new_n444), .C2(new_n446), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n432), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n429), .B1(new_n447), .B2(KEYINPUT29), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(new_n456), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n412), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(G50gat), .B1(new_n459), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n465), .A2(new_n467), .ZN(new_n470));
  INV_X1    g269(.A(new_n412), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(G50gat), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(new_n473), .A3(new_n458), .ZN(new_n474));
  XNOR2_X1  g273(.A(G78gat), .B(G106gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n475), .B(G22gat), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  AND3_X1   g276(.A1(new_n469), .A2(new_n474), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n477), .B1(new_n469), .B2(new_n474), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n411), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR3_X1   g279(.A1(new_n459), .A2(new_n468), .A3(G50gat), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n473), .B1(new_n472), .B2(new_n458), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n476), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n469), .A2(new_n474), .A3(new_n477), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(new_n410), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n480), .A2(new_n485), .ZN(new_n486));
  OR2_X1    g285(.A1(new_n462), .A2(new_n464), .ZN(new_n487));
  NAND2_X1  g286(.A1(G226gat), .A2(G233gat), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n489), .B1(new_n350), .B2(new_n431), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n488), .B1(new_n370), .B2(new_n332), .ZN(new_n491));
  OAI211_X1 g290(.A(KEYINPUT74), .B(new_n487), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n350), .A2(new_n489), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT29), .B1(new_n370), .B2(new_n332), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n494), .B1(new_n495), .B2(new_n489), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT74), .B1(new_n496), .B2(new_n487), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n350), .A2(new_n431), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n488), .ZN(new_n500));
  INV_X1    g299(.A(new_n447), .ZN(new_n501));
  AOI211_X1 g300(.A(KEYINPUT75), .B(new_n488), .C1(new_n370), .C2(new_n332), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT75), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n503), .B1(new_n350), .B2(new_n489), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n500), .B(new_n501), .C1(new_n502), .C2(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(G8gat), .B(G36gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(G64gat), .B(G92gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n498), .A2(KEYINPUT30), .A3(new_n505), .A4(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n487), .B1(new_n490), .B2(new_n491), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT74), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n513), .A2(new_n505), .A3(new_n492), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(new_n508), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n513), .A2(new_n505), .A3(new_n492), .A4(new_n509), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT30), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n510), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(G1gat), .B(G29gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(new_n272), .ZN(new_n521));
  XNOR2_X1  g320(.A(KEYINPUT0), .B(G57gat), .ZN(new_n522));
  XOR2_X1   g321(.A(new_n521), .B(new_n522), .Z(new_n523));
  NAND2_X1  g322(.A1(G225gat), .A2(G233gat), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n456), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n525), .A2(new_n372), .A3(new_n430), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n429), .B1(new_n426), .B2(new_n428), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n527), .A2(KEYINPUT77), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT78), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  OR2_X1    g328(.A1(new_n527), .A2(KEYINPUT77), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n366), .B1(new_n527), .B2(KEYINPUT77), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT78), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n530), .A2(new_n531), .A3(new_n532), .A4(new_n430), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  NOR3_X1   g333(.A1(new_n372), .A2(KEYINPUT4), .A3(new_n456), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT80), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT4), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n537), .B1(new_n457), .B2(new_n366), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n457), .A2(new_n537), .A3(new_n366), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT80), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n536), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n524), .B1(new_n534), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT39), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n523), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n366), .B(new_n456), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(new_n524), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n538), .B1(new_n541), .B2(new_n540), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n529), .A2(new_n533), .B1(new_n549), .B2(new_n536), .ZN(new_n550));
  OAI211_X1 g349(.A(KEYINPUT39), .B(new_n548), .C1(new_n550), .C2(new_n524), .ZN(new_n551));
  AND3_X1   g350(.A1(new_n546), .A2(KEYINPUT40), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT40), .B1(new_n546), .B2(new_n551), .ZN(new_n553));
  AOI21_X1  g352(.A(KEYINPUT5), .B1(G225gat), .B2(G233gat), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n534), .A2(new_n554), .A3(new_n543), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n524), .B1(new_n535), .B2(new_n538), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n556), .B1(new_n529), .B2(new_n533), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n457), .A2(new_n366), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n372), .A2(new_n456), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n524), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT5), .ZN(new_n561));
  OAI21_X1  g360(.A(KEYINPUT79), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT79), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n563), .B(KEYINPUT5), .C1(new_n547), .C2(new_n524), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n555), .B1(new_n557), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(new_n523), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NOR3_X1   g367(.A1(new_n552), .A2(new_n553), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n486), .B1(new_n519), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n500), .B1(new_n502), .B2(new_n504), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(new_n447), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT85), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n496), .A2(new_n487), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT85), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n571), .A2(new_n575), .A3(new_n447), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n573), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT37), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT37), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n513), .A2(new_n579), .A3(new_n505), .A4(new_n492), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n580), .A2(new_n508), .ZN(new_n581));
  AOI21_X1  g380(.A(KEYINPUT38), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n514), .A2(KEYINPUT37), .ZN(new_n583));
  AND4_X1   g382(.A1(KEYINPUT38), .A2(new_n583), .A3(new_n508), .A4(new_n580), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n516), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT81), .B(KEYINPUT6), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n523), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n555), .B(new_n588), .C1(new_n557), .C2(new_n565), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n567), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n566), .A2(new_n523), .A3(new_n586), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT82), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n566), .A2(KEYINPUT82), .A3(new_n523), .A4(new_n586), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n590), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n570), .B1(new_n585), .B2(new_n595), .ZN(new_n596));
  AND3_X1   g395(.A1(new_n510), .A2(new_n515), .A3(new_n518), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(new_n486), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n409), .A2(new_n596), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(KEYINPUT86), .ZN(new_n601));
  AND2_X1   g400(.A1(new_n480), .A2(new_n485), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT86), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n595), .B(new_n597), .C1(new_n603), .C2(KEYINPUT35), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n601), .A2(new_n602), .A3(new_n604), .A4(new_n405), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n602), .A2(new_n402), .ZN(new_n606));
  OAI21_X1  g405(.A(KEYINPUT35), .B1(new_n606), .B2(new_n598), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n600), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n230), .A2(new_n234), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n287), .A2(KEYINPUT99), .ZN(new_n611));
  INV_X1    g410(.A(new_n224), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(new_n288), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT10), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n235), .A2(new_n287), .A3(new_n285), .A4(new_n611), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n289), .A2(KEYINPUT10), .A3(new_n235), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(G230gat), .ZN(new_n620));
  INV_X1    g419(.A(G233gat), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n614), .A2(new_n616), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(new_n622), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G120gat), .B(G148gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT100), .ZN(new_n629));
  XNOR2_X1  g428(.A(G176gat), .B(G204gat), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n629), .B(new_n630), .Z(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n627), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT101), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n624), .A2(new_n626), .A3(new_n631), .ZN(new_n635));
  AND3_X1   g434(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n634), .B1(new_n633), .B2(new_n635), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT89), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n639), .B1(new_n268), .B2(new_n215), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n213), .B(G8gat), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n641), .A2(KEYINPUT89), .A3(new_n295), .A4(new_n264), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(G229gat), .A2(G233gat), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n644), .B(KEYINPUT88), .Z(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n294), .A2(new_n297), .A3(new_n215), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n643), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT18), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n268), .A2(new_n215), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n643), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n645), .B(KEYINPUT13), .Z(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n643), .A2(KEYINPUT18), .A3(new_n647), .A4(new_n646), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n650), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(G113gat), .B(G141gat), .ZN(new_n658));
  INV_X1    g457(.A(G197gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(KEYINPUT11), .B(G169gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT12), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n657), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n650), .A2(new_n655), .A3(new_n656), .A4(new_n663), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n665), .A2(KEYINPUT90), .A3(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT90), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n657), .A2(new_n668), .A3(new_n664), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  AND4_X1   g470(.A1(new_n309), .A2(new_n609), .A3(new_n638), .A4(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n595), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g474(.A1(new_n672), .A2(new_n519), .ZN(new_n676));
  OAI21_X1  g475(.A(KEYINPUT42), .B1(new_n676), .B2(new_n214), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT102), .B(KEYINPUT16), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(new_n214), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  MUX2_X1   g479(.A(KEYINPUT42), .B(new_n677), .S(new_n680), .Z(G1325gat));
  AOI21_X1  g480(.A(G15gat), .B1(new_n672), .B2(new_n405), .ZN(new_n682));
  INV_X1    g481(.A(new_n409), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n672), .A2(G15gat), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n682), .B1(new_n683), .B2(new_n684), .ZN(G1326gat));
  NAND2_X1  g484(.A1(new_n672), .A2(new_n486), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT43), .B(G22gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1327gat));
  AOI21_X1  g487(.A(new_n308), .B1(new_n600), .B2(new_n608), .ZN(new_n689));
  INV_X1    g488(.A(new_n638), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n254), .A2(new_n670), .A3(new_n690), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(G29gat), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n692), .A2(new_n693), .A3(new_n673), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT45), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696));
  INV_X1    g495(.A(new_n308), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n696), .B1(new_n609), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  AOI211_X1 g498(.A(KEYINPUT44), .B(new_n308), .C1(new_n600), .C2(new_n608), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n702), .A2(new_n691), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(new_n673), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n695), .B1(new_n705), .B2(new_n693), .ZN(G1328gat));
  INV_X1    g505(.A(G36gat), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n692), .A2(new_n707), .A3(new_n519), .ZN(new_n708));
  XOR2_X1   g507(.A(new_n708), .B(KEYINPUT46), .Z(new_n709));
  NAND2_X1  g508(.A1(new_n703), .A2(new_n519), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n709), .B1(new_n711), .B2(new_n707), .ZN(G1329gat));
  OAI211_X1 g511(.A(new_n683), .B(new_n691), .C1(new_n698), .C2(new_n700), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(G43gat), .ZN(new_n714));
  INV_X1    g513(.A(G43gat), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n692), .A2(new_n715), .A3(new_n405), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n714), .A2(KEYINPUT47), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n714), .A2(KEYINPUT103), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT103), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n713), .A2(new_n719), .A3(G43gat), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n718), .A2(new_n716), .A3(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT104), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT47), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n722), .B1(new_n721), .B2(new_n723), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n717), .B1(new_n724), .B2(new_n725), .ZN(G1330gat));
  NAND3_X1  g525(.A1(new_n702), .A2(new_n486), .A3(new_n691), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(G50gat), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT105), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT48), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n692), .A2(new_n473), .A3(new_n486), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n730), .B(new_n732), .ZN(G1331gat));
  NAND2_X1  g532(.A1(new_n309), .A2(new_n670), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n734), .A2(new_n638), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n609), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n595), .B(KEYINPUT106), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(new_n222), .ZN(G1332gat));
  AOI211_X1 g538(.A(new_n597), .B(new_n736), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n740));
  NOR2_X1   g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n740), .B(new_n741), .ZN(G1333gat));
  INV_X1    g541(.A(new_n405), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n217), .B1(new_n736), .B2(new_n743), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n609), .A2(G71gat), .A3(new_n683), .A4(new_n735), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g546(.A1(new_n736), .A2(new_n602), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(new_n218), .ZN(G1335gat));
  AOI21_X1  g548(.A(new_n638), .B1(new_n699), .B2(new_n701), .ZN(new_n750));
  INV_X1    g549(.A(new_n254), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n670), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT107), .ZN(new_n753));
  AND4_X1   g552(.A1(G85gat), .A2(new_n750), .A3(new_n673), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n689), .A2(new_n753), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT51), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n689), .A2(KEYINPUT51), .A3(new_n753), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n757), .A2(KEYINPUT108), .A3(new_n758), .ZN(new_n759));
  OR2_X1    g558(.A1(new_n758), .A2(KEYINPUT108), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n759), .A2(new_n690), .A3(new_n760), .ZN(new_n761));
  OR2_X1    g560(.A1(new_n761), .A2(new_n595), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n754), .B1(new_n762), .B2(new_n272), .ZN(G1336gat));
  NAND3_X1  g562(.A1(new_n750), .A2(new_n519), .A3(new_n753), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(G92gat), .ZN(new_n765));
  XNOR2_X1  g564(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n519), .A2(new_n273), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n765), .B(new_n766), .C1(new_n761), .C2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n757), .A2(new_n758), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n597), .A2(G92gat), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n690), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT109), .ZN(new_n773));
  AOI22_X1  g572(.A1(new_n764), .A2(G92gat), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n768), .B1(new_n769), .B2(new_n774), .ZN(G1337gat));
  INV_X1    g574(.A(G99gat), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(new_n761), .B2(new_n743), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n750), .A2(G99gat), .A3(new_n683), .A4(new_n753), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(KEYINPUT111), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT111), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n777), .A2(new_n781), .A3(new_n778), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(G1338gat));
  NAND3_X1  g582(.A1(new_n750), .A2(new_n486), .A3(new_n753), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(G106gat), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n602), .A2(G106gat), .A3(new_n638), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n759), .A2(new_n760), .A3(new_n786), .ZN(new_n787));
  XNOR2_X1  g586(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n785), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n790));
  AOI22_X1  g589(.A1(new_n784), .A2(G106gat), .B1(new_n770), .B2(new_n786), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(G1339gat));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT113), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n617), .A2(new_n794), .A3(new_n622), .A4(new_n618), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n795), .A2(KEYINPUT54), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n617), .A2(new_n622), .A3(new_n618), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n622), .B1(new_n617), .B2(new_n618), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n797), .B1(new_n798), .B2(KEYINPUT113), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n631), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n800), .A2(KEYINPUT55), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT55), .B1(new_n800), .B2(new_n802), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n793), .B1(new_n805), .B2(new_n635), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n795), .A2(KEYINPUT54), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n624), .A2(new_n794), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n808), .B1(new_n809), .B2(new_n797), .ZN(new_n810));
  INV_X1    g609(.A(new_n802), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n807), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n800), .A2(KEYINPUT55), .A3(new_n802), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n812), .A2(new_n813), .A3(new_n793), .A4(new_n635), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n671), .B1(new_n806), .B2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n818), .B1(new_n652), .B2(new_n654), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n643), .A2(KEYINPUT115), .A3(new_n651), .A4(new_n653), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n646), .B1(new_n643), .B2(new_n647), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n662), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n823), .B(new_n666), .C1(new_n636), .C2(new_n637), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n816), .A2(new_n817), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n812), .A2(new_n635), .A3(new_n813), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(KEYINPUT114), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n670), .B1(new_n827), .B2(new_n814), .ZN(new_n828));
  INV_X1    g627(.A(new_n824), .ZN(new_n829));
  OAI21_X1  g628(.A(KEYINPUT116), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n825), .A2(new_n830), .A3(new_n308), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n823), .A2(new_n666), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n308), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n833), .B1(new_n806), .B2(new_n815), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n254), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n309), .A2(new_n638), .A3(new_n670), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n838), .A2(new_n486), .A3(new_n743), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n595), .A2(new_n519), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(G113gat), .B1(new_n841), .B2(new_n670), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n831), .A2(new_n834), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n751), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n836), .ZN(new_n845));
  INV_X1    g644(.A(new_n606), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n737), .A2(new_n519), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n849), .A2(new_n353), .A3(new_n671), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n842), .A2(new_n850), .ZN(G1340gat));
  OAI21_X1  g650(.A(G120gat), .B1(new_n841), .B2(new_n638), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n849), .A2(new_n351), .A3(new_n690), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(G1341gat));
  OR3_X1    g653(.A1(new_n848), .A2(KEYINPUT118), .A3(new_n751), .ZN(new_n855));
  INV_X1    g654(.A(G127gat), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT118), .B1(new_n848), .B2(new_n751), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n839), .A2(G127gat), .A3(new_n254), .A4(new_n840), .ZN(new_n859));
  OR2_X1    g658(.A1(new_n859), .A2(KEYINPUT117), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(KEYINPUT117), .ZN(new_n861));
  AND3_X1   g660(.A1(new_n858), .A2(new_n860), .A3(new_n861), .ZN(G1342gat));
  NOR3_X1   g661(.A1(new_n848), .A2(G134gat), .A3(new_n308), .ZN(new_n863));
  XNOR2_X1  g662(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n863), .B(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(G134gat), .B1(new_n841), .B2(new_n308), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(G1343gat));
  NOR3_X1   g666(.A1(new_n838), .A2(new_n519), .A3(new_n737), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n683), .A2(new_n602), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n413), .B1(new_n870), .B2(new_n670), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n409), .A2(new_n840), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n824), .B1(new_n670), .B2(new_n826), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n308), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n254), .B1(new_n874), .B2(new_n834), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n875), .A2(KEYINPUT120), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n836), .B1(new_n875), .B2(KEYINPUT120), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n486), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n872), .B1(new_n878), .B2(KEYINPUT57), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n880), .B(new_n486), .C1(new_n835), .C2(new_n837), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(G141gat), .A3(new_n671), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n871), .A2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT58), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n871), .A2(new_n883), .A3(KEYINPUT58), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(G1344gat));
  NAND3_X1  g687(.A1(new_n879), .A2(new_n690), .A3(new_n881), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT59), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n889), .A2(new_n890), .A3(G148gat), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(KEYINPUT121), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n889), .A2(new_n893), .A3(new_n890), .A4(G148gat), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n826), .ZN(new_n896));
  AOI22_X1  g695(.A1(new_n873), .A2(new_n308), .B1(new_n833), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n836), .B1(new_n897), .B2(new_n254), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT122), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT122), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n836), .B(new_n900), .C1(new_n897), .C2(new_n254), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n602), .A2(KEYINPUT57), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n899), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n486), .B1(new_n835), .B2(new_n837), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n903), .B1(new_n904), .B2(KEYINPUT57), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n905), .A2(new_n690), .A3(new_n409), .A4(new_n840), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n890), .B1(new_n906), .B2(G148gat), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n690), .A2(new_n415), .ZN(new_n908));
  OAI22_X1  g707(.A1(new_n895), .A2(new_n907), .B1(new_n870), .B2(new_n908), .ZN(G1345gat));
  INV_X1    g708(.A(KEYINPUT123), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n910), .B1(new_n870), .B2(new_n751), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n868), .A2(KEYINPUT123), .A3(new_n254), .A4(new_n869), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n911), .A2(new_n419), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n882), .A2(G155gat), .A3(new_n254), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n913), .A2(new_n914), .ZN(G1346gat));
  OAI21_X1  g714(.A(new_n420), .B1(new_n870), .B2(new_n308), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n882), .A2(G162gat), .A3(new_n697), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n916), .A2(new_n917), .ZN(G1347gat));
  NAND2_X1  g717(.A1(new_n737), .A2(new_n519), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT124), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n839), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(G169gat), .B1(new_n922), .B2(new_n670), .ZN(new_n923));
  NOR4_X1   g722(.A1(new_n838), .A2(new_n673), .A3(new_n597), .A4(new_n606), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n924), .A2(new_n320), .A3(new_n671), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(G1348gat));
  AOI21_X1  g725(.A(G176gat), .B1(new_n924), .B2(new_n690), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n922), .A2(new_n638), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n927), .B1(new_n928), .B2(G176gat), .ZN(G1349gat));
  OAI21_X1  g728(.A(G183gat), .B1(new_n922), .B2(new_n751), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n924), .B(new_n254), .C1(new_n335), .C2(new_n334), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT60), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT60), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n930), .A2(new_n934), .A3(new_n931), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n933), .A2(new_n935), .ZN(G1350gat));
  NAND3_X1  g735(.A1(new_n924), .A2(new_n333), .A3(new_n697), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n839), .A2(new_n697), .A3(new_n921), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT61), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n938), .A2(new_n939), .A3(G190gat), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n939), .B1(new_n938), .B2(G190gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n937), .B1(new_n941), .B2(new_n942), .ZN(G1351gat));
  NAND3_X1  g742(.A1(new_n845), .A2(new_n595), .A3(new_n869), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n944), .A2(new_n597), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n945), .A2(new_n659), .A3(new_n671), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT125), .ZN(new_n947));
  OR2_X1    g746(.A1(new_n905), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n920), .A2(new_n683), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n905), .A2(new_n947), .ZN(new_n950));
  AND4_X1   g749(.A1(new_n671), .A2(new_n948), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n946), .B1(new_n951), .B2(new_n659), .ZN(G1352gat));
  NAND4_X1  g751(.A1(new_n948), .A2(new_n690), .A3(new_n949), .A4(new_n950), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(G204gat), .ZN(new_n954));
  NOR4_X1   g753(.A1(new_n944), .A2(G204gat), .A3(new_n638), .A4(new_n597), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT62), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n955), .B1(KEYINPUT126), .B2(new_n956), .ZN(new_n957));
  XNOR2_X1  g756(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n958));
  OAI211_X1 g757(.A(new_n954), .B(new_n957), .C1(new_n958), .C2(new_n955), .ZN(G1353gat));
  INV_X1    g758(.A(G211gat), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n945), .A2(new_n960), .A3(new_n254), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT63), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n920), .A2(new_n751), .A3(new_n683), .ZN(new_n963));
  AOI211_X1 g762(.A(new_n962), .B(new_n960), .C1(new_n905), .C2(new_n963), .ZN(new_n964));
  INV_X1    g763(.A(new_n903), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n602), .B1(new_n844), .B2(new_n836), .ZN(new_n966));
  OAI211_X1 g765(.A(new_n965), .B(new_n963), .C1(new_n966), .C2(new_n880), .ZN(new_n967));
  AOI21_X1  g766(.A(KEYINPUT63), .B1(new_n967), .B2(G211gat), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n961), .B1(new_n964), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(KEYINPUT127), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT127), .ZN(new_n971));
  OAI211_X1 g770(.A(new_n971), .B(new_n961), .C1(new_n964), .C2(new_n968), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n970), .A2(new_n972), .ZN(G1354gat));
  INV_X1    g772(.A(G218gat), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n945), .A2(new_n974), .A3(new_n697), .ZN(new_n975));
  AND4_X1   g774(.A1(new_n697), .A2(new_n948), .A3(new_n949), .A4(new_n950), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n975), .B1(new_n976), .B2(new_n974), .ZN(G1355gat));
endmodule


