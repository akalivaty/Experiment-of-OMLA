//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 0 0 1 1 0 0 0 1 0 1 0 0 1 0 0 1 1 1 1 1 0 1 1 0 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 1 1 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n770, new_n772,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1007;
  INV_X1    g000(.A(G141gat), .ZN(new_n202));
  NAND3_X1  g001(.A1(new_n202), .A2(KEYINPUT76), .A3(G148gat), .ZN(new_n203));
  INV_X1    g002(.A(G162gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G155gat), .ZN(new_n205));
  INV_X1    g004(.A(G155gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G162gat), .ZN(new_n207));
  AND3_X1   g006(.A1(new_n203), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n202), .A2(G148gat), .ZN(new_n209));
  INV_X1    g008(.A(G148gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G141gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT76), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n209), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT2), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n204), .A2(KEYINPUT77), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT77), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G162gat), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n206), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  OAI211_X1 g017(.A(new_n208), .B(new_n213), .C1(new_n214), .C2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n205), .A2(new_n207), .ZN(new_n220));
  XNOR2_X1  g019(.A(G141gat), .B(G148gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n220), .B1(new_n221), .B2(KEYINPUT2), .ZN(new_n222));
  AND2_X1   g021(.A1(KEYINPUT69), .A2(G134gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(KEYINPUT69), .A2(G134gat), .ZN(new_n224));
  OAI21_X1  g023(.A(G127gat), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  OR2_X1    g024(.A1(G127gat), .A2(G134gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(G113gat), .B(G120gat), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n225), .B(new_n226), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  XOR2_X1   g027(.A(G113gat), .B(G120gat), .Z(new_n229));
  XOR2_X1   g028(.A(KEYINPUT70), .B(KEYINPUT1), .Z(new_n230));
  XNOR2_X1  g029(.A(G127gat), .B(G134gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n219), .A2(new_n222), .A3(new_n228), .A4(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT79), .B1(new_n233), .B2(KEYINPUT4), .ZN(new_n234));
  INV_X1    g033(.A(new_n222), .ZN(new_n235));
  XNOR2_X1  g034(.A(G155gat), .B(G162gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n213), .A2(new_n236), .A3(new_n203), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n215), .A2(new_n217), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n214), .B1(new_n239), .B2(G155gat), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n235), .B1(new_n238), .B2(new_n241), .ZN(new_n242));
  AND2_X1   g041(.A1(new_n228), .A2(new_n232), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT79), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT4), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n242), .A2(new_n243), .A3(new_n244), .A4(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n233), .A2(KEYINPUT4), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n234), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(G225gat), .A2(G233gat), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT78), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n222), .B1(new_n237), .B2(new_n240), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n243), .B1(KEYINPUT3), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT3), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n219), .A2(new_n253), .A3(new_n222), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n250), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n228), .A2(new_n232), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n256), .A2(new_n250), .A3(new_n254), .A4(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n248), .B(new_n249), .C1(new_n255), .C2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT5), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n251), .A2(new_n257), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(new_n233), .ZN(new_n263));
  INV_X1    g062(.A(new_n249), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n261), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n256), .A2(new_n257), .A3(new_n254), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT78), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n242), .A2(new_n243), .A3(new_n245), .ZN(new_n268));
  AOI22_X1  g067(.A1(new_n267), .A2(new_n258), .B1(new_n268), .B2(new_n247), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n264), .A2(KEYINPUT5), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n260), .A2(new_n265), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(G1gat), .B(G29gat), .Z(new_n272));
  XNOR2_X1  g071(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G57gat), .B(G85gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n271), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n268), .A2(new_n247), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n279), .B1(new_n255), .B2(new_n259), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT39), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n280), .A2(new_n281), .A3(new_n264), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(new_n277), .ZN(new_n283));
  OAI21_X1  g082(.A(KEYINPUT39), .B1(new_n263), .B2(new_n264), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n284), .B1(new_n280), .B2(new_n264), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT88), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n278), .B1(new_n286), .B2(KEYINPUT40), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT40), .ZN(new_n288));
  OAI211_X1 g087(.A(KEYINPUT88), .B(new_n288), .C1(new_n283), .C2(new_n285), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT22), .ZN(new_n290));
  AOI22_X1  g089(.A1(new_n290), .A2(KEYINPUT72), .B1(G211gat), .B2(G218gat), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n291), .B1(KEYINPUT72), .B2(new_n290), .ZN(new_n292));
  XNOR2_X1  g091(.A(G197gat), .B(G204gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  XOR2_X1   g093(.A(G211gat), .B(G218gat), .Z(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G169gat), .ZN(new_n298));
  INV_X1    g097(.A(G176gat), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n298), .A2(new_n299), .A3(KEYINPUT68), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT26), .ZN(new_n301));
  AOI22_X1  g100(.A1(new_n300), .A2(new_n301), .B1(G169gat), .B2(G176gat), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n298), .A2(new_n299), .A3(KEYINPUT68), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT26), .ZN(new_n304));
  AOI22_X1  g103(.A1(new_n302), .A2(new_n304), .B1(G183gat), .B2(G190gat), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT28), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n306), .A2(G190gat), .ZN(new_n307));
  AND2_X1   g106(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT67), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n307), .B(KEYINPUT67), .C1(new_n309), .C2(new_n308), .ZN(new_n313));
  AND2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AND2_X1   g113(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT27), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n309), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(G190gat), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT28), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n305), .B1(new_n314), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(G226gat), .A2(G233gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n323), .B(KEYINPUT73), .ZN(new_n324));
  NAND2_X1  g123(.A1(G183gat), .A2(G190gat), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT65), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT24), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT24), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n325), .A2(new_n326), .A3(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT66), .B(G183gat), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n328), .B(new_n330), .C1(new_n331), .C2(G190gat), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n298), .A2(new_n299), .A3(KEYINPUT23), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT23), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n334), .B1(G169gat), .B2(G176gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(G169gat), .A2(G176gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n333), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT25), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n332), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n325), .A2(KEYINPUT24), .ZN(new_n341));
  INV_X1    g140(.A(G183gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(G190gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n320), .A2(G183gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n341), .B1(new_n345), .B2(KEYINPUT24), .ZN(new_n346));
  AND3_X1   g145(.A1(new_n333), .A2(new_n335), .A3(new_n336), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT25), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT64), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n340), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n329), .A2(G183gat), .A3(G190gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(G183gat), .B(G190gat), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n351), .B1(new_n352), .B2(new_n329), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n349), .B(new_n338), .C1(new_n353), .C2(new_n337), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n322), .B(new_n324), .C1(new_n350), .C2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT29), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n324), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n338), .B1(new_n353), .B2(new_n337), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(KEYINPUT64), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n362), .A2(new_n354), .A3(new_n340), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n360), .B1(new_n363), .B2(new_n322), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n297), .B1(new_n357), .B2(new_n364), .ZN(new_n365));
  AOI22_X1  g164(.A1(new_n361), .A2(KEYINPUT64), .B1(new_n332), .B2(new_n339), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n309), .B1(new_n331), .B2(KEYINPUT27), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n306), .B1(new_n367), .B2(G190gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n312), .A2(new_n313), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI22_X1  g169(.A1(new_n366), .A2(new_n354), .B1(new_n370), .B2(new_n305), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n356), .B(new_n296), .C1(new_n371), .C2(new_n360), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n365), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G8gat), .B(G36gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(G64gat), .B(G92gat), .ZN(new_n375));
  XOR2_X1   g174(.A(new_n374), .B(new_n375), .Z(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n365), .A2(KEYINPUT74), .A3(new_n372), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT74), .B1(new_n365), .B2(new_n372), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n377), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n378), .B1(new_n382), .B2(KEYINPUT30), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n365), .A2(KEYINPUT30), .A3(new_n372), .A4(new_n376), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT75), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n384), .B(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n287), .B(new_n289), .C1(new_n383), .C2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT37), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT74), .ZN(new_n390));
  INV_X1    g189(.A(new_n372), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n322), .B1(new_n350), .B2(new_n355), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n359), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n296), .B1(new_n393), .B2(new_n356), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n390), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n389), .B1(new_n395), .B2(new_n379), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n377), .B1(new_n373), .B2(KEYINPUT37), .ZN(new_n397));
  OAI21_X1  g196(.A(KEYINPUT38), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n397), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT38), .B1(new_n373), .B2(KEYINPUT37), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n378), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  XOR2_X1   g200(.A(KEYINPUT82), .B(KEYINPUT6), .Z(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n260), .A2(new_n265), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n269), .A2(new_n270), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(new_n277), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT81), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n404), .A2(new_n405), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n276), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n403), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n404), .A2(KEYINPUT81), .A3(new_n277), .A4(new_n405), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n278), .B1(new_n412), .B2(new_n402), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n398), .B(new_n401), .C1(new_n411), .C2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT87), .B(G22gat), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  XOR2_X1   g215(.A(G78gat), .B(G106gat), .Z(new_n417));
  XNOR2_X1  g216(.A(new_n417), .B(KEYINPUT84), .ZN(new_n418));
  INV_X1    g217(.A(G50gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n418), .B(new_n419), .ZN(new_n420));
  XOR2_X1   g219(.A(KEYINPUT83), .B(KEYINPUT31), .Z(new_n421));
  XNOR2_X1  g220(.A(new_n420), .B(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n296), .B1(new_n358), .B2(new_n254), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n294), .A2(new_n295), .ZN(new_n425));
  INV_X1    g224(.A(new_n295), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n426), .B1(new_n292), .B2(new_n293), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n358), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n242), .B1(new_n428), .B2(new_n253), .ZN(new_n429));
  NAND2_X1  g228(.A1(G228gat), .A2(G233gat), .ZN(new_n430));
  OR3_X1    g229(.A1(new_n424), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  XOR2_X1   g230(.A(new_n430), .B(KEYINPUT85), .Z(new_n432));
  OAI211_X1 g231(.A(KEYINPUT86), .B(new_n432), .C1(new_n424), .C2(new_n429), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n432), .B1(new_n424), .B2(new_n429), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT86), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n423), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n431), .A2(new_n433), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n435), .A2(new_n436), .ZN(new_n440));
  NOR3_X1   g239(.A1(new_n439), .A2(new_n440), .A3(new_n422), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n416), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n434), .A2(new_n423), .A3(new_n437), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n422), .B1(new_n439), .B2(new_n440), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(new_n415), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n388), .A2(new_n414), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT36), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT33), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n257), .B(new_n322), .C1(new_n350), .C2(new_n355), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n257), .B1(new_n363), .B2(new_n322), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(G227gat), .ZN(new_n454));
  INV_X1    g253(.A(G233gat), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT71), .B1(new_n453), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n392), .A2(new_n243), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n458), .A2(KEYINPUT71), .A3(new_n456), .A4(new_n450), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n449), .B1(new_n457), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT34), .B1(new_n453), .B2(new_n456), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n458), .A2(new_n450), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT34), .ZN(new_n464));
  INV_X1    g263(.A(new_n456), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  XOR2_X1   g266(.A(G15gat), .B(G43gat), .Z(new_n468));
  XNOR2_X1  g267(.A(G71gat), .B(G99gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n468), .B(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n461), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n458), .A2(new_n456), .A3(new_n450), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT71), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(new_n459), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT32), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n464), .B1(new_n463), .B2(new_n465), .ZN(new_n478));
  AOI211_X1 g277(.A(KEYINPUT34), .B(new_n456), .C1(new_n458), .C2(new_n450), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT33), .B1(new_n474), .B2(new_n459), .ZN(new_n481));
  INV_X1    g280(.A(new_n470), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n471), .A2(new_n477), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n477), .B1(new_n471), .B2(new_n483), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n448), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NOR3_X1   g285(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n467), .B1(new_n461), .B2(new_n470), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n476), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n471), .A2(new_n477), .A3(new_n483), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n489), .A2(KEYINPUT36), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n446), .ZN(new_n492));
  INV_X1    g291(.A(new_n378), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n376), .B1(new_n395), .B2(new_n379), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT30), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT81), .B1(new_n271), .B2(new_n277), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n402), .B1(new_n497), .B2(new_n278), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n412), .A2(new_n402), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n410), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n496), .A2(new_n498), .A3(new_n500), .A4(new_n386), .ZN(new_n501));
  AOI22_X1  g300(.A1(new_n486), .A2(new_n491), .B1(new_n492), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n489), .A2(new_n446), .A3(new_n490), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT35), .B1(new_n503), .B2(new_n501), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n484), .A2(new_n485), .ZN(new_n505));
  AND4_X1   g304(.A1(new_n500), .A2(new_n496), .A3(new_n498), .A4(new_n386), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT35), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n505), .A2(new_n506), .A3(new_n507), .A4(new_n446), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n447), .A2(new_n502), .B1(new_n504), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT15), .ZN(new_n510));
  XNOR2_X1  g309(.A(G43gat), .B(G50gat), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT91), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(G43gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(new_n419), .ZN(new_n515));
  NAND2_X1  g314(.A1(G43gat), .A2(G50gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(KEYINPUT91), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n511), .A2(KEYINPUT15), .ZN(new_n519));
  INV_X1    g318(.A(G29gat), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n520), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT14), .B(G29gat), .ZN(new_n523));
  INV_X1    g322(.A(G36gat), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n518), .B1(new_n519), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT17), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n523), .A2(new_n524), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n517), .B(new_n513), .C1(new_n528), .C2(new_n522), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n526), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G15gat), .B(G22gat), .ZN(new_n531));
  INV_X1    g330(.A(G1gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(KEYINPUT16), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n534), .B1(G1gat), .B2(new_n531), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(G8gat), .ZN(new_n536));
  INV_X1    g335(.A(G8gat), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n534), .B(new_n537), .C1(G1gat), .C2(new_n531), .ZN(new_n538));
  AND2_X1   g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n530), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n526), .A2(new_n529), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT92), .B1(new_n541), .B2(KEYINPUT17), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT92), .ZN(new_n543));
  AOI211_X1 g342(.A(new_n543), .B(new_n527), .C1(new_n526), .C2(new_n529), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n540), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(G229gat), .A2(G233gat), .ZN(new_n546));
  XOR2_X1   g345(.A(new_n546), .B(KEYINPUT93), .Z(new_n547));
  INV_X1    g346(.A(new_n539), .ZN(new_n548));
  INV_X1    g347(.A(new_n541), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n545), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT18), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n545), .A2(KEYINPUT18), .A3(new_n547), .A4(new_n550), .ZN(new_n554));
  OR3_X1    g353(.A1(new_n548), .A2(new_n549), .A3(KEYINPUT94), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n541), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n550), .A2(KEYINPUT94), .A3(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n547), .B(KEYINPUT13), .Z(new_n558));
  NAND3_X1  g357(.A1(new_n555), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n553), .A2(new_n554), .A3(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(KEYINPUT89), .B(KEYINPUT11), .Z(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT90), .ZN(new_n562));
  XOR2_X1   g361(.A(G113gat), .B(G141gat), .Z(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  XOR2_X1   g363(.A(G169gat), .B(G197gat), .Z(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n566), .B(KEYINPUT12), .Z(new_n567));
  NAND2_X1  g366(.A1(new_n560), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n566), .B(KEYINPUT12), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n569), .A2(new_n553), .A3(new_n554), .A4(new_n559), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n509), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n574));
  NAND2_X1  g373(.A1(G231gat), .A2(G233gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G183gat), .B(G211gat), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n576), .B(new_n577), .Z(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G127gat), .B(G155gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(G57gat), .B(G64gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT95), .ZN(new_n582));
  NAND2_X1  g381(.A1(G71gat), .A2(G78gat), .ZN(new_n583));
  OR2_X1    g382(.A1(G71gat), .A2(G78gat), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT9), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(G64gat), .ZN(new_n587));
  OR3_X1    g386(.A1(new_n587), .A2(KEYINPUT95), .A3(G57gat), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n582), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n583), .B(new_n584), .C1(new_n581), .C2(new_n585), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT96), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n589), .A2(KEYINPUT96), .A3(new_n590), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n580), .B1(new_n595), .B2(KEYINPUT21), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n548), .B1(new_n595), .B2(KEYINPUT21), .ZN(new_n598));
  NOR3_X1   g397(.A1(new_n595), .A2(KEYINPUT21), .A3(new_n580), .ZN(new_n599));
  NOR3_X1   g398(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n595), .A2(KEYINPUT21), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(new_n539), .ZN(new_n602));
  INV_X1    g401(.A(new_n599), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n602), .B1(new_n603), .B2(new_n596), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n579), .B1(new_n600), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n598), .B1(new_n597), .B2(new_n599), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n603), .A2(new_n602), .A3(new_n596), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n606), .A2(new_n607), .A3(new_n578), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(G99gat), .A2(G106gat), .ZN(new_n610));
  OR2_X1    g409(.A1(G99gat), .A2(G106gat), .ZN(new_n611));
  NAND2_X1  g410(.A1(G85gat), .A2(G92gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(G85gat), .ZN(new_n615));
  INV_X1    g414(.A(G92gat), .ZN(new_n616));
  AOI22_X1  g415(.A1(KEYINPUT8), .A2(new_n610), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  OAI211_X1 g417(.A(new_n610), .B(new_n611), .C1(new_n614), .C2(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n612), .B(new_n613), .Z(new_n620));
  NAND2_X1  g419(.A1(new_n611), .A2(new_n610), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n620), .A2(new_n621), .A3(new_n617), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n530), .B(new_n623), .C1(new_n542), .C2(new_n544), .ZN(new_n624));
  XOR2_X1   g423(.A(G190gat), .B(G218gat), .Z(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G232gat), .A2(G233gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT97), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT41), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n619), .A2(new_n622), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n630), .B1(new_n549), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n624), .A2(new_n626), .A3(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n626), .B1(new_n624), .B2(new_n632), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n628), .A2(new_n629), .ZN(new_n636));
  XNOR2_X1  g435(.A(G134gat), .B(G162gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  OAI22_X1  g438(.A1(new_n634), .A2(new_n635), .B1(KEYINPUT99), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n635), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n638), .B(KEYINPUT99), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n641), .A2(new_n633), .A3(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n609), .A2(new_n640), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(KEYINPUT100), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT100), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n609), .A2(new_n640), .A3(new_n644), .A4(new_n647), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(G230gat), .A2(G233gat), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n651), .B(KEYINPUT101), .Z(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n594), .ZN(new_n654));
  AOI21_X1  g453(.A(KEYINPUT96), .B1(new_n589), .B2(new_n590), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n623), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n631), .A2(new_n591), .ZN(new_n657));
  AOI21_X1  g456(.A(KEYINPUT10), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT10), .ZN(new_n659));
  AOI211_X1 g458(.A(new_n659), .B(new_n623), .C1(new_n593), .C2(new_n594), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n653), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  AND3_X1   g460(.A1(new_n591), .A2(new_n622), .A3(new_n619), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n662), .B1(new_n595), .B2(new_n623), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(new_n652), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(G120gat), .B(G148gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(G176gat), .B(G204gat), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n666), .B(new_n667), .Z(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n661), .A2(new_n664), .A3(new_n668), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n650), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n573), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n498), .A2(new_n500), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(new_n532), .ZN(G1324gat));
  NAND2_X1  g477(.A1(new_n496), .A2(new_n386), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT102), .B(KEYINPUT16), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(G8gat), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n684), .B1(new_n537), .B2(new_n681), .ZN(new_n685));
  MUX2_X1   g484(.A(new_n684), .B(new_n685), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g485(.A1(new_n486), .A2(new_n491), .ZN(new_n687));
  OAI21_X1  g486(.A(G15gat), .B1(new_n674), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n505), .ZN(new_n689));
  OR2_X1    g488(.A1(new_n689), .A2(G15gat), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n688), .B1(new_n674), .B2(new_n690), .ZN(G1326gat));
  NOR2_X1   g490(.A1(new_n674), .A2(new_n446), .ZN(new_n692));
  XOR2_X1   g491(.A(KEYINPUT43), .B(G22gat), .Z(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1327gat));
  NOR2_X1   g493(.A1(new_n609), .A2(new_n672), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n640), .A2(new_n644), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n573), .A2(new_n699), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n700), .A2(G29gat), .A3(new_n676), .ZN(new_n701));
  XNOR2_X1  g500(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(new_n703));
  OR2_X1    g502(.A1(new_n697), .A2(KEYINPUT105), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n697), .A2(KEYINPUT105), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n509), .A2(KEYINPUT44), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n504), .A2(new_n508), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n492), .A2(new_n501), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n687), .A2(new_n710), .A3(new_n447), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n698), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n713));
  OAI21_X1  g512(.A(KEYINPUT104), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT104), .ZN(new_n715));
  OAI211_X1 g514(.A(new_n715), .B(KEYINPUT44), .C1(new_n509), .C2(new_n698), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n708), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n572), .A2(new_n696), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n717), .A2(new_n676), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n703), .B1(new_n520), .B2(new_n720), .ZN(G1328gat));
  NAND2_X1  g520(.A1(new_n714), .A2(new_n716), .ZN(new_n722));
  INV_X1    g521(.A(new_n708), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n719), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n524), .B1(new_n724), .B2(new_n679), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n573), .A2(new_n524), .A3(new_n679), .A4(new_n699), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT46), .ZN(new_n727));
  OAI21_X1  g526(.A(KEYINPUT106), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT46), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n726), .B(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT106), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n717), .A2(new_n680), .A3(new_n719), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n730), .B(new_n731), .C1(new_n732), .C2(new_n524), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n728), .A2(new_n733), .ZN(G1329gat));
  NOR2_X1   g533(.A1(new_n687), .A2(new_n514), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n724), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n700), .A2(new_n689), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n737), .A2(G43gat), .ZN(new_n738));
  OAI21_X1  g537(.A(KEYINPUT47), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n735), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT47), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n740), .B(new_n741), .C1(G43gat), .C2(new_n737), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n739), .A2(new_n742), .ZN(G1330gat));
  NOR3_X1   g542(.A1(new_n700), .A2(G50gat), .A3(new_n446), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT48), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n419), .B1(new_n724), .B2(new_n492), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n747), .B1(new_n748), .B2(new_n744), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n717), .A2(new_n446), .A3(new_n719), .ZN(new_n750));
  OAI221_X1 g549(.A(new_n745), .B1(new_n746), .B2(KEYINPUT48), .C1(new_n750), .C2(new_n419), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(G1331gat));
  INV_X1    g551(.A(new_n672), .ZN(new_n753));
  NOR4_X1   g552(.A1(new_n509), .A2(new_n571), .A3(new_n650), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n675), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(G57gat), .ZN(G1332gat));
  OR2_X1    g555(.A1(new_n679), .A2(KEYINPUT108), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n679), .A2(KEYINPUT108), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n760), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n754), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g561(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n762), .B(new_n763), .ZN(new_n764));
  XNOR2_X1  g563(.A(KEYINPUT109), .B(KEYINPUT110), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n764), .B(new_n765), .ZN(G1333gat));
  INV_X1    g565(.A(new_n687), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n754), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n689), .A2(G71gat), .ZN(new_n769));
  AOI22_X1  g568(.A1(new_n768), .A2(G71gat), .B1(new_n754), .B2(new_n769), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g570(.A1(new_n754), .A2(new_n492), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g572(.A1(new_n675), .A2(new_n615), .A3(new_n672), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT114), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT51), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n709), .A2(new_n711), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT112), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n777), .A2(new_n778), .A3(new_n697), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n571), .A2(new_n609), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n712), .A2(new_n778), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n776), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n780), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n784), .B1(new_n712), .B2(new_n778), .ZN(new_n785));
  OAI21_X1  g584(.A(KEYINPUT112), .B1(new_n509), .B2(new_n698), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n785), .A2(KEYINPUT51), .A3(new_n786), .ZN(new_n787));
  AND3_X1   g586(.A1(new_n783), .A2(KEYINPUT113), .A3(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(KEYINPUT113), .B1(new_n783), .B2(new_n787), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n775), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n784), .A2(new_n753), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n717), .A2(new_n676), .A3(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT111), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(G85gat), .B1(new_n793), .B2(new_n794), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n790), .B1(new_n795), .B2(new_n796), .ZN(G1336gat));
  INV_X1    g596(.A(KEYINPUT115), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n760), .A2(G92gat), .A3(new_n753), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  AOI211_X1 g599(.A(new_n798), .B(new_n800), .C1(new_n783), .C2(new_n787), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n792), .B1(new_n722), .B2(new_n723), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n616), .B1(new_n802), .B2(new_n679), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT52), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n787), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT51), .B1(new_n785), .B2(new_n786), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n799), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(KEYINPUT115), .A2(KEYINPUT52), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n717), .A2(new_n760), .A3(new_n792), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n616), .A2(KEYINPUT52), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n807), .B(new_n808), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n804), .A2(new_n811), .ZN(G1337gat));
  NOR3_X1   g611(.A1(new_n689), .A2(G99gat), .A3(new_n753), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n813), .B1(new_n788), .B2(new_n789), .ZN(new_n814));
  INV_X1    g613(.A(new_n802), .ZN(new_n815));
  OAI21_X1  g614(.A(G99gat), .B1(new_n815), .B2(new_n687), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(G1338gat));
  INV_X1    g616(.A(G106gat), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n818), .B1(new_n802), .B2(new_n492), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n753), .A2(G106gat), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n492), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n821), .B1(new_n783), .B2(new_n787), .ZN(new_n822));
  OAI21_X1  g621(.A(KEYINPUT53), .B1(new_n819), .B2(new_n822), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n492), .B(new_n820), .C1(new_n805), .C2(new_n806), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n717), .A2(new_n446), .A3(new_n792), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n824), .B(new_n825), .C1(new_n818), .C2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n823), .A2(new_n827), .ZN(G1339gat));
  NAND4_X1  g627(.A1(new_n572), .A2(new_n646), .A3(new_n648), .A4(new_n753), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n558), .B1(new_n555), .B2(new_n557), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n547), .B1(new_n545), .B2(new_n550), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n566), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n570), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n656), .A2(new_n657), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n659), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n595), .A2(new_n631), .A3(KEYINPUT10), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n652), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n668), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n652), .B(new_n837), .C1(new_n663), .C2(KEYINPUT10), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n661), .A2(new_n841), .A3(KEYINPUT54), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n840), .A2(KEYINPUT55), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n671), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n845));
  INV_X1    g644(.A(new_n842), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n669), .B1(new_n661), .B2(KEYINPUT54), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(KEYINPUT116), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n840), .A2(new_n842), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n850), .A2(new_n851), .A3(new_n845), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n844), .B1(new_n849), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n706), .A2(new_n834), .A3(new_n853), .ZN(new_n854));
  AND3_X1   g653(.A1(new_n570), .A2(new_n672), .A3(new_n833), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n855), .B1(new_n853), .B2(new_n571), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n707), .B1(new_n856), .B2(KEYINPUT117), .ZN(new_n857));
  INV_X1    g656(.A(new_n671), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n846), .A2(new_n847), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n858), .B1(new_n859), .B2(KEYINPUT55), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n851), .B1(new_n850), .B2(new_n845), .ZN(new_n861));
  AOI211_X1 g660(.A(KEYINPUT116), .B(KEYINPUT55), .C1(new_n840), .C2(new_n842), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n571), .B(new_n860), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n855), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT117), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n854), .B1(new_n857), .B2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n609), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n830), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n870), .A2(new_n492), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n871), .A2(new_n675), .A3(new_n505), .A4(new_n760), .ZN(new_n872));
  OAI21_X1  g671(.A(G113gat), .B1(new_n872), .B2(new_n572), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n706), .A2(new_n834), .A3(new_n853), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n706), .B1(new_n865), .B2(new_n866), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n856), .A2(KEYINPUT117), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n829), .B1(new_n877), .B2(new_n609), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n675), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n879), .A2(new_n503), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n760), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n572), .A2(G113gat), .ZN(new_n882));
  XOR2_X1   g681(.A(new_n882), .B(KEYINPUT118), .Z(new_n883));
  OAI21_X1  g682(.A(new_n873), .B1(new_n881), .B2(new_n883), .ZN(G1340gat));
  INV_X1    g683(.A(G120gat), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n872), .A2(new_n885), .A3(new_n753), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n880), .A2(new_n672), .A3(new_n760), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n886), .B1(new_n887), .B2(new_n885), .ZN(G1341gat));
  OAI21_X1  g687(.A(G127gat), .B1(new_n872), .B2(new_n869), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n869), .A2(G127gat), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n889), .B1(new_n881), .B2(new_n890), .ZN(G1342gat));
  NAND2_X1  g690(.A1(new_n680), .A2(new_n697), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT119), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n893), .A2(new_n224), .A3(new_n223), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n880), .A2(new_n894), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n895), .A2(KEYINPUT56), .ZN(new_n896));
  OAI21_X1  g695(.A(G134gat), .B1(new_n872), .B2(new_n698), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n895), .A2(KEYINPUT56), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(G1343gat));
  NOR3_X1   g698(.A1(new_n767), .A2(new_n676), .A3(new_n759), .ZN(new_n900));
  AOI21_X1  g699(.A(KEYINPUT57), .B1(new_n878), .B2(new_n492), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT57), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n446), .A2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  AND3_X1   g703(.A1(new_n571), .A2(new_n860), .A3(new_n848), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n698), .B1(new_n905), .B2(new_n855), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n854), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n869), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n904), .B1(new_n908), .B2(new_n829), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n571), .B(new_n900), .C1(new_n901), .C2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(G141gat), .ZN(new_n911));
  AND2_X1   g710(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n687), .A2(new_n492), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n879), .A2(new_n759), .A3(new_n913), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n572), .A2(G141gat), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n912), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g715(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n911), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(new_n911), .B2(new_n916), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n919), .A2(new_n920), .ZN(G1344gat));
  INV_X1    g720(.A(KEYINPUT59), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n900), .B1(new_n901), .B2(new_n909), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n922), .B(G148gat), .C1(new_n923), .C2(new_n753), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n853), .A2(new_n697), .A3(new_n834), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n609), .B1(new_n906), .B2(new_n925), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n649), .A2(KEYINPUT121), .A3(new_n572), .A4(new_n753), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT121), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n829), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n492), .B1(new_n926), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(new_n902), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n932), .B1(new_n870), .B2(new_n904), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n900), .A2(new_n672), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n210), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT122), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n936), .A2(new_n937), .A3(new_n922), .ZN(new_n938));
  AOI22_X1  g737(.A1(new_n878), .A2(new_n903), .B1(new_n902), .B2(new_n931), .ZN(new_n939));
  OAI21_X1  g738(.A(G148gat), .B1(new_n939), .B2(new_n934), .ZN(new_n940));
  AOI21_X1  g739(.A(KEYINPUT122), .B1(new_n940), .B2(KEYINPUT59), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n924), .B1(new_n938), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n914), .A2(new_n210), .A3(new_n672), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1345gat));
  OAI21_X1  g743(.A(G155gat), .B1(new_n923), .B2(new_n869), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n914), .A2(new_n206), .A3(new_n609), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1346gat));
  OAI21_X1  g746(.A(new_n239), .B1(new_n923), .B2(new_n707), .ZN(new_n948));
  OR4_X1    g747(.A1(new_n239), .A2(new_n879), .A3(new_n893), .A4(new_n913), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(G1347gat));
  NOR2_X1   g749(.A1(new_n680), .A2(new_n675), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n951), .A2(new_n505), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n871), .A2(new_n952), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n953), .A2(new_n298), .A3(new_n572), .ZN(new_n954));
  OAI21_X1  g753(.A(KEYINPUT123), .B1(new_n870), .B2(new_n675), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT123), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n878), .A2(new_n956), .A3(new_n676), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n760), .A2(new_n503), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n958), .A2(new_n571), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n954), .B1(new_n960), .B2(new_n298), .ZN(G1348gat));
  OAI21_X1  g760(.A(G176gat), .B1(new_n953), .B2(new_n753), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n958), .A2(new_n959), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n672), .A2(new_n299), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(G1349gat));
  INV_X1    g764(.A(new_n308), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n869), .B1(new_n318), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n958), .A2(new_n959), .A3(new_n967), .ZN(new_n968));
  OR2_X1    g767(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n878), .A2(new_n446), .A3(new_n609), .A4(new_n952), .ZN(new_n970));
  AOI22_X1  g769(.A1(new_n970), .A2(new_n331), .B1(KEYINPUT124), .B2(KEYINPUT60), .ZN(new_n971));
  AND3_X1   g770(.A1(new_n968), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n969), .B1(new_n968), .B2(new_n971), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n972), .A2(new_n973), .ZN(G1350gat));
  OAI21_X1  g773(.A(G190gat), .B1(new_n953), .B2(new_n698), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n975), .A2(KEYINPUT61), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n975), .A2(KEYINPUT61), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n706), .A2(new_n320), .ZN(new_n978));
  OAI22_X1  g777(.A1(new_n976), .A2(new_n977), .B1(new_n963), .B2(new_n978), .ZN(G1351gat));
  AND2_X1   g778(.A1(new_n687), .A2(new_n951), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n933), .A2(new_n980), .ZN(new_n981));
  INV_X1    g780(.A(G197gat), .ZN(new_n982));
  NOR3_X1   g781(.A1(new_n981), .A2(new_n982), .A3(new_n572), .ZN(new_n983));
  AOI211_X1 g782(.A(new_n760), .B(new_n913), .C1(new_n955), .C2(new_n957), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n984), .A2(new_n571), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n983), .B1(new_n985), .B2(new_n982), .ZN(G1352gat));
  AND2_X1   g785(.A1(new_n933), .A2(new_n980), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT126), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n987), .A2(new_n988), .A3(new_n672), .ZN(new_n989));
  OAI21_X1  g788(.A(KEYINPUT126), .B1(new_n981), .B2(new_n753), .ZN(new_n990));
  XNOR2_X1  g789(.A(KEYINPUT125), .B(G204gat), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n753), .A2(new_n991), .ZN(new_n993));
  AND3_X1   g792(.A1(new_n984), .A2(KEYINPUT62), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g793(.A(KEYINPUT62), .B1(new_n984), .B2(new_n993), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n992), .B1(new_n994), .B2(new_n995), .ZN(G1353gat));
  NAND3_X1  g795(.A1(new_n933), .A2(new_n609), .A3(new_n980), .ZN(new_n997));
  AND3_X1   g796(.A1(new_n997), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n998));
  AOI21_X1  g797(.A(KEYINPUT63), .B1(new_n997), .B2(G211gat), .ZN(new_n999));
  NOR2_X1   g798(.A1(new_n913), .A2(new_n760), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n958), .A2(new_n1000), .ZN(new_n1001));
  OR2_X1    g800(.A1(new_n869), .A2(G211gat), .ZN(new_n1002));
  OAI22_X1  g801(.A1(new_n998), .A2(new_n999), .B1(new_n1001), .B2(new_n1002), .ZN(G1354gat));
  OAI21_X1  g802(.A(new_n697), .B1(new_n987), .B2(KEYINPUT127), .ZN(new_n1004));
  AND3_X1   g803(.A1(new_n933), .A2(KEYINPUT127), .A3(new_n980), .ZN(new_n1005));
  OAI21_X1  g804(.A(G218gat), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  OR3_X1    g805(.A1(new_n1001), .A2(G218gat), .A3(new_n707), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1006), .A2(new_n1007), .ZN(G1355gat));
endmodule


