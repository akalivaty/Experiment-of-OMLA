//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 1 1 1 1 0 1 0 0 1 1 1 0 0 0 1 0 0 0 1 0 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 0 0 0 0 1 0 1 0 0 1 0 0 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n538, new_n539, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n600, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187, new_n1188, new_n1189;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT64), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI211_X1 g040(.A(G137), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G101), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n463), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g044(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n463), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n469), .A2(new_n472), .ZN(G160));
  INV_X1    g048(.A(new_n464), .ZN(new_n474));
  INV_X1    g049(.A(new_n465), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n463), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n463), .A2(G112), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G136), .ZN(new_n480));
  XNOR2_X1  g055(.A(KEYINPUT3), .B(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(new_n463), .ZN(new_n482));
  OAI221_X1 g057(.A(new_n477), .B1(new_n478), .B2(new_n479), .C1(new_n480), .C2(new_n482), .ZN(new_n483));
  XOR2_X1   g058(.A(new_n483), .B(KEYINPUT66), .Z(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  OAI211_X1 g060(.A(G126), .B(G2105), .C1(new_n464), .C2(new_n465), .ZN(new_n486));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n487), .A2(new_n489), .A3(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n493), .B1(new_n464), .B2(new_n465), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n493), .B(new_n496), .C1(new_n465), .C2(new_n464), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n491), .B1(new_n495), .B2(new_n497), .ZN(G164));
  OR2_X1    g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n501), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT6), .B(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G88), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G50), .ZN(new_n509));
  OAI22_X1  g084(.A1(new_n506), .A2(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n504), .A2(new_n510), .ZN(G166));
  NAND3_X1  g086(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n512));
  XNOR2_X1  g087(.A(new_n512), .B(KEYINPUT7), .ZN(new_n513));
  INV_X1    g088(.A(G51), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n513), .B1(new_n508), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n500), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n505), .A2(G89), .ZN(new_n519));
  NAND2_X1  g094(.A1(G63), .A2(G651), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n515), .A2(new_n521), .ZN(G168));
  AOI22_X1  g097(.A1(new_n501), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n523), .A2(new_n503), .ZN(new_n524));
  INV_X1    g099(.A(G90), .ZN(new_n525));
  INV_X1    g100(.A(G52), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n506), .A2(new_n525), .B1(new_n508), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n524), .A2(new_n527), .ZN(G171));
  AOI22_X1  g103(.A1(new_n501), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(new_n503), .ZN(new_n530));
  XOR2_X1   g105(.A(KEYINPUT67), .B(G81), .Z(new_n531));
  INV_X1    g106(.A(G43), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n506), .A2(new_n531), .B1(new_n508), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G860), .ZN(new_n535));
  XOR2_X1   g110(.A(new_n535), .B(KEYINPUT68), .Z(G153));
  NAND4_X1  g111(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g112(.A1(G1), .A2(G3), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT8), .ZN(new_n539));
  NAND4_X1  g114(.A1(G319), .A2(G483), .A3(G661), .A4(new_n539), .ZN(G188));
  AND2_X1   g115(.A1(KEYINPUT6), .A2(G651), .ZN(new_n541));
  NOR2_X1   g116(.A1(KEYINPUT6), .A2(G651), .ZN(new_n542));
  OAI211_X1 g117(.A(G53), .B(G543), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT69), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n543), .A2(new_n544), .A3(KEYINPUT9), .ZN(new_n545));
  INV_X1    g120(.A(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(KEYINPUT6), .A2(G651), .ZN(new_n547));
  NAND2_X1  g122(.A1(KEYINPUT6), .A2(G651), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n544), .A2(KEYINPUT9), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n549), .A2(G53), .A3(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n499), .A2(new_n500), .B1(new_n547), .B2(new_n548), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n545), .A2(new_n551), .B1(new_n552), .B2(G91), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT70), .ZN(new_n554));
  INV_X1    g129(.A(G65), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n555), .B1(new_n499), .B2(new_n500), .ZN(new_n556));
  NAND2_X1  g131(.A1(G78), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n554), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  OAI211_X1 g134(.A(KEYINPUT70), .B(new_n557), .C1(new_n518), .C2(new_n555), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n559), .A2(new_n560), .A3(G651), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n553), .A2(new_n561), .ZN(G299));
  INV_X1    g137(.A(G171), .ZN(G301));
  INV_X1    g138(.A(G168), .ZN(G286));
  INV_X1    g139(.A(G166), .ZN(G303));
  NAND2_X1  g140(.A1(new_n552), .A2(G87), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n501), .B2(G74), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n549), .A2(G49), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(G288));
  INV_X1    g144(.A(G86), .ZN(new_n570));
  INV_X1    g145(.A(G48), .ZN(new_n571));
  OAI22_X1  g146(.A1(new_n506), .A2(new_n570), .B1(new_n508), .B2(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n501), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n573));
  OAI21_X1  g148(.A(KEYINPUT71), .B1(new_n573), .B2(new_n503), .ZN(new_n574));
  OAI21_X1  g149(.A(G61), .B1(new_n516), .B2(new_n517), .ZN(new_n575));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT71), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n577), .A2(new_n578), .A3(G651), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n572), .B1(new_n574), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G305));
  AOI22_X1  g156(.A1(new_n552), .A2(G85), .B1(new_n549), .B2(G47), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT72), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n501), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n584), .A2(new_n503), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n583), .A2(new_n585), .ZN(G290));
  NAND2_X1  g161(.A1(G301), .A2(G868), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n552), .A2(G92), .ZN(new_n588));
  XOR2_X1   g163(.A(new_n588), .B(KEYINPUT10), .Z(new_n589));
  NAND2_X1  g164(.A1(G79), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G66), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n518), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n592), .A2(G651), .B1(G54), .B2(new_n549), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n587), .B1(new_n595), .B2(G868), .ZN(G284));
  OAI21_X1  g171(.A(new_n587), .B1(new_n595), .B2(G868), .ZN(G321));
  MUX2_X1   g172(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g173(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n595), .B1(new_n600), .B2(G860), .ZN(G148));
  NAND2_X1  g176(.A1(new_n595), .A2(new_n600), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G868), .B2(new_n534), .ZN(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g180(.A(new_n481), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n606), .A2(new_n468), .ZN(new_n607));
  XOR2_X1   g182(.A(new_n607), .B(KEYINPUT12), .Z(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT13), .ZN(new_n609));
  XOR2_X1   g184(.A(KEYINPUT73), .B(G2100), .Z(new_n610));
  OR2_X1    g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n609), .A2(new_n610), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n476), .A2(G123), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n463), .A2(G111), .ZN(new_n614));
  OAI21_X1  g189(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n615));
  INV_X1    g190(.A(G135), .ZN(new_n616));
  OAI221_X1 g191(.A(new_n613), .B1(new_n614), .B2(new_n615), .C1(new_n616), .C2(new_n482), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(G2096), .Z(new_n618));
  NAND3_X1  g193(.A1(new_n611), .A2(new_n612), .A3(new_n618), .ZN(G156));
  XNOR2_X1  g194(.A(G2427), .B(G2438), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2430), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT15), .B(G2435), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n623), .A2(KEYINPUT14), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(G1341), .B(G1348), .Z(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n625), .B(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(G2451), .B(G2454), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT75), .ZN(new_n632));
  XOR2_X1   g207(.A(G2443), .B(G2446), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  OAI21_X1  g210(.A(G14), .B1(new_n630), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n636), .B1(new_n635), .B2(new_n630), .ZN(G401));
  XOR2_X1   g212(.A(G2072), .B(G2078), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT76), .ZN(new_n639));
  XOR2_X1   g214(.A(KEYINPUT78), .B(KEYINPUT17), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2067), .B(G2678), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(KEYINPUT77), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2084), .B(G2090), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(new_n639), .B2(new_n642), .ZN(new_n646));
  OAI22_X1  g221(.A1(new_n641), .A2(new_n643), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n647), .B1(new_n644), .B2(new_n646), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT79), .Z(new_n649));
  NOR2_X1   g224(.A1(new_n643), .A2(new_n645), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n639), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT18), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n645), .A2(new_n642), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n652), .B1(new_n641), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n649), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2096), .B(G2100), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(G227));
  XOR2_X1   g233(.A(G1956), .B(G2474), .Z(new_n659));
  XOR2_X1   g234(.A(G1961), .B(G1966), .Z(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n661), .A2(KEYINPUT80), .ZN(new_n662));
  XOR2_X1   g237(.A(G1971), .B(G1976), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n661), .A2(KEYINPUT80), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n662), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(KEYINPUT81), .B(KEYINPUT20), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n659), .A2(new_n660), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n664), .A2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n669), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(new_n661), .ZN(new_n672));
  OAI211_X1 g247(.A(new_n668), .B(new_n670), .C1(new_n664), .C2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G1991), .B(G1996), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1981), .B(G1986), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(G229));
  NOR2_X1   g255(.A1(G16), .A2(G24), .ZN(new_n681));
  XNOR2_X1  g256(.A(G290), .B(KEYINPUT83), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n681), .B1(new_n682), .B2(G16), .ZN(new_n683));
  INV_X1    g258(.A(G1986), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n476), .A2(G119), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n463), .A2(G107), .ZN(new_n687));
  OAI21_X1  g262(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n688));
  INV_X1    g263(.A(G131), .ZN(new_n689));
  OAI221_X1 g264(.A(new_n686), .B1(new_n687), .B2(new_n688), .C1(new_n689), .C2(new_n482), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT82), .Z(new_n691));
  MUX2_X1   g266(.A(G25), .B(new_n691), .S(G29), .Z(new_n692));
  XOR2_X1   g267(.A(KEYINPUT35), .B(G1991), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G22), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(G166), .B2(new_n695), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(G1971), .Z(new_n698));
  NAND2_X1  g273(.A1(new_n695), .A2(G6), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(new_n580), .B2(new_n695), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT32), .B(G1981), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n695), .A2(G23), .ZN(new_n704));
  INV_X1    g279(.A(G288), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n704), .B1(new_n705), .B2(new_n695), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT33), .B(G1976), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT84), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n706), .B(new_n708), .ZN(new_n709));
  NAND4_X1  g284(.A1(new_n698), .A2(new_n702), .A3(new_n703), .A4(new_n709), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n685), .B(new_n694), .C1(KEYINPUT34), .C2(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT85), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(KEYINPUT34), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT36), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n715), .A2(KEYINPUT86), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n712), .B(new_n713), .C1(KEYINPUT86), .C2(new_n715), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G32), .ZN(new_n721));
  NAND3_X1  g296(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT26), .Z(new_n723));
  NAND2_X1  g298(.A1(new_n481), .A2(G2105), .ZN(new_n724));
  INV_X1    g299(.A(G129), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G141), .ZN(new_n727));
  INV_X1    g302(.A(G105), .ZN(new_n728));
  OAI22_X1  g303(.A1(new_n482), .A2(new_n727), .B1(new_n728), .B2(new_n468), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n721), .B1(new_n730), .B2(new_n720), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT27), .B(G1996), .Z(new_n732));
  NAND2_X1  g307(.A1(new_n695), .A2(G5), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G171), .B2(new_n695), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n731), .A2(new_n732), .B1(new_n734), .B2(G1961), .ZN(new_n735));
  INV_X1    g310(.A(G1966), .ZN(new_n736));
  NOR2_X1   g311(.A1(G168), .A2(new_n695), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n695), .B2(G21), .ZN(new_n738));
  INV_X1    g313(.A(G34), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n739), .A2(KEYINPUT24), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n739), .A2(KEYINPUT24), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n720), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G160), .B2(new_n720), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT94), .Z(new_n744));
  INV_X1    g319(.A(G2084), .ZN(new_n745));
  OAI221_X1 g320(.A(new_n735), .B1(new_n736), .B2(new_n738), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n738), .A2(new_n736), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT31), .B(G11), .ZN(new_n748));
  INV_X1    g323(.A(G28), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n749), .A2(KEYINPUT30), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT30), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n720), .B1(new_n751), .B2(G28), .ZN(new_n752));
  OAI221_X1 g327(.A(new_n748), .B1(new_n750), .B2(new_n752), .C1(new_n617), .C2(new_n720), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n734), .A2(G1961), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n731), .A2(new_n732), .ZN(new_n755));
  NOR4_X1   g330(.A1(new_n747), .A2(new_n753), .A3(new_n754), .A4(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n695), .A2(G20), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT23), .Z(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G299), .B2(G16), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(G1956), .ZN(new_n760));
  NOR2_X1   g335(.A1(G27), .A2(G29), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G164), .B2(G29), .ZN(new_n762));
  INV_X1    g337(.A(G2078), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n756), .A2(new_n760), .A3(new_n764), .ZN(new_n765));
  AOI211_X1 g340(.A(new_n746), .B(new_n765), .C1(new_n745), .C2(new_n744), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT25), .Z(new_n768));
  INV_X1    g343(.A(G139), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n769), .B2(new_n482), .ZN(new_n770));
  NAND2_X1  g345(.A1(G115), .A2(G2104), .ZN(new_n771));
  INV_X1    g346(.A(G127), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n771), .B1(new_n606), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n770), .B1(G2105), .B2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT92), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT93), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n777), .A2(G29), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G29), .B2(G33), .ZN(new_n779));
  INV_X1    g354(.A(G2072), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n720), .A2(G35), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT95), .Z(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n484), .B2(G29), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT29), .Z(new_n785));
  AOI22_X1  g360(.A1(new_n779), .A2(new_n780), .B1(G2090), .B2(new_n785), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n785), .A2(G2090), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n766), .A2(new_n781), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(G16), .A2(G19), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n534), .B2(G16), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT88), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(G1341), .Z(new_n792));
  NAND2_X1  g367(.A1(new_n720), .A2(G26), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT28), .Z(new_n794));
  OR2_X1    g369(.A1(G104), .A2(G2105), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n795), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT89), .ZN(new_n797));
  INV_X1    g372(.A(G128), .ZN(new_n798));
  INV_X1    g373(.A(G140), .ZN(new_n799));
  OAI22_X1  g374(.A1(new_n798), .A2(new_n724), .B1(new_n482), .B2(new_n799), .ZN(new_n800));
  OR3_X1    g375(.A1(new_n797), .A2(new_n800), .A3(KEYINPUT90), .ZN(new_n801));
  OAI21_X1  g376(.A(KEYINPUT90), .B1(new_n797), .B2(new_n800), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n794), .B1(new_n803), .B2(G29), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G2067), .ZN(new_n805));
  NOR2_X1   g380(.A1(G4), .A2(G16), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT87), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n594), .B2(new_n695), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G1348), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n792), .A2(new_n805), .A3(new_n809), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT91), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n788), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n719), .A2(new_n812), .ZN(G150));
  INV_X1    g388(.A(G150), .ZN(G311));
  NAND2_X1  g389(.A1(new_n595), .A2(G559), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT96), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT38), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n501), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n818), .A2(new_n503), .ZN(new_n819));
  INV_X1    g394(.A(G93), .ZN(new_n820));
  INV_X1    g395(.A(G55), .ZN(new_n821));
  OAI22_X1  g396(.A1(new_n506), .A2(new_n820), .B1(new_n508), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n534), .B(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n817), .B(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT39), .ZN(new_n826));
  AOI21_X1  g401(.A(G860), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(new_n826), .B2(new_n825), .ZN(new_n828));
  OAI21_X1  g403(.A(G860), .B1(new_n819), .B2(new_n822), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT37), .Z(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n830), .ZN(G145));
  XOR2_X1   g406(.A(new_n690), .B(KEYINPUT100), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(new_n608), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n476), .A2(G130), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n481), .A2(G142), .A3(new_n463), .ZN(new_n836));
  OR2_X1    g411(.A1(G106), .A2(G2105), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n837), .B(G2104), .C1(G118), .C2(new_n463), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n835), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n803), .A2(G164), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n803), .A2(G164), .ZN(new_n842));
  OAI22_X1  g417(.A1(new_n841), .A2(new_n842), .B1(new_n729), .B2(new_n726), .ZN(new_n843));
  INV_X1    g418(.A(new_n842), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n844), .A2(new_n730), .A3(new_n840), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(new_n777), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT99), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n843), .A2(new_n845), .A3(new_n848), .A4(new_n776), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n843), .A2(new_n845), .A3(new_n776), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(KEYINPUT99), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n839), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n853), .ZN(new_n855));
  INV_X1    g430(.A(new_n839), .ZN(new_n856));
  NOR3_X1   g431(.A1(new_n855), .A2(new_n850), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n834), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n851), .A2(new_n839), .A3(new_n853), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n856), .B1(new_n855), .B2(new_n850), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n859), .A2(new_n833), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n484), .B(new_n617), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(G160), .Z(new_n864));
  XNOR2_X1  g439(.A(KEYINPUT97), .B(KEYINPUT98), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(G37), .B1(new_n862), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n866), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n858), .A2(new_n868), .A3(new_n861), .ZN(new_n869));
  AOI21_X1  g444(.A(KEYINPUT40), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  AND3_X1   g445(.A1(new_n859), .A2(new_n833), .A3(new_n860), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n833), .B1(new_n859), .B2(new_n860), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n866), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(G37), .ZN(new_n874));
  AND4_X1   g449(.A1(KEYINPUT40), .A2(new_n873), .A3(new_n874), .A4(new_n869), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n870), .A2(new_n875), .ZN(G395));
  XNOR2_X1  g451(.A(G290), .B(new_n580), .ZN(new_n877));
  XNOR2_X1  g452(.A(G166), .B(new_n705), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n880), .A2(KEYINPUT42), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n879), .B(KEYINPUT102), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n881), .B1(new_n882), .B2(KEYINPUT42), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n594), .B(G299), .ZN(new_n884));
  XOR2_X1   g459(.A(KEYINPUT101), .B(KEYINPUT41), .Z(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n887), .B1(KEYINPUT41), .B2(new_n884), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n602), .B(new_n824), .Z(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n890), .B1(new_n889), .B2(new_n884), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n883), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n883), .A2(new_n891), .ZN(new_n893));
  OAI21_X1  g468(.A(G868), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n823), .A2(G868), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n894), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n895), .B1(new_n894), .B2(new_n897), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(G295));
  NAND2_X1  g475(.A1(new_n894), .A2(new_n897), .ZN(G331));
  XNOR2_X1  g476(.A(new_n824), .B(G171), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(G168), .ZN(new_n903));
  OR2_X1    g478(.A1(new_n903), .A2(new_n884), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n888), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(G37), .B1(new_n906), .B2(new_n882), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT43), .ZN(new_n908));
  INV_X1    g483(.A(new_n882), .ZN(new_n909));
  MUX2_X1   g484(.A(new_n885), .B(KEYINPUT41), .S(new_n884), .Z(new_n910));
  NAND3_X1  g485(.A1(new_n903), .A2(new_n910), .A3(KEYINPUT104), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n904), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(KEYINPUT104), .B1(new_n903), .B2(new_n910), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n909), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n907), .A2(new_n908), .A3(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n906), .A2(new_n882), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n904), .A2(new_n905), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n874), .B1(new_n917), .B2(new_n909), .ZN(new_n918));
  OAI21_X1  g493(.A(KEYINPUT43), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n915), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n907), .A2(KEYINPUT43), .A3(new_n914), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n908), .B1(new_n916), .B2(new_n918), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  MUX2_X1   g498(.A(new_n920), .B(new_n923), .S(KEYINPUT44), .Z(G397));
  XOR2_X1   g499(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n925));
  OAI21_X1  g500(.A(new_n925), .B1(G164), .B2(G1384), .ZN(new_n926));
  NAND2_X1  g501(.A1(G160), .A2(G40), .ZN(new_n927));
  NOR3_X1   g502(.A1(new_n926), .A2(G1996), .A3(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(KEYINPUT46), .ZN(new_n929));
  INV_X1    g504(.A(G2067), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n803), .B(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n730), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n926), .A2(new_n927), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n929), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n934), .B(KEYINPUT47), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n730), .B(G1996), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n931), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n693), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n937), .A2(new_n691), .A3(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n803), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n939), .B1(new_n930), .B2(new_n940), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n941), .A2(new_n927), .A3(new_n926), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n690), .B(new_n938), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n933), .B1(new_n937), .B2(new_n943), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n933), .A2(new_n684), .A3(new_n585), .A4(new_n583), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n945), .B(KEYINPUT48), .ZN(new_n946));
  AOI211_X1 g521(.A(new_n935), .B(new_n942), .C1(new_n944), .C2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(G290), .A2(G1986), .A3(new_n933), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n945), .ZN(new_n949));
  XOR2_X1   g524(.A(new_n949), .B(KEYINPUT106), .Z(new_n950));
  AND2_X1   g525(.A1(new_n950), .A2(new_n944), .ZN(new_n951));
  INV_X1    g526(.A(G1981), .ZN(new_n952));
  AOI22_X1  g527(.A1(new_n552), .A2(G86), .B1(new_n549), .B2(G48), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n577), .A2(G651), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n955), .B1(new_n580), .B2(new_n952), .ZN(new_n956));
  XOR2_X1   g531(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n957));
  OAI21_X1  g532(.A(KEYINPUT111), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT111), .ZN(new_n959));
  INV_X1    g534(.A(new_n957), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n578), .B1(new_n577), .B2(G651), .ZN(new_n961));
  AOI211_X1 g536(.A(KEYINPUT71), .B(new_n503), .C1(new_n575), .C2(new_n576), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n952), .B(new_n953), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n959), .B(new_n960), .C1(new_n964), .C2(new_n955), .ZN(new_n965));
  INV_X1    g540(.A(G8), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n495), .A2(new_n497), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n486), .A2(new_n490), .ZN(new_n968));
  AOI21_X1  g543(.A(G1384), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(G40), .ZN(new_n970));
  NOR3_X1   g545(.A1(new_n469), .A2(new_n472), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n966), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n956), .A2(KEYINPUT49), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n958), .A2(new_n965), .A3(new_n972), .A4(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n705), .A2(G1976), .ZN(new_n975));
  INV_X1    g550(.A(G1976), .ZN(new_n976));
  AOI21_X1  g551(.A(KEYINPUT52), .B1(G288), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n972), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n972), .A2(KEYINPUT109), .A3(new_n975), .A4(new_n977), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n972), .A2(new_n975), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT108), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT108), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n972), .A2(new_n985), .A3(new_n975), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n984), .A2(KEYINPUT52), .A3(new_n986), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n974), .A2(new_n982), .A3(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n925), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n969), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n992), .B1(G164), .B2(G1384), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n991), .A2(new_n993), .A3(new_n971), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n736), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n967), .A2(new_n968), .ZN(new_n997));
  INV_X1    g572(.A(G1384), .ZN(new_n998));
  XNOR2_X1  g573(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n996), .A2(new_n1000), .A3(new_n745), .A4(new_n971), .ZN(new_n1001));
  AOI211_X1 g576(.A(new_n966), .B(G286), .C1(new_n995), .C2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n997), .A2(KEYINPUT45), .A3(new_n998), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n926), .A2(new_n1003), .A3(new_n971), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n996), .A2(new_n1000), .A3(new_n971), .ZN(new_n1005));
  OAI22_X1  g580(.A1(new_n1004), .A2(G1971), .B1(new_n1005), .B2(G2090), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n1006), .A2(G8), .ZN(new_n1007));
  NOR2_X1   g582(.A1(G166), .A2(new_n966), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n1008), .B(KEYINPUT55), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1002), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(KEYINPUT63), .B1(new_n989), .B2(new_n1010), .ZN(new_n1011));
  AND3_X1   g586(.A1(new_n974), .A2(new_n976), .A3(new_n705), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n972), .B1(new_n1012), .B2(new_n964), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT50), .ZN(new_n1015));
  INV_X1    g590(.A(new_n497), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n496), .B1(new_n481), .B2(new_n493), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1015), .B(new_n998), .C1(new_n1018), .C2(new_n491), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT112), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n969), .A2(KEYINPUT112), .A3(new_n1015), .ZN(new_n1022));
  INV_X1    g597(.A(new_n999), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(G164), .B2(G1384), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1021), .A2(new_n1022), .A3(new_n971), .A4(new_n1024), .ZN(new_n1025));
  OAI22_X1  g600(.A1(new_n1025), .A2(G2090), .B1(new_n1004), .B2(G1971), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(G8), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1009), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT63), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1029), .A2(new_n1030), .A3(new_n1002), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1006), .A2(new_n1009), .A3(G8), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n989), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1014), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n1035));
  INV_X1    g610(.A(G1956), .ZN(new_n1036));
  XNOR2_X1  g611(.A(KEYINPUT56), .B(G2072), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n1025), .A2(new_n1036), .B1(new_n1004), .B2(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g613(.A(KEYINPUT113), .B(KEYINPUT57), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n553), .A2(new_n561), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1039), .B1(new_n553), .B2(new_n561), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT114), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1039), .ZN(new_n1043));
  NAND2_X1  g618(.A1(G299), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT114), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n553), .A2(new_n561), .A3(new_n1039), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n1042), .A2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1035), .B1(new_n1038), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1042), .A2(new_n1047), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n971), .B1(new_n969), .B2(new_n999), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT112), .B1(new_n969), .B2(new_n1015), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(G1956), .B1(new_n1053), .B2(new_n1022), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n926), .A2(new_n1003), .A3(new_n971), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1037), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g632(.A(KEYINPUT115), .B(new_n1050), .C1(new_n1054), .C2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1049), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G1348), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n969), .A2(new_n971), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  AOI22_X1  g637(.A1(new_n1005), .A2(new_n1060), .B1(new_n1062), .B2(new_n930), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1063), .A2(new_n594), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1059), .A2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1038), .A2(new_n1067), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1005), .A2(new_n1060), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1062), .A2(new_n930), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(KEYINPUT60), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(new_n595), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT118), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1063), .A2(KEYINPUT117), .A3(KEYINPUT60), .A4(new_n594), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1070), .A2(KEYINPUT60), .A3(new_n594), .A4(new_n1071), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT117), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT118), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1072), .A2(new_n1079), .A3(new_n595), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1074), .A2(new_n1075), .A3(new_n1078), .A4(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1063), .A2(KEYINPUT60), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1081), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1082), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  OAI22_X1  g662(.A1(new_n1054), .A2(new_n1057), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(new_n1068), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT61), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT58), .B(G1341), .ZN(new_n1092));
  OAI22_X1  g667(.A1(new_n1055), .A2(G1996), .B1(new_n1062), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n534), .ZN(new_n1094));
  XNOR2_X1  g669(.A(new_n1094), .B(KEYINPUT59), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1091), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1090), .B1(new_n1038), .B2(new_n1067), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1059), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT116), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1059), .A2(KEYINPUT116), .A3(new_n1097), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1096), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1069), .B1(new_n1087), .B2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n926), .A2(new_n1003), .A3(new_n763), .A4(new_n971), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT122), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1104), .A2(KEYINPUT122), .A3(new_n1105), .ZN(new_n1108));
  INV_X1    g683(.A(G1961), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1107), .A2(new_n1108), .B1(new_n1109), .B2(new_n1005), .ZN(new_n1110));
  OR3_X1    g685(.A1(new_n994), .A2(new_n1105), .A3(G2078), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1110), .A2(G301), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT125), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1110), .A2(KEYINPUT125), .A3(G301), .A4(new_n1111), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1005), .A2(new_n1109), .ZN(new_n1118));
  AOI211_X1 g693(.A(new_n1105), .B(G2078), .C1(new_n927), .C2(KEYINPUT123), .ZN(new_n1119));
  OR2_X1    g694(.A1(new_n927), .A2(KEYINPUT123), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1119), .A2(new_n926), .A3(new_n1003), .A4(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1108), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1118), .B(new_n1121), .C1(new_n1122), .C2(new_n1106), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1117), .B1(new_n1123), .B2(G171), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1116), .A2(new_n1124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1032), .A2(new_n974), .A3(new_n982), .A4(new_n987), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1009), .B1(new_n1026), .B2(G8), .ZN(new_n1127));
  OAI21_X1  g702(.A(KEYINPUT124), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n988), .A2(new_n1029), .A3(new_n1129), .A4(new_n1032), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(G301), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1123), .A2(G171), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1117), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT121), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n995), .A2(new_n1001), .A3(G168), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT51), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n966), .A2(KEYINPUT120), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n995), .A2(new_n1001), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1140), .A2(G8), .A3(G286), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1137), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1135), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(KEYINPUT51), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1146), .A2(KEYINPUT121), .A3(new_n1141), .A4(new_n1139), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1125), .A2(new_n1131), .A3(new_n1134), .A4(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1034), .B1(new_n1103), .B2(new_n1149), .ZN(new_n1150));
  AND3_X1   g725(.A1(new_n1128), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1148), .A2(KEYINPUT62), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT62), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1144), .A2(new_n1153), .A3(new_n1147), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1151), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT126), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1151), .A2(new_n1152), .A3(KEYINPUT126), .A4(new_n1154), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  OAI211_X1 g734(.A(KEYINPUT127), .B(new_n951), .C1(new_n1150), .C2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1069), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1078), .A2(new_n1075), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1079), .B1(new_n1072), .B2(new_n595), .ZN(new_n1164));
  AOI211_X1 g739(.A(KEYINPUT118), .B(new_n594), .C1(new_n1063), .C2(KEYINPUT60), .ZN(new_n1165));
  NOR3_X1   g740(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(KEYINPUT119), .B1(new_n1166), .B2(new_n1083), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1081), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT59), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1094), .B(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1171), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1172));
  AND3_X1   g747(.A1(new_n1059), .A2(KEYINPUT116), .A3(new_n1097), .ZN(new_n1173));
  AOI21_X1  g748(.A(KEYINPUT116), .B1(new_n1059), .B2(new_n1097), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1172), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1162), .B1(new_n1169), .B2(new_n1175), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1148), .A2(new_n1134), .A3(new_n1128), .A4(new_n1130), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1124), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1178), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1176), .A2(new_n1180), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1181), .A2(new_n1034), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1182));
  AOI21_X1  g757(.A(KEYINPUT127), .B1(new_n1182), .B2(new_n951), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n947), .B1(new_n1161), .B2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g759(.A1(new_n867), .A2(new_n869), .ZN(new_n1186));
  NOR2_X1   g760(.A1(G401), .A2(new_n461), .ZN(new_n1187));
  NAND3_X1  g761(.A1(new_n679), .A2(new_n657), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g762(.A(new_n1188), .B1(new_n915), .B2(new_n919), .ZN(new_n1189));
  NAND2_X1  g763(.A1(new_n1186), .A2(new_n1189), .ZN(G225));
  INV_X1    g764(.A(G225), .ZN(G308));
endmodule


