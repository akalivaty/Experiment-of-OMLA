//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 1 1 1 1 0 1 0 1 0 0 1 1 0 0 0 0 0 1 0 0 1 1 0 0 0 0 1 0 0 0 1 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n494, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n593, new_n594,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n654, new_n657, new_n659, new_n660, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1214,
    new_n1215;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT64), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  NAND2_X1  g032(.A1(G113), .A2(G2104), .ZN(new_n458));
  INV_X1    g033(.A(G125), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT65), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n461), .A2(new_n463), .A3(KEYINPUT65), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n459), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n458), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AND3_X1   g045(.A1(new_n461), .A2(new_n463), .A3(KEYINPUT65), .ZN(new_n471));
  AOI21_X1  g046(.A(KEYINPUT65), .B1(new_n461), .B2(new_n463), .ZN(new_n472));
  OAI21_X1  g047(.A(G125), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(KEYINPUT66), .ZN(new_n474));
  OAI21_X1  g049(.A(G2105), .B1(new_n470), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT67), .ZN(new_n476));
  AOI22_X1  g051(.A1(new_n473), .A2(KEYINPUT66), .B1(G113), .B2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n468), .A2(new_n469), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n479), .A2(new_n480), .A3(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g057(.A(KEYINPUT68), .B(G2104), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  AND3_X1   g059(.A1(new_n484), .A2(KEYINPUT69), .A3(G101), .ZN(new_n485));
  AOI21_X1  g060(.A(KEYINPUT69), .B1(new_n484), .B2(G101), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n461), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n488), .B1(new_n483), .B2(KEYINPUT3), .ZN(new_n489));
  INV_X1    g064(.A(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n487), .B1(G137), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n482), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G160));
  NAND2_X1  g070(.A1(new_n492), .A2(G136), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n489), .A2(G2105), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G124), .ZN(new_n498));
  OR2_X1    g073(.A1(G100), .A2(G2105), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n499), .B(G2104), .C1(G112), .C2(new_n490), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n496), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G162));
  NAND2_X1  g077(.A1(new_n466), .A2(new_n467), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n490), .A2(G138), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g080(.A(KEYINPUT4), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G114), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n462), .B1(new_n507), .B2(G2105), .ZN(new_n508));
  NOR2_X1   g083(.A1(G102), .A2(G2105), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n508), .A2(KEYINPUT70), .A3(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT70), .ZN(new_n512));
  OAI21_X1  g087(.A(G2104), .B1(new_n490), .B2(G114), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n512), .B1(new_n513), .B2(new_n509), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(G126), .A2(G2105), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT4), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n516), .B1(new_n504), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n462), .A2(KEYINPUT68), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT68), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G2104), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n519), .A2(new_n521), .A3(KEYINPUT3), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n518), .A2(new_n522), .A3(new_n461), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n515), .A2(new_n523), .ZN(new_n524));
  NOR3_X1   g099(.A1(new_n506), .A2(new_n524), .A3(KEYINPUT71), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT71), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n471), .A2(new_n472), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n517), .B1(new_n527), .B2(new_n504), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n489), .A2(new_n518), .B1(new_n511), .B2(new_n514), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n526), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n525), .A2(new_n530), .ZN(G164));
  INV_X1    g106(.A(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT72), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT72), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT5), .ZN(new_n537));
  OAI21_X1  g112(.A(G543), .B1(new_n537), .B2(KEYINPUT73), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT73), .ZN(new_n539));
  INV_X1    g114(.A(G543), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n539), .A2(new_n540), .A3(KEYINPUT5), .ZN(new_n541));
  AND2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n542), .A2(G62), .ZN(new_n543));
  NAND2_X1  g118(.A1(G75), .A2(G543), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT74), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n536), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(KEYINPUT6), .A2(G651), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n547), .B1(new_n536), .B2(KEYINPUT6), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n538), .A2(new_n541), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G88), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n548), .A2(new_n540), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G50), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n546), .A2(new_n551), .A3(new_n553), .ZN(G303));
  INV_X1    g129(.A(G303), .ZN(G166));
  INV_X1    g130(.A(KEYINPUT76), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n556), .B1(new_n548), .B2(new_n540), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT6), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n558), .B1(new_n533), .B2(new_n535), .ZN(new_n559));
  OAI211_X1 g134(.A(KEYINPUT76), .B(G543), .C1(new_n559), .C2(new_n547), .ZN(new_n560));
  AND2_X1   g135(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  AND2_X1   g136(.A1(new_n561), .A2(G51), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n550), .A2(G89), .ZN(new_n563));
  NAND3_X1  g138(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT7), .ZN(new_n565));
  AND3_X1   g140(.A1(new_n538), .A2(new_n541), .A3(KEYINPUT75), .ZN(new_n566));
  AOI21_X1  g141(.A(KEYINPUT75), .B1(new_n538), .B2(new_n541), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(G63), .A2(G651), .ZN(new_n569));
  OAI211_X1 g144(.A(new_n563), .B(new_n565), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n562), .A2(new_n570), .ZN(G168));
  INV_X1    g146(.A(G64), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n549), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n538), .A2(new_n541), .A3(KEYINPUT75), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n572), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AND2_X1   g151(.A1(G77), .A2(G543), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n536), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n557), .A2(G52), .A3(new_n560), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n550), .A2(G90), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G301));
  INV_X1    g156(.A(G301), .ZN(G171));
  INV_X1    g157(.A(G56), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n583), .B1(new_n574), .B2(new_n575), .ZN(new_n584));
  AND2_X1   g159(.A1(G68), .A2(G543), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n536), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n557), .A2(G43), .A3(new_n560), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n550), .A2(G81), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(G860), .ZN(G153));
  NAND4_X1  g166(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g167(.A1(G1), .A2(G3), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n593), .B(KEYINPUT8), .ZN(new_n594));
  NAND4_X1  g169(.A1(G319), .A2(G483), .A3(G661), .A4(new_n594), .ZN(G188));
  INV_X1    g170(.A(G53), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n596), .B1(KEYINPUT77), .B2(KEYINPUT9), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n552), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g173(.A1(KEYINPUT77), .A2(KEYINPUT9), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g175(.A(new_n552), .B(new_n597), .C1(KEYINPUT77), .C2(KEYINPUT9), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n542), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n602), .A2(new_n532), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n550), .A2(G91), .ZN(new_n604));
  NAND4_X1  g179(.A1(new_n600), .A2(new_n601), .A3(new_n603), .A4(new_n604), .ZN(G299));
  INV_X1    g180(.A(G168), .ZN(G286));
  INV_X1    g181(.A(G74), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n574), .A2(new_n607), .A3(new_n575), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G651), .ZN(new_n609));
  OAI211_X1 g184(.A(new_n542), .B(G87), .C1(new_n559), .C2(new_n547), .ZN(new_n610));
  OAI211_X1 g185(.A(G49), .B(G543), .C1(new_n559), .C2(new_n547), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(G288));
  OAI211_X1 g187(.A(G48), .B(G543), .C1(new_n559), .C2(new_n547), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT78), .ZN(new_n614));
  NAND2_X1  g189(.A1(G73), .A2(G543), .ZN(new_n615));
  INV_X1    g190(.A(G61), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n549), .B2(new_n616), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n550), .A2(G86), .B1(new_n536), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n614), .A2(new_n618), .ZN(G305));
  INV_X1    g194(.A(G60), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n620), .B1(new_n574), .B2(new_n575), .ZN(new_n621));
  AND2_X1   g196(.A1(G72), .A2(G543), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n536), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(KEYINPUT79), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI211_X1 g200(.A(KEYINPUT79), .B(new_n536), .C1(new_n621), .C2(new_n622), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n557), .A2(G47), .A3(new_n560), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n550), .A2(G85), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(KEYINPUT80), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT80), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n628), .A2(new_n632), .A3(new_n629), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n627), .A2(new_n631), .A3(new_n633), .ZN(G290));
  INV_X1    g209(.A(G868), .ZN(new_n635));
  NOR2_X1   g210(.A1(G301), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n550), .A2(G92), .ZN(new_n637));
  INV_X1    g212(.A(KEYINPUT10), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n550), .A2(KEYINPUT10), .A3(G92), .ZN(new_n640));
  NAND2_X1  g215(.A1(G79), .A2(G543), .ZN(new_n641));
  INV_X1    g216(.A(G66), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n641), .B1(new_n549), .B2(new_n642), .ZN(new_n643));
  AOI22_X1  g218(.A1(new_n639), .A2(new_n640), .B1(G651), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n561), .A2(G54), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(KEYINPUT81), .ZN(new_n647));
  INV_X1    g222(.A(KEYINPUT81), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n644), .A2(new_n648), .A3(new_n645), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n636), .B1(new_n651), .B2(new_n635), .ZN(G284));
  AOI21_X1  g227(.A(new_n636), .B1(new_n651), .B2(new_n635), .ZN(G321));
  NAND2_X1  g228(.A1(G299), .A2(new_n635), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(G168), .B2(new_n635), .ZN(G297));
  OAI21_X1  g230(.A(new_n654), .B1(G168), .B2(new_n635), .ZN(G280));
  INV_X1    g231(.A(G559), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n651), .B1(new_n657), .B2(G860), .ZN(G148));
  NAND3_X1  g233(.A1(new_n647), .A2(new_n657), .A3(new_n649), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(G868), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n660), .B1(G868), .B2(new_n590), .ZN(G323));
  XNOR2_X1  g236(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g237(.A1(new_n503), .A2(new_n484), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT12), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT13), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT82), .B(G2100), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n492), .A2(G135), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n497), .A2(G123), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT83), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n670), .A2(new_n490), .A3(G111), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n670), .B1(new_n490), .B2(G111), .ZN(new_n672));
  OR2_X1    g247(.A1(G99), .A2(G2105), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n672), .A2(G2104), .A3(new_n673), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n668), .B(new_n669), .C1(new_n671), .C2(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(KEYINPUT84), .B(G2096), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n667), .A2(new_n677), .ZN(G156));
  XNOR2_X1  g253(.A(G2427), .B(G2438), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(G2430), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT15), .B(G2435), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n680), .A2(new_n681), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n682), .A2(KEYINPUT14), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G1341), .B(G1348), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G2451), .B(G2454), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n687), .B(new_n688), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n686), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G2443), .B(G2446), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT86), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n690), .A2(new_n692), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n693), .A2(G14), .A3(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(G401));
  XOR2_X1   g271(.A(G2084), .B(G2090), .Z(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(G2072), .A2(G2078), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n442), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G2067), .B(G2678), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  NOR3_X1   g277(.A1(new_n698), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT18), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n701), .B1(KEYINPUT87), .B2(new_n700), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(KEYINPUT87), .B2(new_n700), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n700), .B(KEYINPUT17), .ZN(new_n707));
  OAI211_X1 g282(.A(new_n706), .B(new_n698), .C1(new_n707), .C2(new_n702), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n707), .A2(new_n702), .A3(new_n697), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n704), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(G2096), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(G2100), .ZN(G227));
  XOR2_X1   g287(.A(G1971), .B(G1976), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT19), .ZN(new_n714));
  XNOR2_X1  g289(.A(G1956), .B(G2474), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  XOR2_X1   g291(.A(G1961), .B(G1966), .Z(new_n717));
  AND2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT20), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n716), .A2(new_n717), .ZN(new_n721));
  NOR3_X1   g296(.A1(new_n714), .A2(new_n718), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n714), .B2(new_n721), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT88), .Z(new_n726));
  XNOR2_X1  g301(.A(new_n724), .B(new_n726), .ZN(new_n727));
  XOR2_X1   g302(.A(G1981), .B(G1986), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(G1991), .B(G1996), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(G229));
  INV_X1    g306(.A(G29), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G33), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n490), .A2(G103), .A3(G2104), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT97), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT25), .Z(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G139), .B2(new_n492), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n503), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n738), .A2(new_n490), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n733), .B1(new_n741), .B2(new_n732), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G2072), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n675), .A2(new_n732), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n744), .A2(KEYINPUT102), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n744), .A2(KEYINPUT102), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT30), .ZN(new_n747));
  AND2_X1   g322(.A1(new_n747), .A2(G28), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n732), .B1(new_n747), .B2(G28), .ZN(new_n749));
  AND2_X1   g324(.A1(KEYINPUT31), .A2(G11), .ZN(new_n750));
  NOR2_X1   g325(.A1(KEYINPUT31), .A2(G11), .ZN(new_n751));
  OAI22_X1  g326(.A1(new_n748), .A2(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NOR4_X1   g327(.A1(new_n743), .A2(new_n745), .A3(new_n746), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n732), .A2(G32), .ZN(new_n754));
  AOI22_X1  g329(.A1(new_n492), .A2(G141), .B1(G105), .B2(new_n484), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n497), .A2(G129), .ZN(new_n756));
  NAND3_X1  g331(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT99), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT26), .ZN(new_n759));
  AND3_X1   g334(.A1(new_n755), .A2(new_n756), .A3(new_n759), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT100), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n754), .B1(new_n762), .B2(new_n732), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT27), .B(G1996), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n732), .A2(G35), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G162), .B2(new_n732), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT29), .B(G2090), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(G16), .ZN(new_n770));
  NOR2_X1   g345(.A1(G168), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n770), .B2(G21), .ZN(new_n772));
  INV_X1    g347(.A(G1966), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n769), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n753), .A2(new_n765), .A3(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(G4), .A2(G16), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT93), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n650), .B2(new_n770), .ZN(new_n778));
  INV_X1    g353(.A(G1348), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n772), .A2(new_n773), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT101), .ZN(new_n782));
  NOR3_X1   g357(.A1(new_n775), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n732), .B1(KEYINPUT24), .B2(G34), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(KEYINPUT24), .B2(G34), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n494), .B2(G29), .ZN(new_n786));
  INV_X1    g361(.A(G2084), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT98), .Z(new_n789));
  NAND2_X1  g364(.A1(new_n770), .A2(G20), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT23), .ZN(new_n791));
  INV_X1    g366(.A(G299), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(new_n770), .ZN(new_n793));
  INV_X1    g368(.A(G1956), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n770), .A2(G19), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT94), .Z(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n590), .B2(new_n770), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT95), .B(G1341), .Z(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n770), .A2(G5), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G171), .B2(new_n770), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n795), .B(new_n800), .C1(G1961), .C2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n732), .A2(G26), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT28), .Z(new_n805));
  NAND2_X1  g380(.A1(new_n497), .A2(G128), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT96), .Z(new_n807));
  OR2_X1    g382(.A1(G104), .A2(G2105), .ZN(new_n808));
  INV_X1    g383(.A(G116), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n462), .B1(new_n809), .B2(G2105), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n492), .A2(G140), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n805), .B1(new_n812), .B2(G29), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G2067), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n732), .A2(G27), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G164), .B2(new_n732), .ZN(new_n816));
  INV_X1    g391(.A(G2078), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n802), .A2(G1961), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n798), .A2(new_n799), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n814), .A2(new_n818), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  AOI211_X1 g396(.A(new_n803), .B(new_n821), .C1(new_n787), .C2(new_n786), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n783), .A2(new_n789), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n770), .A2(G23), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n532), .B1(new_n568), .B2(new_n607), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n610), .A2(new_n611), .ZN(new_n826));
  OAI21_X1  g401(.A(KEYINPUT92), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT92), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n609), .A2(new_n828), .A3(new_n610), .A4(new_n611), .ZN(new_n829));
  AND2_X1   g404(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n824), .B1(new_n830), .B2(new_n770), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT33), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(G1976), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n770), .A2(G6), .ZN(new_n834));
  INV_X1    g409(.A(G305), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n835), .B2(new_n770), .ZN(new_n836));
  XNOR2_X1  g411(.A(KEYINPUT32), .B(G1981), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(KEYINPUT91), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n838), .A2(KEYINPUT91), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n770), .A2(G22), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(G166), .B2(new_n770), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(G1971), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n833), .A2(new_n839), .A3(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT34), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  MUX2_X1   g422(.A(G24), .B(G290), .S(G16), .Z(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(KEYINPUT90), .Z(new_n849));
  AND2_X1   g424(.A1(new_n849), .A2(G1986), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n849), .A2(G1986), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n732), .A2(G25), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n492), .A2(G131), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n497), .A2(G119), .ZN(new_n854));
  OR2_X1    g429(.A1(G95), .A2(G2105), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n855), .B(G2104), .C1(G107), .C2(new_n490), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n852), .B1(new_n858), .B2(new_n732), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT89), .ZN(new_n860));
  XOR2_X1   g435(.A(KEYINPUT35), .B(G1991), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  NOR3_X1   g437(.A1(new_n850), .A2(new_n851), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n847), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(KEYINPUT36), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT36), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n847), .A2(new_n866), .A3(new_n863), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n823), .B1(new_n865), .B2(new_n867), .ZN(G311));
  INV_X1    g443(.A(new_n823), .ZN(new_n869));
  INV_X1    g444(.A(new_n867), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n866), .B1(new_n847), .B2(new_n863), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(G150));
  INV_X1    g447(.A(G67), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n873), .B1(new_n574), .B2(new_n575), .ZN(new_n874));
  AND2_X1   g449(.A1(G80), .A2(G543), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n536), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n557), .A2(G55), .A3(new_n560), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n550), .A2(G93), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(G860), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n880), .B(KEYINPUT37), .Z(new_n881));
  NAND2_X1  g456(.A1(new_n589), .A2(new_n879), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n589), .A2(new_n879), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT38), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n650), .A2(new_n657), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n886), .B(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT39), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT103), .ZN(new_n891));
  INV_X1    g466(.A(G860), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n892), .B1(new_n888), .B2(new_n889), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n881), .B1(new_n891), .B2(new_n893), .ZN(G145));
  NAND2_X1  g469(.A1(new_n761), .A2(new_n741), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n740), .A2(new_n760), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n528), .A2(new_n529), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n812), .B(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n506), .A2(new_n524), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n812), .B(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n902), .A2(new_n895), .A3(new_n896), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n492), .A2(G142), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n497), .A2(G130), .ZN(new_n906));
  NOR2_X1   g481(.A1(G106), .A2(G2105), .ZN(new_n907));
  OAI21_X1  g482(.A(G2104), .B1(new_n490), .B2(G118), .ZN(new_n908));
  OAI211_X1 g483(.A(new_n905), .B(new_n906), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(new_n664), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(new_n857), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n904), .B(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n494), .B(new_n675), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(new_n501), .ZN(new_n915));
  AOI21_X1  g490(.A(G37), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n904), .A2(new_n912), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n911), .B1(new_n900), .B2(new_n903), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(KEYINPUT104), .B1(new_n904), .B2(new_n912), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  XOR2_X1   g497(.A(new_n915), .B(KEYINPUT105), .Z(new_n923));
  OAI21_X1  g498(.A(new_n916), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g500(.A(KEYINPUT109), .ZN(new_n926));
  OR2_X1    g501(.A1(new_n659), .A2(new_n885), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n659), .A2(new_n885), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n646), .A2(new_n792), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n644), .A2(G299), .A3(new_n645), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT41), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n929), .A2(KEYINPUT41), .A3(new_n930), .ZN(new_n934));
  AOI22_X1  g509(.A1(new_n927), .A2(new_n928), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n931), .B(new_n936), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n927), .A2(new_n928), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n935), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  XNOR2_X1  g514(.A(G166), .B(G305), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n827), .A2(new_n829), .ZN(new_n943));
  NOR2_X1   g518(.A1(G290), .A2(new_n943), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n628), .A2(new_n632), .A3(new_n629), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n632), .B1(new_n628), .B2(new_n629), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n830), .B1(new_n947), .B2(new_n627), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n942), .B1(new_n944), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(G290), .A2(new_n943), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n830), .A2(new_n627), .A3(new_n633), .A4(new_n631), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(new_n951), .A3(KEYINPUT107), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n941), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n952), .A2(new_n941), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n953), .A2(KEYINPUT108), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n950), .A2(new_n951), .A3(KEYINPUT107), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT107), .B1(new_n950), .B2(new_n951), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n940), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n952), .A2(new_n941), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n956), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT42), .B1(new_n955), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT42), .B1(new_n959), .B2(new_n960), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n939), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT42), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT108), .B1(new_n953), .B2(new_n954), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n959), .A2(new_n956), .A3(new_n960), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n937), .A2(new_n927), .A3(new_n928), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n933), .A2(new_n934), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n970), .B1(new_n938), .B2(new_n972), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n969), .A2(new_n973), .A3(new_n963), .ZN(new_n974));
  OAI21_X1  g549(.A(G868), .B1(new_n965), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n879), .A2(new_n635), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n926), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n973), .B1(new_n969), .B2(new_n963), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n962), .A2(new_n964), .A3(new_n939), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n635), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n976), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n980), .A2(KEYINPUT109), .A3(new_n981), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n977), .A2(new_n982), .ZN(G295));
  NAND2_X1  g558(.A1(new_n975), .A2(new_n976), .ZN(G331));
  NAND2_X1  g559(.A1(G301), .A2(KEYINPUT110), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT110), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n578), .A2(new_n579), .A3(new_n986), .A4(new_n580), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n985), .B(new_n987), .C1(new_n883), .C2(new_n884), .ZN(new_n988));
  INV_X1    g563(.A(new_n884), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n985), .A2(new_n987), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n989), .A2(new_n990), .A3(new_n882), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n988), .A2(new_n991), .A3(G168), .ZN(new_n992));
  AOI21_X1  g567(.A(G168), .B1(new_n988), .B2(new_n991), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n971), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT111), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n971), .B(KEYINPUT111), .C1(new_n992), .C2(new_n993), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n992), .A2(new_n993), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n931), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n996), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n967), .A2(new_n968), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(G37), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n996), .A2(new_n997), .A3(new_n999), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n1001), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT43), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G37), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(new_n1004), .B2(new_n1001), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT112), .ZN(new_n1009));
  OR2_X1    g584(.A1(new_n994), .A2(new_n1009), .ZN(new_n1010));
  AOI22_X1  g585(.A1(new_n994), .A2(new_n1009), .B1(new_n998), .B2(new_n937), .ZN(new_n1011));
  AOI22_X1  g586(.A1(new_n1010), .A2(new_n1011), .B1(new_n967), .B2(new_n968), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT43), .ZN(new_n1013));
  NOR3_X1   g588(.A1(new_n1008), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT44), .B1(new_n1006), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT44), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1013), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1017));
  NOR3_X1   g592(.A1(new_n1008), .A2(new_n1012), .A3(KEYINPUT43), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1016), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1015), .A2(new_n1019), .ZN(G397));
  OR2_X1    g595(.A1(G290), .A2(G1986), .ZN(new_n1021));
  NAND2_X1  g596(.A1(G290), .A2(G1986), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(KEYINPUT113), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G137), .ZN(new_n1024));
  OAI221_X1 g599(.A(G40), .B1(new_n491), .B2(new_n1024), .C1(new_n485), .C2(new_n486), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1025), .B1(new_n476), .B2(new_n481), .ZN(new_n1026));
  INV_X1    g601(.A(G1384), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n898), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT45), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1026), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1023), .B(new_n1033), .C1(KEYINPUT113), .C2(new_n1022), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n1034), .B(KEYINPUT114), .ZN(new_n1035));
  XNOR2_X1  g610(.A(new_n1032), .B(KEYINPUT115), .ZN(new_n1036));
  OR2_X1    g611(.A1(new_n812), .A2(G2067), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n812), .A2(G2067), .ZN(new_n1038));
  INV_X1    g613(.A(G1996), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1037), .B(new_n1038), .C1(new_n1039), .C2(new_n760), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1032), .A2(G1996), .ZN(new_n1041));
  AOI22_X1  g616(.A1(new_n1036), .A2(new_n1040), .B1(new_n762), .B2(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g617(.A(new_n857), .B(new_n861), .ZN(new_n1043));
  XOR2_X1   g618(.A(new_n1043), .B(KEYINPUT116), .Z(new_n1044));
  NAND2_X1  g619(.A1(new_n1036), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1042), .A2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1035), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G8), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1027), .B1(new_n525), .B2(new_n530), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1030), .B1(new_n1049), .B2(new_n1029), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1025), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n480), .B1(new_n479), .B2(G2105), .ZN(new_n1052));
  AOI211_X1 g627(.A(KEYINPUT67), .B(new_n490), .C1(new_n477), .C2(new_n478), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1051), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n773), .B1(new_n1050), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT50), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1028), .A2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1057), .B1(new_n1049), .B2(new_n1056), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1058), .A2(new_n1026), .A3(new_n787), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1048), .B1(new_n1055), .B2(new_n1059), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1060), .A2(KEYINPUT124), .B1(G8), .B2(G286), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT51), .ZN(new_n1062));
  AOI22_X1  g637(.A1(G286), .A2(G8), .B1(KEYINPUT124), .B2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1064));
  AOI211_X1 g639(.A(new_n1048), .B(G286), .C1(new_n1055), .C2(new_n1059), .ZN(new_n1065));
  OAI22_X1  g640(.A1(new_n1061), .A2(KEYINPUT51), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT62), .ZN(new_n1067));
  NAND2_X1  g642(.A1(G303), .A2(G8), .ZN(new_n1068));
  XOR2_X1   g643(.A(new_n1068), .B(KEYINPUT55), .Z(new_n1069));
  XNOR2_X1  g644(.A(KEYINPUT117), .B(G2090), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1058), .A2(new_n1026), .A3(new_n1070), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n901), .A2(new_n1029), .A3(G1384), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1072), .B1(new_n1049), .B2(new_n1029), .ZN(new_n1073));
  AOI21_X1  g648(.A(G1971), .B1(new_n1073), .B2(new_n1026), .ZN(new_n1074));
  OAI211_X1 g649(.A(G8), .B(new_n1069), .C1(new_n1071), .C2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1028), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1051), .B(new_n1076), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n830), .A2(G1976), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(G8), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT52), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1080), .A2(KEYINPUT118), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1079), .A2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1077), .A2(new_n1078), .A3(G8), .A4(new_n1081), .ZN(new_n1084));
  INV_X1    g659(.A(G1976), .ZN(new_n1085));
  NAND3_X1  g660(.A1(G288), .A2(new_n1080), .A3(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1083), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1077), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1088), .A2(new_n1048), .ZN(new_n1089));
  INV_X1    g664(.A(G1981), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n835), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT49), .ZN(new_n1092));
  NOR2_X1   g667(.A1(G305), .A2(G1981), .ZN(new_n1093));
  OR3_X1    g668(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1092), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1089), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1075), .A2(new_n1087), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1074), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1028), .A2(KEYINPUT50), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n1049), .B2(KEYINPUT50), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1100), .A2(new_n1054), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n1070), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1048), .B1(new_n1098), .B2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(KEYINPUT119), .B1(new_n1103), .B2(new_n1069), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT119), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1069), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1074), .B1(new_n1070), .B2(new_n1101), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1105), .B(new_n1106), .C1(new_n1107), .C2(new_n1048), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1097), .B1(new_n1104), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1073), .A2(new_n1026), .A3(new_n817), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT53), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1058), .A2(new_n1026), .ZN(new_n1112));
  INV_X1    g687(.A(G1961), .ZN(new_n1113));
  AOI22_X1  g688(.A1(new_n1110), .A2(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n817), .A2(KEYINPUT53), .ZN(new_n1115));
  OR3_X1    g690(.A1(new_n1050), .A2(new_n1054), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(G301), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1055), .A2(new_n1059), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1118), .A2(G8), .A3(G168), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1119), .B1(new_n1060), .B2(new_n1063), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT62), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1120), .B(new_n1121), .C1(KEYINPUT51), .C2(new_n1061), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1067), .A2(new_n1109), .A3(new_n1117), .A4(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(G288), .A2(G1976), .ZN(new_n1124));
  AND2_X1   g699(.A1(new_n1096), .A2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1089), .B1(new_n1125), .B2(new_n1093), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n794), .B1(new_n1100), .B2(new_n1054), .ZN(new_n1127));
  NAND2_X1  g702(.A1(KEYINPUT121), .A2(KEYINPUT57), .ZN(new_n1128));
  NAND2_X1  g703(.A1(G299), .A2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(KEYINPUT121), .A2(KEYINPUT57), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NOR3_X1   g706(.A1(G299), .A2(KEYINPUT121), .A3(KEYINPUT57), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g708(.A(KEYINPUT56), .B(G2072), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1073), .A2(new_n1026), .A3(new_n1134), .ZN(new_n1135));
  AND3_X1   g710(.A1(new_n1127), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1127), .A2(new_n1135), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1133), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n646), .ZN(new_n1140));
  AOI21_X1  g715(.A(G1348), .B1(new_n1058), .B2(new_n1026), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1077), .A2(G2067), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1140), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1136), .B1(new_n1139), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1141), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1142), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1145), .A2(new_n1146), .A3(KEYINPUT60), .A4(new_n646), .ZN(new_n1147));
  XOR2_X1   g722(.A(KEYINPUT123), .B(KEYINPUT61), .Z(new_n1148));
  AOI21_X1  g723(.A(new_n1133), .B1(new_n1127), .B2(new_n1135), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1148), .B1(new_n1136), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1145), .A2(new_n1146), .A3(KEYINPUT60), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT60), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1152), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1151), .A2(new_n1153), .A3(new_n1140), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1127), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1139), .A2(KEYINPUT61), .A3(new_n1155), .ZN(new_n1156));
  AND4_X1   g731(.A1(new_n1147), .A2(new_n1150), .A3(new_n1154), .A4(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1073), .A2(new_n1026), .A3(new_n1039), .ZN(new_n1158));
  XOR2_X1   g733(.A(KEYINPUT58), .B(G1341), .Z(new_n1159));
  NAND2_X1  g734(.A1(new_n1077), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(KEYINPUT122), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT122), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1158), .A2(new_n1163), .A3(new_n1160), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(KEYINPUT59), .B1(new_n1165), .B2(new_n590), .ZN(new_n1166));
  AND3_X1   g741(.A1(new_n1158), .A2(new_n1163), .A3(new_n1160), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1163), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1168));
  OAI211_X1 g743(.A(KEYINPUT59), .B(new_n590), .C1(new_n1167), .C2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1166), .A2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1144), .B1(new_n1157), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1031), .A2(new_n1072), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1025), .A2(new_n1115), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1175), .A2(new_n475), .A3(new_n1176), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1173), .A2(new_n1174), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(G171), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1114), .A2(G301), .A3(new_n1116), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1179), .A2(new_n1180), .A3(KEYINPUT54), .ZN(new_n1181));
  XOR2_X1   g756(.A(KEYINPUT125), .B(KEYINPUT54), .Z(new_n1182));
  NOR2_X1   g757(.A1(new_n1178), .A2(G171), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1182), .B1(new_n1183), .B2(new_n1117), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1109), .A2(new_n1181), .A3(new_n1184), .A4(new_n1066), .ZN(new_n1185));
  OAI211_X1 g760(.A(new_n1123), .B(new_n1126), .C1(new_n1172), .C2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1065), .A2(KEYINPUT63), .ZN(new_n1187));
  OAI21_X1  g762(.A(G8), .B1(new_n1071), .B2(new_n1074), .ZN(new_n1188));
  AOI211_X1 g763(.A(new_n1187), .B(new_n1097), .C1(new_n1106), .C2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1119), .B1(new_n1104), .B2(new_n1108), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1075), .ZN(new_n1191));
  OAI211_X1 g766(.A(new_n1096), .B(new_n1087), .C1(new_n1190), .C2(new_n1191), .ZN(new_n1192));
  XOR2_X1   g767(.A(KEYINPUT120), .B(KEYINPUT63), .Z(new_n1193));
  AOI21_X1  g768(.A(new_n1189), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1047), .B1(new_n1186), .B2(new_n1194), .ZN(new_n1195));
  OR2_X1    g770(.A1(new_n1046), .A2(KEYINPUT127), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1046), .A2(KEYINPUT127), .ZN(new_n1197));
  NOR2_X1   g772(.A1(new_n1021), .A2(new_n1032), .ZN(new_n1198));
  XOR2_X1   g773(.A(new_n1198), .B(KEYINPUT48), .Z(new_n1199));
  NAND3_X1  g774(.A1(new_n1196), .A2(new_n1197), .A3(new_n1199), .ZN(new_n1200));
  XOR2_X1   g775(.A(new_n1041), .B(KEYINPUT46), .Z(new_n1201));
  NAND3_X1  g776(.A1(new_n1037), .A2(new_n760), .A3(new_n1038), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1036), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1201), .A2(new_n1203), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n1204), .B(KEYINPUT47), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n858), .A2(new_n861), .ZN(new_n1206));
  XOR2_X1   g781(.A(new_n1206), .B(KEYINPUT126), .Z(new_n1207));
  NAND2_X1  g782(.A1(new_n1042), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1208), .A2(new_n1037), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1209), .A2(new_n1036), .ZN(new_n1210));
  AND3_X1   g785(.A1(new_n1200), .A2(new_n1205), .A3(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1195), .A2(new_n1211), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g787(.A(G319), .ZN(new_n1214));
  NOR4_X1   g788(.A1(G229), .A2(new_n1214), .A3(G401), .A4(G227), .ZN(new_n1215));
  OAI211_X1 g789(.A(new_n924), .B(new_n1215), .C1(new_n1017), .C2(new_n1018), .ZN(G225));
  INV_X1    g790(.A(G225), .ZN(G308));
endmodule


