//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1 0 0 1 0 1 1 1 1 0 0 1 0 1 1 0 1 1 0 1 0 1 1 0 0 1 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 0 0 0 1 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n551, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n614, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1222, new_n1223, new_n1224, new_n1225;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT66), .Z(G173));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  OAI21_X1  g035(.A(KEYINPUT68), .B1(new_n460), .B2(G2105), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n462), .A2(new_n463), .A3(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(G137), .A3(new_n463), .ZN(new_n468));
  INV_X1    g043(.A(G113), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(new_n460), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n470), .B1(new_n467), .B2(G125), .ZN(new_n471));
  OAI211_X1 g046(.A(new_n466), .B(new_n468), .C1(new_n471), .C2(new_n463), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n477), .A2(new_n463), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  NAND4_X1  g060(.A1(new_n474), .A2(new_n476), .A3(G126), .A4(G2105), .ZN(new_n486));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n487), .A2(new_n489), .A3(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n463), .A2(KEYINPUT69), .A3(G138), .ZN(new_n492));
  OAI21_X1  g067(.A(KEYINPUT4), .B1(new_n477), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  AND3_X1   g069(.A1(new_n463), .A2(KEYINPUT69), .A3(G138), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n467), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n491), .B1(new_n493), .B2(new_n496), .ZN(G164));
  INV_X1    g072(.A(G543), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT6), .ZN(new_n499));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n498), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT70), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n503), .A2(new_n504), .A3(G50), .ZN(new_n505));
  INV_X1    g080(.A(new_n502), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  OAI211_X1 g082(.A(G50), .B(G543), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT70), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n512), .B2(G543), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n498), .A2(KEYINPUT71), .A3(KEYINPUT5), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n513), .A2(new_n514), .B1(new_n512), .B2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n501), .A2(new_n502), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n515), .A2(G88), .A3(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  OAI211_X1 g093(.A(new_n510), .B(new_n517), .C1(new_n518), .C2(new_n500), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND3_X1  g095(.A1(new_n515), .A2(G89), .A3(new_n516), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT72), .B(G51), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT7), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n525), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n503), .A2(new_n522), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n513), .A2(new_n514), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n512), .A2(G543), .ZN(new_n529));
  NAND4_X1  g104(.A1(new_n528), .A2(G63), .A3(G651), .A4(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n521), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT73), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n521), .A2(new_n527), .A3(KEYINPUT73), .A4(new_n530), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(G168));
  AOI22_X1  g110(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n500), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n503), .A2(G52), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n515), .A2(new_n516), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n537), .A2(new_n541), .ZN(G171));
  NAND2_X1  g117(.A1(new_n503), .A2(G43), .ZN(new_n543));
  INV_X1    g118(.A(G81), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n539), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n515), .A2(G56), .ZN(new_n546));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n500), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(G188));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n528), .A2(new_n529), .ZN(new_n557));
  INV_X1    g132(.A(G65), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT76), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OAI211_X1 g136(.A(KEYINPUT76), .B(new_n556), .C1(new_n557), .C2(new_n558), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n561), .A2(G651), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n516), .A2(G53), .A3(G543), .ZN(new_n564));
  XNOR2_X1  g139(.A(KEYINPUT74), .B(KEYINPUT9), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT74), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n503), .A2(new_n567), .A3(KEYINPUT9), .A4(G53), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(G91), .ZN(new_n570));
  OAI21_X1  g145(.A(KEYINPUT75), .B1(new_n539), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT75), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n515), .A2(new_n572), .A3(G91), .A4(new_n516), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n569), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n563), .A2(new_n574), .ZN(G299));
  INV_X1    g150(.A(G171), .ZN(G301));
  INV_X1    g151(.A(G168), .ZN(G286));
  NAND3_X1  g152(.A1(new_n515), .A2(G87), .A3(new_n516), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n503), .A2(G49), .ZN(new_n579));
  AND2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(G288));
  NAND3_X1  g157(.A1(new_n528), .A2(G61), .A3(new_n529), .ZN(new_n583));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n500), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n528), .A2(G86), .A3(new_n529), .A4(new_n516), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n503), .A2(G48), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G305));
  NAND2_X1  g165(.A1(new_n503), .A2(G47), .ZN(new_n591));
  INV_X1    g166(.A(G85), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OAI221_X1 g168(.A(new_n591), .B1(new_n539), .B2(new_n592), .C1(new_n593), .C2(new_n500), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n515), .A2(G92), .A3(new_n516), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n557), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G54), .ZN(new_n602));
  INV_X1    g177(.A(new_n503), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT77), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n503), .A2(KEYINPUT77), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n601), .A2(G651), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n598), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n595), .B1(new_n609), .B2(G868), .ZN(G284));
  OAI21_X1  g185(.A(new_n595), .B1(new_n609), .B2(G868), .ZN(G321));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NOR2_X1   g187(.A1(G286), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g188(.A(G299), .B(KEYINPUT78), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(new_n612), .ZN(G297));
  AOI21_X1  g190(.A(new_n613), .B1(new_n614), .B2(new_n612), .ZN(G280));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n609), .B1(new_n617), .B2(G860), .ZN(G148));
  INV_X1    g193(.A(new_n549), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n619), .A2(G868), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n609), .A2(new_n617), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT79), .Z(new_n622));
  AOI21_X1  g197(.A(new_n620), .B1(new_n622), .B2(G868), .ZN(G323));
  XOR2_X1   g198(.A(KEYINPUT80), .B(KEYINPUT11), .Z(new_n624));
  XNOR2_X1  g199(.A(G323), .B(new_n624), .ZN(G282));
  NAND2_X1  g200(.A1(new_n465), .A2(new_n467), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  INV_X1    g203(.A(G2100), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n478), .A2(G135), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n480), .A2(G123), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n463), .A2(G111), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n632), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NAND3_X1  g212(.A1(new_n630), .A2(new_n631), .A3(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2427), .B(G2430), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(KEYINPUT14), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT82), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n644), .A2(KEYINPUT82), .A3(KEYINPUT14), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n642), .A2(new_n643), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2451), .B(G2454), .Z(new_n653));
  XOR2_X1   g228(.A(G2443), .B(G2446), .Z(new_n654));
  XOR2_X1   g229(.A(new_n653), .B(new_n654), .Z(new_n655));
  NAND2_X1  g230(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n657));
  INV_X1    g232(.A(new_n655), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n649), .A2(new_n651), .A3(new_n658), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n656), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n657), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n658), .B1(new_n649), .B2(new_n651), .ZN(new_n662));
  AOI211_X1 g237(.A(new_n650), .B(new_n655), .C1(new_n647), .C2(new_n648), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n640), .B1(new_n660), .B2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT84), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(G14), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n660), .A2(new_n664), .A3(new_n640), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(KEYINPUT83), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT83), .ZN(new_n671));
  NAND4_X1  g246(.A1(new_n660), .A2(new_n664), .A3(new_n671), .A4(new_n640), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n668), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  AND3_X1   g248(.A1(new_n667), .A2(KEYINPUT85), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(KEYINPUT85), .B1(new_n667), .B2(new_n673), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(G401));
  INV_X1    g251(.A(KEYINPUT18), .ZN(new_n677));
  XOR2_X1   g252(.A(G2084), .B(G2090), .Z(new_n678));
  XNOR2_X1  g253(.A(G2067), .B(G2678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(KEYINPUT17), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n678), .A2(new_n679), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n677), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G2072), .B(G2078), .Z(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(new_n680), .B2(KEYINPUT18), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n683), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(G2096), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT86), .B(G2100), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(G227));
  XOR2_X1   g266(.A(G1971), .B(G1976), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT19), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1956), .B(G2474), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1961), .B(G1966), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(KEYINPUT87), .ZN(new_n697));
  OR3_X1    g272(.A1(new_n694), .A2(new_n695), .A3(KEYINPUT87), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n693), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n694), .A2(new_n695), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n696), .A2(new_n702), .ZN(new_n703));
  MUX2_X1   g278(.A(new_n703), .B(new_n702), .S(new_n693), .Z(new_n704));
  NAND2_X1  g279(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT89), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n705), .B(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(G1991), .B(G1996), .Z(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n708), .A2(new_n710), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1981), .B(G1986), .ZN(new_n713));
  AND3_X1   g288(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n713), .B1(new_n711), .B2(new_n712), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n714), .A2(new_n715), .ZN(G229));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n717), .A2(G33), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n478), .A2(G139), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT25), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(G115), .A2(G2104), .ZN(new_n724));
  INV_X1    g299(.A(G127), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n724), .B1(new_n477), .B2(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n723), .B1(G2105), .B2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n718), .B1(new_n728), .B2(G29), .ZN(new_n729));
  INV_X1    g304(.A(G2072), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT98), .Z(new_n732));
  NAND2_X1  g307(.A1(new_n717), .A2(G32), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n480), .A2(G129), .ZN(new_n734));
  NAND3_X1  g309(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT26), .Z(new_n736));
  NAND2_X1  g311(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n478), .A2(G141), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n465), .A2(G105), .ZN(new_n739));
  NOR3_X1   g314(.A1(new_n737), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n733), .B1(new_n740), .B2(new_n717), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT27), .B(G1996), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(G34), .ZN(new_n744));
  AOI21_X1  g319(.A(G29), .B1(new_n744), .B2(KEYINPUT24), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(KEYINPUT24), .B2(new_n744), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n472), .B2(new_n717), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G2084), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n732), .A2(new_n743), .A3(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(G27), .A2(G29), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G164), .B2(G29), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT103), .B(G2078), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n751), .B(new_n752), .Z(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n730), .B2(new_n729), .ZN(new_n754));
  INV_X1    g329(.A(G5), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n755), .A2(G16), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G301), .B2(G16), .ZN(new_n757));
  INV_X1    g332(.A(G1961), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n717), .A2(G35), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G162), .B2(new_n717), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT29), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n754), .B(new_n759), .C1(G2090), .C2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n717), .A2(G26), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT28), .Z(new_n765));
  NOR2_X1   g340(.A1(G104), .A2(G2105), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT96), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n767), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n478), .A2(G140), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n480), .A2(G128), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n771), .A2(KEYINPUT97), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(KEYINPUT97), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n765), .B1(new_n774), .B2(G29), .ZN(new_n775));
  INV_X1    g350(.A(G2067), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NOR3_X1   g352(.A1(new_n749), .A2(new_n763), .A3(new_n777), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n757), .A2(new_n758), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT101), .ZN(new_n780));
  MUX2_X1   g355(.A(G21), .B(G286), .S(G16), .Z(new_n781));
  OR2_X1    g356(.A1(new_n781), .A2(G1966), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT30), .ZN(new_n783));
  AND3_X1   g358(.A1(new_n783), .A2(KEYINPUT100), .A3(G28), .ZN(new_n784));
  AOI21_X1  g359(.A(KEYINPUT100), .B1(new_n783), .B2(G28), .ZN(new_n785));
  OAI221_X1 g360(.A(new_n717), .B1(new_n783), .B2(G28), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT31), .B(G11), .Z(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT99), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n786), .B(new_n788), .C1(new_n636), .C2(new_n717), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n781), .B2(G1966), .ZN(new_n790));
  AND3_X1   g365(.A1(new_n780), .A2(new_n782), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(KEYINPUT102), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT93), .B(G16), .Z(new_n793));
  MUX2_X1   g368(.A(new_n619), .B(G19), .S(new_n793), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT95), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(G1341), .Z(new_n796));
  NOR2_X1   g371(.A1(G4), .A2(G16), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n609), .B2(G16), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT94), .B(G1348), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n778), .A2(new_n792), .A3(new_n796), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n762), .A2(G2090), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT104), .B(G1956), .Z(new_n803));
  NAND2_X1  g378(.A1(new_n793), .A2(G20), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT23), .Z(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G299), .B2(G16), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n802), .B1(new_n803), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(new_n803), .B2(new_n806), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n808), .A2(KEYINPUT105), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(KEYINPUT105), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n809), .B(new_n810), .C1(KEYINPUT102), .C2(new_n791), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n801), .A2(new_n811), .ZN(new_n812));
  MUX2_X1   g387(.A(G23), .B(G288), .S(G16), .Z(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT33), .B(G1976), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(G6), .A2(G16), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(new_n589), .B2(G16), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT32), .B(G1981), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  MUX2_X1   g396(.A(G303), .B(G22), .S(new_n793), .Z(new_n822));
  INV_X1    g397(.A(G1971), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n813), .A2(new_n815), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n818), .A2(new_n819), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n821), .A2(new_n824), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n827), .A2(KEYINPUT34), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n717), .A2(G25), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n478), .A2(G131), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n480), .A2(G119), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n463), .A2(G107), .ZN(new_n832));
  OAI21_X1  g407(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n830), .B(new_n831), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT90), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT91), .Z(new_n836));
  AOI21_X1  g411(.A(new_n829), .B1(new_n836), .B2(G29), .ZN(new_n837));
  XNOR2_X1  g412(.A(KEYINPUT35), .B(G1991), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT92), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n827), .A2(KEYINPUT34), .ZN(new_n842));
  MUX2_X1   g417(.A(G290), .B(G24), .S(new_n793), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(G1986), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(new_n837), .B2(new_n840), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n828), .A2(new_n841), .A3(new_n842), .A4(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT36), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n812), .A2(new_n847), .ZN(G150));
  INV_X1    g423(.A(G150), .ZN(G311));
  AOI22_X1  g424(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT106), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(G651), .B1(new_n850), .B2(new_n851), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n515), .A2(G93), .A3(new_n516), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n503), .A2(G55), .ZN(new_n856));
  AND3_X1   g431(.A1(new_n855), .A2(KEYINPUT107), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(KEYINPUT107), .B1(new_n855), .B2(new_n856), .ZN(new_n858));
  OAI22_X1  g433(.A1(new_n853), .A2(new_n854), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(G860), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(KEYINPUT37), .Z(new_n861));
  NAND3_X1  g436(.A1(new_n859), .A2(KEYINPUT108), .A3(new_n619), .ZN(new_n862));
  INV_X1    g437(.A(new_n545), .ZN(new_n863));
  INV_X1    g438(.A(new_n548), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT108), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n858), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n855), .A2(KEYINPUT107), .A3(new_n856), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(G80), .A2(G543), .ZN(new_n870));
  INV_X1    g445(.A(G67), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n870), .B1(new_n557), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n500), .B1(new_n872), .B2(KEYINPUT106), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(new_n852), .ZN(new_n874));
  OAI21_X1  g449(.A(KEYINPUT108), .B1(new_n545), .B2(new_n548), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n866), .A2(new_n869), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n862), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT38), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n608), .A2(new_n617), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  AND2_X1   g455(.A1(new_n880), .A2(KEYINPUT39), .ZN(new_n881));
  INV_X1    g456(.A(G860), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n882), .B1(new_n880), .B2(KEYINPUT39), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n861), .B1(new_n881), .B2(new_n883), .ZN(G145));
  NAND3_X1  g459(.A1(new_n772), .A2(G164), .A3(new_n773), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(G164), .B1(new_n772), .B2(new_n773), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n740), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n887), .ZN(new_n889));
  INV_X1    g464(.A(new_n740), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(new_n890), .A3(new_n885), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n888), .A2(new_n891), .A3(new_n727), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n727), .B1(new_n888), .B2(new_n891), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n478), .A2(G142), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n480), .A2(G130), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n463), .A2(G118), .ZN(new_n897));
  OAI21_X1  g472(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n895), .B(new_n896), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n627), .B(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(new_n835), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  OAI22_X1  g477(.A1(new_n893), .A2(new_n894), .B1(KEYINPUT109), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n902), .A2(KEYINPUT109), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n888), .A2(new_n891), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(new_n728), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n904), .A2(new_n906), .A3(new_n892), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n636), .B(G160), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(G162), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n903), .A2(new_n907), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n901), .B1(new_n893), .B2(new_n894), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n906), .A2(new_n892), .A3(new_n902), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(new_n909), .A3(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(G37), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n911), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g492(.A(new_n621), .B(KEYINPUT79), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n918), .A2(new_n877), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n877), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n563), .A2(new_n574), .A3(new_n598), .A4(new_n607), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  AOI22_X1  g497(.A1(new_n563), .A2(new_n574), .B1(new_n598), .B2(new_n607), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT41), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(G299), .A2(new_n608), .ZN(new_n926));
  AOI21_X1  g501(.A(KEYINPUT41), .B1(new_n926), .B2(new_n921), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  OR3_X1    g503(.A1(new_n919), .A2(new_n920), .A3(new_n928), .ZN(new_n929));
  OR2_X1    g504(.A1(G166), .A2(G290), .ZN(new_n930));
  NAND2_X1  g505(.A1(G166), .A2(G290), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(G288), .B(new_n589), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(G305), .B(G288), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n935), .A2(new_n930), .A3(new_n931), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT110), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n937), .B1(new_n938), .B2(KEYINPUT42), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n938), .A2(KEYINPUT42), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n939), .B(new_n940), .ZN(new_n941));
  OAI22_X1  g516(.A1(new_n919), .A2(new_n920), .B1(new_n923), .B2(new_n922), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n929), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n941), .B1(new_n929), .B2(new_n942), .ZN(new_n944));
  OAI21_X1  g519(.A(G868), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n859), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n945), .B1(G868), .B2(new_n946), .ZN(G295));
  OAI21_X1  g522(.A(new_n945), .B1(G868), .B2(new_n946), .ZN(G331));
  INV_X1    g523(.A(KEYINPUT112), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n533), .A2(new_n949), .A3(new_n534), .ZN(new_n950));
  NAND2_X1  g525(.A1(G301), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n949), .B1(new_n533), .B2(new_n534), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(G168), .A2(KEYINPUT112), .A3(G171), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n877), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(G168), .A2(KEYINPUT112), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n957), .A2(G301), .A3(new_n950), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n958), .A2(new_n862), .A3(new_n876), .A4(new_n954), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n928), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n922), .A2(new_n923), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n956), .A2(new_n962), .A3(new_n959), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n961), .A2(new_n937), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(new_n915), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n937), .B1(new_n961), .B2(new_n963), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT43), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n961), .A2(new_n963), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n937), .B1(new_n963), .B2(KEYINPUT113), .ZN(new_n969));
  AOI21_X1  g544(.A(G37), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT43), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n961), .B(new_n963), .C1(KEYINPUT113), .C2(new_n937), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n967), .A2(new_n973), .ZN(new_n974));
  XOR2_X1   g549(.A(KEYINPUT111), .B(KEYINPUT44), .Z(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n970), .A2(KEYINPUT115), .A3(new_n972), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT115), .B1(new_n970), .B2(new_n972), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n977), .A2(new_n978), .A3(new_n971), .ZN(new_n979));
  INV_X1    g554(.A(new_n965), .ZN(new_n980));
  INV_X1    g555(.A(new_n937), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n924), .B1(new_n922), .B2(new_n923), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n926), .A2(KEYINPUT41), .A3(new_n921), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n984), .B1(new_n959), .B2(new_n956), .ZN(new_n985));
  INV_X1    g560(.A(new_n963), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n981), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n980), .A2(KEYINPUT114), .A3(new_n971), .A4(new_n987), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n987), .A2(new_n971), .A3(new_n915), .A4(new_n964), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT114), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n988), .A2(new_n991), .A3(KEYINPUT44), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n976), .B1(new_n979), .B2(new_n992), .ZN(G397));
  INV_X1    g568(.A(KEYINPUT116), .ZN(new_n994));
  INV_X1    g569(.A(G40), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n994), .B1(new_n472), .B2(new_n995), .ZN(new_n996));
  AND2_X1   g571(.A1(new_n466), .A2(new_n468), .ZN(new_n997));
  INV_X1    g572(.A(G125), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n477), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(G2105), .B1(new_n999), .B2(new_n470), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n997), .A2(new_n1000), .A3(KEYINPUT116), .A4(G40), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n996), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1003), .B1(G164), .B2(G1384), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n774), .B(G2067), .ZN(new_n1008));
  INV_X1    g583(.A(G1996), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n740), .B(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1007), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n835), .B(new_n840), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1011), .B1(new_n1006), .B2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g588(.A(G290), .B(G1986), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1013), .B1(new_n1007), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n493), .A2(new_n496), .ZN(new_n1016));
  INV_X1    g591(.A(new_n491), .ZN(new_n1017));
  AOI21_X1  g592(.A(G1384), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n996), .A2(new_n1001), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT118), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n580), .A2(new_n1020), .A3(G1976), .A4(new_n581), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n581), .A2(new_n578), .A3(G1976), .A4(new_n579), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT118), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1019), .A2(G8), .A3(new_n1021), .A4(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT52), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT119), .ZN(new_n1026));
  INV_X1    g601(.A(new_n585), .ZN(new_n1027));
  INV_X1    g602(.A(new_n588), .ZN(new_n1028));
  INV_X1    g603(.A(G1981), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(G1981), .B1(new_n585), .B2(new_n588), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1030), .A2(KEYINPUT49), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT120), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT120), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1030), .A2(new_n1031), .A3(new_n1034), .A4(KEYINPUT49), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1019), .A2(G8), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT49), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1024), .ZN(new_n1041));
  INV_X1    g616(.A(G1976), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT52), .B1(G288), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT119), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1024), .A2(new_n1045), .A3(KEYINPUT52), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1026), .A2(new_n1040), .A3(new_n1044), .A4(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1050));
  OR2_X1    g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT50), .ZN(new_n1052));
  INV_X1    g627(.A(G1384), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n477), .A2(KEYINPUT4), .A3(new_n492), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n494), .B1(new_n467), .B2(new_n495), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1052), .B(new_n1053), .C1(new_n1056), .C2(new_n491), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT117), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1018), .A2(new_n1059), .A3(new_n1052), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1062), .A2(new_n996), .A3(new_n1001), .ZN(new_n1063));
  NOR3_X1   g638(.A1(new_n1061), .A2(G2090), .A3(new_n1063), .ZN(new_n1064));
  OAI211_X1 g639(.A(KEYINPUT45), .B(new_n1053), .C1(new_n1056), .C2(new_n491), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n1004), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(G1971), .B1(new_n1066), .B2(new_n1002), .ZN(new_n1067));
  OAI211_X1 g642(.A(G8), .B(new_n1051), .C1(new_n1064), .C2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(G288), .A2(G1976), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1040), .A2(new_n1069), .B1(new_n1029), .B2(new_n589), .ZN(new_n1070));
  OAI22_X1  g645(.A1(new_n1047), .A2(new_n1068), .B1(new_n1070), .B2(new_n1037), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT121), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1059), .B1(new_n1018), .B2(new_n1052), .ZN(new_n1073));
  NOR4_X1   g648(.A1(G164), .A2(KEYINPUT117), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(G2090), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1062), .A2(new_n996), .A3(new_n1001), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1004), .A2(new_n996), .A3(new_n1065), .A4(new_n1001), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n823), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1051), .B1(new_n1081), .B2(G8), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1072), .B1(new_n1047), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(G8), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AOI22_X1  g661(.A1(new_n1036), .A2(new_n1039), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1024), .A2(new_n1045), .A3(KEYINPUT52), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1045), .B1(new_n1024), .B2(KEYINPUT52), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1086), .A2(KEYINPUT121), .A3(new_n1087), .A4(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(G8), .ZN(new_n1092));
  INV_X1    g667(.A(G2084), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1075), .A2(new_n1093), .A3(new_n1077), .ZN(new_n1094));
  INV_X1    g669(.A(G1966), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1079), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1092), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  AND4_X1   g672(.A1(KEYINPUT63), .A2(new_n1068), .A3(G168), .A4(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1083), .A2(new_n1091), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT63), .ZN(new_n1100));
  AND4_X1   g675(.A1(new_n996), .A2(new_n1062), .A3(new_n1001), .A4(new_n1057), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1101), .A2(new_n1076), .B1(new_n823), .B2(new_n1079), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1085), .B1(new_n1102), .B2(new_n1092), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1090), .A2(new_n1087), .A3(new_n1103), .A4(new_n1068), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1097), .A2(G168), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1100), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1071), .B1(new_n1099), .B2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n758), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1108));
  INV_X1    g683(.A(G2078), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1066), .A2(new_n1002), .A3(KEYINPUT53), .A4(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT53), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1111), .B1(new_n1079), .B2(G2078), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1108), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(G171), .ZN(new_n1114));
  NOR4_X1   g689(.A1(new_n472), .A2(new_n1111), .A3(new_n995), .A4(G2078), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1066), .A2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1108), .A2(new_n1112), .A3(new_n1116), .A4(G301), .ZN(new_n1117));
  AOI21_X1  g692(.A(KEYINPUT54), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1108), .A2(new_n1112), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1119), .A2(KEYINPUT127), .A3(G301), .A4(new_n1110), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT127), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1121), .B1(new_n1113), .B2(G171), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT54), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1108), .A2(new_n1112), .A3(new_n1116), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1124), .B1(new_n1125), .B2(G171), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1118), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1061), .A2(G2084), .A3(new_n1063), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1096), .ZN(new_n1129));
  OAI211_X1 g704(.A(G8), .B(G286), .C1(new_n1128), .C2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT124), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT124), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1097), .A2(new_n1132), .A3(G286), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1094), .A2(G168), .A3(new_n1096), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT125), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT51), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .A4(G8), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1135), .A2(G8), .ZN(new_n1139));
  NAND2_X1  g714(.A1(KEYINPUT125), .A2(KEYINPUT51), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1134), .A2(new_n1138), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT126), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1103), .A2(new_n1068), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1144), .B1(new_n1145), .B2(new_n1047), .ZN(new_n1146));
  AND2_X1   g721(.A1(new_n1103), .A2(new_n1068), .ZN(new_n1147));
  AND4_X1   g722(.A1(new_n1040), .A2(new_n1026), .A3(new_n1044), .A4(new_n1046), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1147), .A2(new_n1148), .A3(KEYINPUT126), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1127), .A2(new_n1143), .A3(new_n1146), .A4(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1079), .ZN(new_n1151));
  XNOR2_X1  g726(.A(KEYINPUT56), .B(G2072), .ZN(new_n1152));
  INV_X1    g727(.A(G1956), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1062), .A2(new_n996), .A3(new_n1057), .A4(new_n1001), .ZN(new_n1154));
  AOI22_X1  g729(.A1(new_n1151), .A2(new_n1152), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT57), .ZN(new_n1156));
  AND3_X1   g731(.A1(new_n563), .A2(new_n574), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1156), .B1(new_n563), .B2(new_n574), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(KEYINPUT122), .B1(new_n1155), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1158), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n563), .A2(new_n574), .A3(new_n1156), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT122), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1154), .A2(new_n1153), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1152), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1079), .A2(new_n1167), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1163), .B(new_n1164), .C1(new_n1166), .C2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(G1348), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1019), .A2(G2067), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n609), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1160), .A2(new_n1169), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1174), .A2(new_n1159), .A3(new_n1165), .ZN(new_n1175));
  AND2_X1   g750(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  XOR2_X1   g751(.A(KEYINPUT123), .B(G1996), .Z(new_n1177));
  NOR2_X1   g752(.A1(new_n1079), .A2(new_n1177), .ZN(new_n1178));
  XOR2_X1   g753(.A(KEYINPUT58), .B(G1341), .Z(new_n1179));
  AND2_X1   g754(.A1(new_n1019), .A2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n549), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT59), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1171), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n608), .A2(KEYINPUT60), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1186));
  OAI211_X1 g761(.A(new_n1184), .B(new_n1185), .C1(new_n1186), .C2(G1348), .ZN(new_n1187));
  OAI211_X1 g762(.A(KEYINPUT59), .B(new_n549), .C1(new_n1178), .C2(new_n1180), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1183), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT60), .ZN(new_n1190));
  OAI211_X1 g765(.A(new_n608), .B(new_n1184), .C1(new_n1186), .C2(G1348), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1190), .B1(new_n1172), .B2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1163), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1193));
  AOI21_X1  g768(.A(KEYINPUT61), .B1(new_n1193), .B2(new_n1175), .ZN(new_n1194));
  NOR3_X1   g769(.A1(new_n1189), .A2(new_n1192), .A3(new_n1194), .ZN(new_n1195));
  NAND4_X1  g770(.A1(new_n1160), .A2(new_n1169), .A3(KEYINPUT61), .A4(new_n1175), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1176), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1107), .B1(new_n1150), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT62), .ZN(new_n1199));
  AND2_X1   g774(.A1(new_n1142), .A2(new_n1138), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1199), .B1(new_n1200), .B2(new_n1134), .ZN(new_n1201));
  AND4_X1   g776(.A1(new_n1199), .A2(new_n1134), .A3(new_n1138), .A4(new_n1142), .ZN(new_n1202));
  INV_X1    g777(.A(new_n1114), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1149), .A2(new_n1146), .A3(new_n1203), .ZN(new_n1204));
  NOR3_X1   g779(.A1(new_n1201), .A2(new_n1202), .A3(new_n1204), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1015), .B1(new_n1198), .B2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1007), .B1(new_n1008), .B2(new_n890), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT46), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1208), .B1(new_n1006), .B2(G1996), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1007), .A2(KEYINPUT46), .A3(new_n1009), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1207), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  XOR2_X1   g786(.A(new_n1211), .B(KEYINPUT47), .Z(new_n1212));
  NOR2_X1   g787(.A1(new_n774), .A2(G2067), .ZN(new_n1213));
  NOR2_X1   g788(.A1(new_n836), .A2(new_n839), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1213), .B1(new_n1214), .B2(new_n1011), .ZN(new_n1215));
  NOR3_X1   g790(.A1(new_n1006), .A2(G1986), .A3(G290), .ZN(new_n1216));
  XNOR2_X1  g791(.A(new_n1216), .B(KEYINPUT48), .ZN(new_n1217));
  OAI22_X1  g792(.A1(new_n1215), .A2(new_n1006), .B1(new_n1013), .B2(new_n1217), .ZN(new_n1218));
  NOR2_X1   g793(.A1(new_n1212), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1206), .A2(new_n1219), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g795(.A(G319), .B1(new_n689), .B2(new_n690), .ZN(new_n1222));
  NOR3_X1   g796(.A1(new_n714), .A2(new_n715), .A3(new_n1222), .ZN(new_n1223));
  OAI211_X1 g797(.A(new_n1223), .B(new_n916), .C1(new_n674), .C2(new_n675), .ZN(new_n1224));
  INV_X1    g798(.A(new_n974), .ZN(new_n1225));
  NOR2_X1   g799(.A1(new_n1224), .A2(new_n1225), .ZN(G308));
  OR2_X1    g800(.A1(new_n1224), .A2(new_n1225), .ZN(G225));
endmodule


