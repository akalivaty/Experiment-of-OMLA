//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 1 0 0 0 1 0 0 0 0 1 0 0 0 1 0 1 0 1 0 0 0 1 1 0 0 0 1 0 1 1 0 0 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 1 1 0 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n761, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n871, new_n872, new_n873, new_n874, new_n876, new_n877, new_n878,
    new_n879, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962, new_n963;
  INV_X1    g000(.A(KEYINPUT70), .ZN(new_n202));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT24), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  NOR2_X1   g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  OR2_X1    g007(.A1(new_n208), .A2(KEYINPUT23), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(KEYINPUT23), .ZN(new_n210));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n207), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n210), .A2(new_n211), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n214), .B(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G183gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n217), .A2(G190gat), .ZN(new_n218));
  OAI211_X1 g017(.A(KEYINPUT25), .B(new_n209), .C1(new_n218), .C2(new_n205), .ZN(new_n219));
  OAI22_X1  g018(.A1(new_n213), .A2(KEYINPUT25), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(KEYINPUT27), .B(G183gat), .ZN(new_n221));
  INV_X1    g020(.A(G190gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT28), .ZN(new_n224));
  AND2_X1   g023(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT27), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  OR2_X1    g026(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n228));
  AND2_X1   g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT28), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(new_n222), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n224), .B(KEYINPUT66), .C1(new_n229), .C2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n231), .B1(new_n227), .B2(new_n228), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n230), .B1(new_n221), .B2(new_n222), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n208), .A2(KEYINPUT26), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(new_n203), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n208), .A2(KEYINPUT26), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n238), .B1(new_n211), .B2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n232), .A2(new_n236), .A3(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G113gat), .B(G120gat), .ZN(new_n242));
  OR2_X1    g041(.A1(new_n242), .A2(KEYINPUT69), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(KEYINPUT69), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT1), .ZN(new_n245));
  INV_X1    g044(.A(G127gat), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n245), .B1(new_n246), .B2(G134gat), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n247), .B1(new_n246), .B2(G134gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n243), .A2(new_n244), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n246), .A2(KEYINPUT68), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT68), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(G127gat), .ZN(new_n252));
  AND3_X1   g051(.A1(new_n250), .A2(new_n252), .A3(G134gat), .ZN(new_n253));
  OAI21_X1  g052(.A(KEYINPUT67), .B1(new_n246), .B2(G134gat), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n255));
  INV_X1    g054(.A(G134gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(new_n256), .A3(G127gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  OAI22_X1  g057(.A1(new_n253), .A2(new_n258), .B1(KEYINPUT1), .B2(new_n242), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n249), .A2(new_n259), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n220), .A2(new_n241), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n260), .B1(new_n220), .B2(new_n241), .ZN(new_n262));
  NAND2_X1  g061(.A1(G227gat), .A2(G233gat), .ZN(new_n263));
  NOR3_X1   g062(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT32), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n202), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n220), .A2(new_n241), .ZN(new_n267));
  AND2_X1   g066(.A1(new_n249), .A2(new_n259), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n263), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n220), .A2(new_n241), .A3(new_n260), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n272), .A2(KEYINPUT70), .A3(KEYINPUT32), .ZN(new_n273));
  XNOR2_X1  g072(.A(G15gat), .B(G43gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(G71gat), .B(G99gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT33), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n276), .B1(new_n272), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n266), .A2(new_n273), .A3(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n266), .A2(new_n278), .A3(KEYINPUT71), .A4(new_n273), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n264), .A2(new_n265), .ZN(new_n284));
  OR2_X1    g083(.A1(new_n276), .A2(new_n277), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n269), .A2(new_n271), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(new_n263), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT34), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT34), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n288), .A2(new_n291), .A3(new_n263), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n287), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n293), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n283), .A2(new_n286), .A3(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT31), .B(G50gat), .ZN(new_n297));
  INV_X1    g096(.A(G106gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(G78gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(KEYINPUT75), .B(G155gat), .ZN(new_n301));
  INV_X1    g100(.A(G162gat), .ZN(new_n302));
  OAI21_X1  g101(.A(KEYINPUT2), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  XOR2_X1   g102(.A(G141gat), .B(G148gat), .Z(new_n304));
  XNOR2_X1  g103(.A(G155gat), .B(G162gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT2), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n305), .B1(new_n304), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G197gat), .B(G204gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT22), .ZN(new_n312));
  INV_X1    g111(.A(G211gat), .ZN(new_n313));
  INV_X1    g112(.A(G218gat), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G211gat), .B(G218gat), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n317), .A2(new_n311), .A3(new_n315), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT29), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT81), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT3), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n325), .B1(new_n321), .B2(new_n322), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n310), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n319), .A2(new_n320), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n306), .A2(new_n309), .A3(new_n325), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT29), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n327), .A2(new_n332), .ZN(new_n333));
  AND2_X1   g132(.A1(G228gat), .A2(G233gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n334), .B(KEYINPUT80), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(G22gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n310), .A2(new_n321), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n310), .A2(KEYINPUT3), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n338), .A2(new_n339), .A3(new_n334), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n340), .A2(new_n331), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n336), .A2(new_n337), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n335), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n344), .B1(new_n327), .B2(new_n332), .ZN(new_n345));
  OAI21_X1  g144(.A(G22gat), .B1(new_n345), .B2(new_n341), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n300), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n343), .A2(new_n346), .A3(new_n300), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n299), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n349), .ZN(new_n351));
  INV_X1    g150(.A(new_n299), .ZN(new_n352));
  NOR3_X1   g151(.A1(new_n351), .A2(new_n347), .A3(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n294), .A2(new_n296), .A3(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(G8gat), .B(G36gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(G64gat), .B(G92gat), .ZN(new_n358));
  XOR2_X1   g157(.A(new_n357), .B(new_n358), .Z(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n328), .ZN(new_n361));
  INV_X1    g160(.A(G226gat), .ZN(new_n362));
  INV_X1    g161(.A(G233gat), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n364), .B1(new_n267), .B2(new_n330), .ZN(new_n365));
  INV_X1    g164(.A(new_n364), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n366), .B1(new_n220), .B2(new_n241), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n361), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n267), .A2(new_n364), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT29), .B1(new_n220), .B2(new_n241), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n369), .B(new_n328), .C1(new_n364), .C2(new_n370), .ZN(new_n371));
  AND3_X1   g170(.A1(new_n368), .A2(KEYINPUT72), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT72), .B1(new_n368), .B2(new_n371), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n360), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n368), .A2(KEYINPUT30), .A3(new_n371), .A4(new_n359), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n368), .A2(new_n371), .A3(new_n359), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT74), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT73), .B(KEYINPUT30), .ZN(new_n378));
  AND3_X1   g177(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n377), .B1(new_n376), .B2(new_n378), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n374), .B(new_n375), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(G1gat), .B(G29gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(KEYINPUT0), .ZN(new_n383));
  XNOR2_X1  g182(.A(G57gat), .B(G85gat), .ZN(new_n384));
  XOR2_X1   g183(.A(new_n383), .B(new_n384), .Z(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G225gat), .A2(G233gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(KEYINPUT76), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n249), .A2(new_n306), .A3(new_n309), .A4(new_n259), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  AOI22_X1  g189(.A1(new_n259), .A2(new_n249), .B1(new_n306), .B2(new_n309), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n388), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT78), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(new_n393), .A3(KEYINPUT5), .ZN(new_n394));
  INV_X1    g193(.A(new_n388), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n260), .A2(new_n310), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n395), .B1(new_n396), .B2(new_n389), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT5), .ZN(new_n398));
  OAI21_X1  g197(.A(KEYINPUT78), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n306), .A2(new_n309), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n268), .A2(new_n400), .A3(KEYINPUT4), .ZN(new_n401));
  XNOR2_X1  g200(.A(KEYINPUT77), .B(KEYINPUT4), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n389), .A2(new_n402), .ZN(new_n403));
  AND3_X1   g202(.A1(new_n401), .A2(new_n403), .A3(new_n395), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n339), .A2(new_n329), .A3(new_n260), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n394), .A2(new_n399), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OR2_X1    g205(.A1(new_n389), .A2(new_n402), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n407), .B(new_n405), .C1(KEYINPUT4), .C2(new_n390), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n395), .A2(new_n398), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n386), .B1(new_n406), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT6), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NOR3_X1   g213(.A1(new_n406), .A2(new_n386), .A3(new_n410), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n411), .B1(new_n415), .B2(KEYINPUT6), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NOR3_X1   g216(.A1(new_n381), .A2(new_n417), .A3(KEYINPUT35), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n356), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT79), .B1(new_n415), .B2(KEYINPUT6), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n394), .A2(new_n399), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n405), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n410), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n423), .A2(new_n424), .A3(new_n385), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT79), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n425), .A2(new_n426), .A3(new_n413), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n420), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n411), .ZN(new_n429));
  INV_X1    g228(.A(new_n381), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n429), .A2(new_n430), .A3(new_n414), .ZN(new_n431));
  OAI211_X1 g230(.A(KEYINPUT84), .B(KEYINPUT35), .C1(new_n355), .C2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n295), .B1(new_n283), .B2(new_n286), .ZN(new_n434));
  INV_X1    g233(.A(new_n286), .ZN(new_n435));
  AOI211_X1 g234(.A(new_n293), .B(new_n435), .C1(new_n281), .C2(new_n282), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n412), .B1(new_n420), .B2(new_n427), .ZN(new_n438));
  INV_X1    g237(.A(new_n414), .ZN(new_n439));
  NOR3_X1   g238(.A1(new_n438), .A2(new_n381), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n437), .A2(new_n440), .A3(new_n354), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT84), .B1(new_n441), .B2(KEYINPUT35), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n419), .B1(new_n433), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n294), .A2(KEYINPUT36), .A3(new_n296), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT36), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n445), .B1(new_n434), .B2(new_n436), .ZN(new_n446));
  INV_X1    g245(.A(new_n354), .ZN(new_n447));
  AOI22_X1  g246(.A1(new_n444), .A2(new_n446), .B1(new_n431), .B2(new_n447), .ZN(new_n448));
  AND2_X1   g247(.A1(new_n448), .A2(KEYINPUT82), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT37), .ZN(new_n450));
  INV_X1    g249(.A(new_n373), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n368), .A2(KEYINPUT72), .A3(new_n371), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  XOR2_X1   g252(.A(KEYINPUT83), .B(KEYINPUT37), .Z(new_n454));
  NAND3_X1  g253(.A1(new_n368), .A2(new_n371), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n360), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT38), .B1(new_n453), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n450), .B1(new_n368), .B2(new_n371), .ZN(new_n458));
  OR3_X1    g257(.A1(new_n456), .A2(KEYINPUT38), .A3(new_n458), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n457), .A2(new_n417), .A3(new_n376), .A4(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n408), .A2(new_n388), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n385), .B1(new_n461), .B2(KEYINPUT39), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n396), .A2(new_n389), .A3(new_n395), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n463), .A2(KEYINPUT39), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n462), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n412), .B1(new_n465), .B2(KEYINPUT40), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n381), .B(new_n466), .C1(KEYINPUT40), .C2(new_n465), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n460), .A2(new_n467), .A3(new_n354), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n468), .B1(new_n448), .B2(KEYINPUT82), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n443), .B1(new_n449), .B2(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(G169gat), .B(G197gat), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n471), .B(KEYINPUT86), .ZN(new_n472));
  INV_X1    g271(.A(G113gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n472), .B(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n475));
  INV_X1    g274(.A(G141gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n475), .B(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n474), .B(new_n477), .ZN(new_n478));
  XOR2_X1   g277(.A(KEYINPUT87), .B(KEYINPUT12), .Z(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  OR2_X1    g280(.A1(new_n474), .A2(new_n477), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n474), .A2(new_n477), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n482), .A2(new_n479), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(G15gat), .B(G22gat), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n487), .A2(G1gat), .ZN(new_n488));
  OAI21_X1  g287(.A(G8gat), .B1(new_n488), .B2(KEYINPUT91), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT16), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n487), .B1(new_n490), .B2(G1gat), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n491), .B1(G1gat), .B2(new_n487), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n489), .B(new_n492), .ZN(new_n493));
  AND2_X1   g292(.A1(G43gat), .A2(G50gat), .ZN(new_n494));
  NOR2_X1   g293(.A1(G43gat), .A2(G50gat), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT15), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(G29gat), .ZN(new_n498));
  INV_X1    g297(.A(G36gat), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n502));
  NOR3_X1   g301(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT88), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT14), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n506), .A2(new_n498), .A3(new_n499), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n507), .A2(KEYINPUT88), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n501), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(G43gat), .ZN(new_n510));
  INV_X1    g309(.A(G50gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT15), .ZN(new_n513));
  NAND2_X1  g312(.A1(G43gat), .A2(G50gat), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n496), .A2(new_n515), .A3(new_n501), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT89), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n507), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT89), .B1(new_n519), .B2(new_n499), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n502), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  AOI22_X1  g320(.A1(new_n497), .A2(new_n509), .B1(new_n516), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n493), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n498), .A2(new_n499), .ZN(new_n524));
  AOI22_X1  g323(.A1(new_n507), .A2(KEYINPUT88), .B1(new_n524), .B2(KEYINPUT14), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n503), .A2(new_n504), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n500), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n507), .A2(new_n517), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n503), .A2(KEYINPUT89), .ZN(new_n529));
  AOI22_X1  g328(.A1(new_n528), .A2(new_n529), .B1(KEYINPUT14), .B2(new_n524), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n496), .A2(new_n515), .A3(new_n501), .ZN(new_n531));
  OAI22_X1  g330(.A1(new_n527), .A2(new_n496), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT17), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT90), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n535), .B1(new_n522), .B2(KEYINPUT17), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n532), .A2(KEYINPUT90), .A3(new_n533), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n523), .B1(new_n538), .B2(new_n493), .ZN(new_n539));
  NAND2_X1  g338(.A1(G229gat), .A2(G233gat), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT18), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n522), .A2(KEYINPUT17), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n509), .A2(new_n497), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n516), .A2(new_n521), .ZN(new_n544));
  AOI211_X1 g343(.A(new_n535), .B(KEYINPUT17), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT90), .B1(new_n532), .B2(new_n533), .ZN(new_n546));
  OAI211_X1 g345(.A(new_n493), .B(new_n542), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(new_n489), .B(new_n492), .Z(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(new_n532), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n547), .A2(KEYINPUT18), .A3(new_n540), .A4(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n493), .A2(new_n522), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(new_n540), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n486), .B1(new_n541), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n547), .A2(new_n540), .A3(new_n549), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT18), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n561), .A2(new_n485), .A3(new_n550), .A4(new_n556), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  AND2_X1   g362(.A1(new_n470), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT93), .B1(G71gat), .B2(G78gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(G71gat), .A2(G78gat), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT94), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT9), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  OR2_X1    g368(.A1(G57gat), .A2(G64gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(G57gat), .A2(G64gat), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n567), .B1(new_n566), .B2(new_n568), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n565), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(G71gat), .B(G78gat), .Z(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n575), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n577), .B(new_n565), .C1(new_n572), .C2(new_n573), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT95), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n576), .A2(KEYINPUT95), .A3(new_n578), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n548), .B1(new_n583), .B2(KEYINPUT21), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT96), .ZN(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(G155gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n585), .B(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n579), .A2(KEYINPUT21), .ZN(new_n589));
  AND2_X1   g388(.A1(G231gat), .A2(G233gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(new_n246), .ZN(new_n592));
  XOR2_X1   g391(.A(G183gat), .B(G211gat), .Z(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n591), .B(G127gat), .ZN(new_n595));
  INV_X1    g394(.A(new_n593), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n588), .B(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(G85gat), .A2(G92gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT7), .ZN(new_n601));
  NAND2_X1  g400(.A1(G99gat), .A2(G106gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT8), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT97), .ZN(new_n604));
  OR2_X1    g403(.A1(G85gat), .A2(G92gat), .ZN(new_n605));
  AND3_X1   g404(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n604), .B1(new_n603), .B2(new_n605), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n601), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(G99gat), .B(G106gat), .Z(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n609), .ZN(new_n611));
  OAI211_X1 g410(.A(new_n611), .B(new_n601), .C1(new_n606), .C2(new_n607), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n542), .B(new_n613), .C1(new_n545), .C2(new_n546), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n610), .A2(new_n612), .ZN(new_n615));
  AND2_X1   g414(.A1(G232gat), .A2(G233gat), .ZN(new_n616));
  AOI22_X1  g415(.A1(new_n615), .A2(new_n532), .B1(KEYINPUT41), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(G190gat), .B(G218gat), .Z(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n616), .A2(KEYINPUT41), .ZN(new_n621));
  XNOR2_X1  g420(.A(G134gat), .B(G162gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n619), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n614), .A2(new_n624), .A3(new_n617), .ZN(new_n625));
  AND3_X1   g424(.A1(new_n620), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n623), .B1(new_n620), .B2(new_n625), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n599), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(KEYINPUT98), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT98), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n599), .A2(new_n632), .A3(new_n629), .ZN(new_n633));
  INV_X1    g432(.A(G230gat), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n634), .A2(new_n363), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT99), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n612), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n579), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n615), .ZN(new_n640));
  AOI22_X1  g439(.A1(new_n576), .A2(new_n578), .B1(new_n612), .B2(new_n637), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(new_n613), .ZN(new_n642));
  AOI21_X1  g441(.A(KEYINPUT10), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT10), .ZN(new_n644));
  AOI211_X1 g443(.A(new_n644), .B(new_n613), .C1(new_n581), .C2(new_n582), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n636), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n640), .A2(new_n635), .A3(new_n642), .ZN(new_n647));
  XNOR2_X1  g446(.A(G120gat), .B(G148gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(G176gat), .B(G204gat), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n648), .B(new_n649), .Z(new_n650));
  NAND3_X1  g449(.A1(new_n646), .A2(new_n647), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n650), .B1(new_n646), .B2(new_n647), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n631), .A2(new_n633), .A3(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n564), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n438), .A2(new_n439), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g461(.A1(new_n657), .A2(new_n430), .ZN(new_n663));
  XOR2_X1   g462(.A(KEYINPUT16), .B(G8gat), .Z(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(G8gat), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n665), .B1(new_n666), .B2(new_n663), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(KEYINPUT42), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT42), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n668), .A2(new_n670), .ZN(G1325gat));
  INV_X1    g470(.A(KEYINPUT101), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n444), .A2(new_n446), .A3(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n672), .B1(new_n444), .B2(new_n446), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n658), .A2(G15gat), .A3(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n564), .A2(new_n437), .A3(new_n656), .ZN(new_n679));
  INV_X1    g478(.A(G15gat), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n679), .A2(KEYINPUT100), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(KEYINPUT100), .B1(new_n679), .B2(new_n680), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n678), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(KEYINPUT102), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT102), .ZN(new_n685));
  OAI211_X1 g484(.A(new_n678), .B(new_n685), .C1(new_n681), .C2(new_n682), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(G1326gat));
  NOR2_X1   g486(.A1(new_n657), .A2(new_n354), .ZN(new_n688));
  XOR2_X1   g487(.A(KEYINPUT43), .B(G22gat), .Z(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1327gat));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n691));
  OAI21_X1  g490(.A(KEYINPUT35), .B1(new_n355), .B2(new_n431), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT84), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI22_X1  g493(.A1(new_n694), .A2(new_n432), .B1(new_n356), .B2(new_n418), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n431), .A2(new_n447), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(new_n468), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n674), .A2(new_n697), .A3(new_n675), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n628), .B1(new_n695), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n629), .A2(new_n691), .ZN(new_n700));
  AOI22_X1  g499(.A1(new_n691), .A2(new_n699), .B1(new_n470), .B2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n599), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(new_n654), .ZN(new_n703));
  INV_X1    g502(.A(new_n563), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(G29gat), .B1(new_n706), .B2(new_n659), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n703), .A2(new_n629), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n470), .A2(new_n563), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n660), .A2(new_n498), .ZN(new_n710));
  OR3_X1    g509(.A1(new_n709), .A2(KEYINPUT103), .A3(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT45), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT103), .B1(new_n709), .B2(new_n710), .ZN(new_n713));
  AND3_X1   g512(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n712), .B1(new_n711), .B2(new_n713), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n707), .B1(new_n714), .B2(new_n715), .ZN(G1328gat));
  OAI21_X1  g515(.A(G36gat), .B1(new_n706), .B2(new_n430), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n564), .A2(new_n499), .A3(new_n381), .A4(new_n708), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT46), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n718), .A2(KEYINPUT46), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n720), .A2(KEYINPUT104), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n720), .A2(KEYINPUT104), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n717), .B(new_n719), .C1(new_n721), .C2(new_n722), .ZN(G1329gat));
  INV_X1    g522(.A(KEYINPUT106), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n724), .A2(KEYINPUT47), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n437), .A2(new_n510), .ZN(new_n726));
  OR3_X1    g525(.A1(new_n709), .A2(KEYINPUT105), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(KEYINPUT105), .B1(new_n709), .B2(new_n726), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n725), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(G43gat), .B1(new_n706), .B2(new_n676), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n724), .A2(KEYINPUT47), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n732), .B(KEYINPUT107), .Z(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n729), .A2(new_n730), .A3(new_n733), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(G1330gat));
  OAI21_X1  g536(.A(G50gat), .B1(new_n706), .B2(new_n354), .ZN(new_n738));
  OR2_X1    g537(.A1(new_n709), .A2(KEYINPUT108), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n709), .A2(KEYINPUT108), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n739), .A2(new_n511), .A3(new_n447), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT48), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(G1331gat));
  INV_X1    g543(.A(new_n654), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n631), .A2(new_n704), .A3(new_n633), .A4(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n675), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n747), .A2(new_n696), .A3(new_n468), .A4(new_n673), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n746), .B1(new_n443), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(new_n660), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n381), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n752), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n753));
  XOR2_X1   g552(.A(KEYINPUT49), .B(G64gat), .Z(new_n754));
  OAI21_X1  g553(.A(new_n753), .B1(new_n752), .B2(new_n754), .ZN(G1333gat));
  NAND2_X1  g554(.A1(new_n749), .A2(new_n677), .ZN(new_n756));
  INV_X1    g555(.A(new_n437), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(G71gat), .ZN(new_n758));
  AOI22_X1  g557(.A1(new_n756), .A2(G71gat), .B1(new_n749), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g559(.A1(new_n749), .A2(new_n447), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g561(.A1(new_n699), .A2(new_n691), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n449), .A2(new_n469), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n700), .B1(new_n764), .B2(new_n695), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n599), .A2(new_n563), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n767), .A2(new_n654), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n763), .A2(new_n660), .A3(new_n765), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(KEYINPUT109), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT109), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n701), .A2(new_n771), .A3(new_n660), .A4(new_n768), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n770), .A2(new_n772), .A3(G85gat), .ZN(new_n773));
  NAND2_X1  g572(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT111), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT51), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  OAI211_X1 g576(.A(KEYINPUT110), .B(new_n628), .C1(new_n695), .C2(new_n698), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n766), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n443), .A2(new_n748), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT110), .B1(new_n780), .B2(new_n628), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n774), .B(new_n777), .C1(new_n779), .C2(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n629), .B1(new_n443), .B2(new_n748), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n767), .B1(new_n783), .B2(KEYINPUT110), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT110), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n699), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n784), .A2(new_n775), .A3(new_n776), .A4(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n659), .A2(G85gat), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n782), .A2(new_n787), .A3(new_n745), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT112), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n773), .A2(new_n789), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(G1336gat));
  AND2_X1   g593(.A1(new_n782), .A2(new_n787), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n430), .A2(G92gat), .A3(new_n654), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n701), .A2(new_n768), .ZN(new_n799));
  OAI21_X1  g598(.A(G92gat), .B1(new_n799), .B2(new_n430), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n797), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(KEYINPUT113), .B1(new_n779), .B2(new_n781), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n776), .ZN(new_n803));
  OAI211_X1 g602(.A(KEYINPUT113), .B(KEYINPUT51), .C1(new_n779), .C2(new_n781), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n803), .A2(new_n804), .A3(new_n796), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n805), .A2(new_n800), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n801), .B1(new_n806), .B2(new_n798), .ZN(G1337gat));
  NOR2_X1   g606(.A1(new_n757), .A2(G99gat), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n795), .A2(new_n745), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(G99gat), .B1(new_n799), .B2(new_n676), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(G1338gat));
  NAND4_X1  g610(.A1(new_n763), .A2(new_n447), .A3(new_n765), .A4(new_n768), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(G106gat), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n354), .A2(G106gat), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n782), .A2(new_n787), .A3(new_n745), .A4(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT114), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n815), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n795), .A2(KEYINPUT114), .A3(new_n745), .A4(new_n816), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n354), .A2(G106gat), .A3(new_n654), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n803), .A2(new_n804), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n813), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(KEYINPUT53), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n821), .A2(new_n825), .ZN(G1339gat));
  NAND4_X1  g625(.A1(new_n631), .A2(new_n704), .A3(new_n633), .A4(new_n654), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT55), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n641), .A2(new_n613), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n641), .A2(new_n613), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n644), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n583), .A2(KEYINPUT10), .A3(new_n615), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n831), .A2(new_n635), .A3(new_n832), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n646), .A2(new_n833), .A3(KEYINPUT54), .ZN(new_n834));
  XNOR2_X1  g633(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n636), .B(new_n835), .C1(new_n643), .C2(new_n645), .ZN(new_n836));
  INV_X1    g635(.A(new_n650), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n828), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n646), .A2(new_n833), .A3(KEYINPUT54), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n840), .A2(KEYINPUT55), .A3(new_n837), .A4(new_n836), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n563), .A2(new_n839), .A3(new_n651), .A4(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n552), .A2(new_n555), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n540), .B1(new_n547), .B2(new_n549), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n478), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n562), .B(new_n845), .C1(new_n652), .C2(new_n653), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n628), .B1(new_n842), .B2(new_n846), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n628), .A2(new_n839), .A3(new_n651), .A4(new_n841), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n562), .A2(new_n845), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(KEYINPUT116), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n562), .A2(new_n852), .A3(new_n845), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n847), .B1(new_n849), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n827), .B1(new_n599), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(new_n660), .A3(new_n356), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n381), .B1(new_n858), .B2(KEYINPUT117), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n859), .B1(KEYINPUT117), .B2(new_n858), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n860), .A2(new_n704), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n858), .A2(new_n381), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n704), .A2(new_n473), .ZN(new_n863));
  AOI22_X1  g662(.A1(new_n861), .A2(new_n473), .B1(new_n862), .B2(new_n863), .ZN(G1340gat));
  NOR3_X1   g663(.A1(new_n860), .A2(G120gat), .A3(new_n654), .ZN(new_n865));
  INV_X1    g664(.A(G120gat), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n866), .B1(new_n862), .B2(new_n745), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n868), .B(new_n869), .ZN(G1341gat));
  NAND2_X1  g669(.A1(new_n250), .A2(new_n252), .ZN(new_n871));
  INV_X1    g670(.A(new_n862), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n871), .B1(new_n872), .B2(new_n702), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n599), .A2(new_n250), .A3(new_n252), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n873), .B1(new_n860), .B2(new_n874), .ZN(G1342gat));
  OR3_X1    g674(.A1(new_n860), .A2(G134gat), .A3(new_n629), .ZN(new_n876));
  OR2_X1    g675(.A1(new_n876), .A2(KEYINPUT56), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(KEYINPUT56), .ZN(new_n878));
  OAI21_X1  g677(.A(G134gat), .B1(new_n872), .B2(new_n629), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(G1343gat));
  NOR3_X1   g679(.A1(new_n677), .A2(new_n659), .A3(new_n381), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n857), .A2(new_n447), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n882), .A2(KEYINPUT57), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n857), .A2(KEYINPUT57), .A3(new_n447), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(G141gat), .B1(new_n885), .B2(new_n704), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n881), .A2(new_n882), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(new_n476), .A3(new_n563), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  XOR2_X1   g688(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n890));
  XNOR2_X1  g689(.A(new_n889), .B(new_n890), .ZN(G1344gat));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n892), .B(G148gat), .C1(new_n885), .C2(new_n654), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT123), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n854), .B1(KEYINPUT120), .B2(new_n848), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n839), .A2(new_n651), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n896), .A2(new_n897), .A3(new_n628), .A4(new_n841), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n847), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT121), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n702), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AOI211_X1 g700(.A(KEYINPUT121), .B(new_n847), .C1(new_n898), .C2(new_n895), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n827), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n354), .B1(new_n903), .B2(KEYINPUT122), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n905), .B(new_n827), .C1(new_n901), .C2(new_n902), .ZN(new_n906));
  AOI21_X1  g705(.A(KEYINPUT57), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n745), .B(new_n881), .C1(new_n907), .C2(new_n884), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(G148gat), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n894), .B1(new_n909), .B2(KEYINPUT59), .ZN(new_n910));
  AOI211_X1 g709(.A(KEYINPUT123), .B(new_n892), .C1(new_n908), .C2(G148gat), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n893), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(G148gat), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n887), .A2(new_n913), .A3(new_n745), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n914), .ZN(G1345gat));
  INV_X1    g714(.A(new_n301), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n916), .B1(new_n885), .B2(new_n702), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n887), .A2(new_n301), .A3(new_n599), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(G1346gat));
  OAI21_X1  g718(.A(G162gat), .B1(new_n885), .B2(new_n629), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n887), .A2(new_n302), .A3(new_n628), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1347gat));
  NOR3_X1   g721(.A1(new_n355), .A2(new_n660), .A3(new_n430), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n857), .A2(new_n563), .A3(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(G169gat), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n925), .A2(KEYINPUT124), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n925), .A2(KEYINPUT124), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n924), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n928), .B1(new_n924), .B2(new_n926), .ZN(G1348gat));
  NAND2_X1  g728(.A1(new_n857), .A2(new_n923), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n930), .A2(new_n654), .ZN(new_n931));
  XOR2_X1   g730(.A(new_n931), .B(G176gat), .Z(G1349gat));
  NOR2_X1   g731(.A1(new_n930), .A2(new_n702), .ZN(new_n933));
  MUX2_X1   g732(.A(new_n217), .B(new_n221), .S(new_n933), .Z(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT60), .ZN(G1350gat));
  NOR2_X1   g734(.A1(new_n930), .A2(new_n629), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT61), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n937), .B2(new_n222), .ZN(new_n938));
  XOR2_X1   g737(.A(KEYINPUT61), .B(G190gat), .Z(new_n939));
  OAI21_X1  g738(.A(new_n938), .B1(new_n936), .B2(new_n939), .ZN(G1351gat));
  NOR2_X1   g739(.A1(new_n660), .A2(new_n430), .ZN(new_n941));
  AND3_X1   g740(.A1(new_n882), .A2(new_n676), .A3(new_n941), .ZN(new_n942));
  XNOR2_X1  g741(.A(KEYINPUT125), .B(G197gat), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n942), .A2(new_n563), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n676), .A2(new_n941), .ZN(new_n945));
  INV_X1    g744(.A(new_n907), .ZN(new_n946));
  INV_X1    g745(.A(new_n884), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n948), .A2(new_n563), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n944), .B1(new_n949), .B2(new_n943), .ZN(G1352gat));
  XNOR2_X1  g749(.A(KEYINPUT126), .B(G204gat), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n942), .A2(new_n745), .A3(new_n951), .ZN(new_n952));
  XOR2_X1   g751(.A(new_n952), .B(KEYINPUT62), .Z(new_n953));
  AOI211_X1 g752(.A(new_n654), .B(new_n945), .C1(new_n946), .C2(new_n947), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n953), .B1(new_n954), .B2(new_n951), .ZN(G1353gat));
  NAND3_X1  g754(.A1(new_n942), .A2(new_n313), .A3(new_n599), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n948), .A2(new_n599), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n957), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n958));
  AOI21_X1  g757(.A(KEYINPUT63), .B1(new_n957), .B2(G211gat), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(G1354gat));
  AOI21_X1  g759(.A(G218gat), .B1(new_n942), .B2(new_n628), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n628), .A2(G218gat), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n962), .B(KEYINPUT127), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n961), .B1(new_n948), .B2(new_n963), .ZN(G1355gat));
endmodule


