

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765;

  NAND2_X1 U374 ( .A1(n353), .A2(n641), .ZN(n757) );
  XNOR2_X1 U375 ( .A(n629), .B(n628), .ZN(n353) );
  AND2_X1 U376 ( .A1(n764), .A2(n671), .ZN(n367) );
  XOR2_X1 U377 ( .A(n585), .B(KEYINPUT38), .Z(n710) );
  XNOR2_X1 U378 ( .A(n607), .B(n509), .ZN(n597) );
  XNOR2_X1 U379 ( .A(n678), .B(n418), .ZN(n631) );
  XNOR2_X1 U380 ( .A(n520), .B(KEYINPUT4), .ZN(n499) );
  XNOR2_X1 U381 ( .A(n457), .B(G131), .ZN(n532) );
  INV_X1 U382 ( .A(KEYINPUT70), .ZN(n457) );
  NOR2_X2 U383 ( .A1(n352), .A2(n651), .ZN(n653) );
  AND2_X2 U384 ( .A1(n648), .A2(n647), .ZN(n352) );
  XNOR2_X2 U385 ( .A(n539), .B(n540), .ZN(n566) );
  NAND2_X1 U386 ( .A1(n517), .A2(n552), .ZN(n395) );
  XNOR2_X2 U387 ( .A(n492), .B(n369), .ZN(n517) );
  XNOR2_X2 U388 ( .A(n699), .B(n461), .ZN(n603) );
  NAND2_X1 U389 ( .A1(n402), .A2(n354), .ZN(n406) );
  NAND2_X1 U390 ( .A1(n363), .A2(n436), .ZN(n354) );
  OR2_X2 U391 ( .A1(n661), .A2(G902), .ZN(n460) );
  NOR2_X2 U392 ( .A1(n566), .A2(n565), .ZN(n678) );
  XOR2_X1 U393 ( .A(KEYINPUT16), .B(KEYINPUT77), .Z(n355) );
  XNOR2_X2 U394 ( .A(n622), .B(KEYINPUT1), .ZN(n633) );
  OR2_X1 U395 ( .A1(n555), .A2(n549), .ZN(n691) );
  INV_X1 U396 ( .A(n753), .ZN(n407) );
  NOR2_X1 U397 ( .A1(n740), .A2(n646), .ZN(n648) );
  AND2_X1 U398 ( .A1(n404), .A2(n403), .ZN(n402) );
  XNOR2_X1 U399 ( .A(n476), .B(n475), .ZN(n555) );
  OR2_X1 U400 ( .A1(n729), .A2(G902), .ZN(n490) );
  XNOR2_X1 U401 ( .A(n410), .B(n407), .ZN(n736) );
  XNOR2_X1 U402 ( .A(n412), .B(n411), .ZN(n410) );
  XNOR2_X1 U403 ( .A(n751), .B(n459), .ZN(n487) );
  XNOR2_X1 U404 ( .A(n499), .B(n435), .ZN(n751) );
  XNOR2_X1 U405 ( .A(n409), .B(n536), .ZN(n753) );
  XNOR2_X1 U406 ( .A(n467), .B(KEYINPUT23), .ZN(n411) );
  XNOR2_X1 U407 ( .A(n532), .B(n458), .ZN(n435) );
  XNOR2_X1 U408 ( .A(n500), .B(n408), .ZN(n536) );
  INV_X2 U409 ( .A(G122), .ZN(n438) );
  INV_X2 U410 ( .A(G953), .ZN(n759) );
  XNOR2_X1 U411 ( .A(KEYINPUT15), .B(G902), .ZN(n646) );
  NOR2_X2 U412 ( .A1(n687), .A2(n653), .ZN(n356) );
  NOR2_X1 U413 ( .A1(n687), .A2(n653), .ZN(n357) );
  XNOR2_X1 U414 ( .A(n516), .B(KEYINPUT0), .ZN(n358) );
  INV_X1 U415 ( .A(n439), .ZN(n359) );
  NOR2_X1 U416 ( .A1(n687), .A2(n653), .ZN(n735) );
  XNOR2_X1 U417 ( .A(n516), .B(KEYINPUT0), .ZN(n552) );
  XNOR2_X1 U418 ( .A(n544), .B(n370), .ZN(n546) );
  XNOR2_X1 U419 ( .A(KEYINPUT67), .B(G101), .ZN(n497) );
  XOR2_X1 U420 ( .A(G125), .B(G146), .Z(n500) );
  XNOR2_X1 U421 ( .A(n454), .B(n453), .ZN(n493) );
  XNOR2_X1 U422 ( .A(KEYINPUT74), .B(KEYINPUT3), .ZN(n453) );
  XNOR2_X1 U423 ( .A(n422), .B(n419), .ZN(n654) );
  XNOR2_X1 U424 ( .A(n421), .B(n522), .ZN(n419) );
  XNOR2_X1 U425 ( .A(n525), .B(n523), .ZN(n422) );
  XNOR2_X1 U426 ( .A(n521), .B(n458), .ZN(n421) );
  INV_X1 U427 ( .A(n654), .ZN(n385) );
  XOR2_X1 U428 ( .A(KEYINPUT97), .B(G140), .Z(n530) );
  XOR2_X1 U429 ( .A(KEYINPUT91), .B(KEYINPUT24), .Z(n469) );
  XNOR2_X1 U430 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n496) );
  NAND2_X1 U431 ( .A1(n584), .A2(n514), .ZN(n515) );
  NAND2_X1 U432 ( .A1(G898), .A2(G953), .ZN(n514) );
  XOR2_X1 U433 ( .A(KEYINPUT5), .B(G137), .Z(n448) );
  XNOR2_X1 U434 ( .A(n495), .B(n394), .ZN(n423) );
  XNOR2_X1 U435 ( .A(n437), .B(n494), .ZN(n495) );
  XNOR2_X1 U436 ( .A(n533), .B(n355), .ZN(n437) );
  INV_X1 U437 ( .A(n484), .ZN(n409) );
  NOR2_X1 U438 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U439 ( .A1(n413), .A2(n555), .ZN(n442) );
  NOR2_X1 U440 ( .A1(n381), .A2(n739), .ZN(n380) );
  NAND2_X1 U441 ( .A1(n356), .A2(n375), .ZN(n382) );
  NAND2_X1 U442 ( .A1(n689), .A2(n759), .ZN(n428) );
  XNOR2_X1 U443 ( .A(n688), .B(KEYINPUT85), .ZN(n429) );
  INV_X1 U444 ( .A(KEYINPUT68), .ZN(n426) );
  INV_X1 U445 ( .A(n638), .ZN(n585) );
  XNOR2_X1 U446 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n521) );
  XOR2_X1 U447 ( .A(G122), .B(KEYINPUT99), .Z(n519) );
  XNOR2_X1 U448 ( .A(n420), .B(G107), .ZN(n522) );
  INV_X1 U449 ( .A(G116), .ZN(n420) );
  XNOR2_X1 U450 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U451 ( .A(G143), .B(G113), .ZN(n529) );
  XNOR2_X1 U452 ( .A(KEYINPUT11), .B(KEYINPUT96), .ZN(n527) );
  XOR2_X1 U453 ( .A(KEYINPUT98), .B(KEYINPUT12), .Z(n528) );
  INV_X1 U454 ( .A(KEYINPUT10), .ZN(n408) );
  NOR2_X1 U455 ( .A1(n439), .A2(n562), .ZN(n563) );
  NOR2_X1 U456 ( .A1(n416), .A2(n691), .ZN(n611) );
  OR2_X1 U457 ( .A1(n596), .A2(n591), .ZN(n416) );
  NAND2_X1 U458 ( .A1(n622), .A2(n414), .ZN(n413) );
  AND2_X1 U459 ( .A1(n585), .A2(n415), .ZN(n414) );
  NOR2_X1 U460 ( .A1(n549), .A2(n591), .ZN(n415) );
  XNOR2_X1 U461 ( .A(n441), .B(n440), .ZN(n612) );
  XNOR2_X1 U462 ( .A(KEYINPUT107), .B(KEYINPUT30), .ZN(n440) );
  XNOR2_X1 U463 ( .A(n471), .B(n470), .ZN(n412) );
  XNOR2_X1 U464 ( .A(G128), .B(KEYINPUT93), .ZN(n468) );
  XNOR2_X1 U465 ( .A(n482), .B(G110), .ZN(n494) );
  XNOR2_X1 U466 ( .A(KEYINPUT71), .B(G140), .ZN(n464) );
  XNOR2_X1 U467 ( .A(G107), .B(G104), .ZN(n481) );
  XNOR2_X1 U468 ( .A(n423), .B(n503), .ZN(n659) );
  INV_X1 U469 ( .A(KEYINPUT100), .ZN(n418) );
  INV_X1 U470 ( .A(KEYINPUT87), .ZN(n507) );
  XNOR2_X1 U471 ( .A(n606), .B(KEYINPUT106), .ZN(n635) );
  XNOR2_X1 U472 ( .A(KEYINPUT81), .B(KEYINPUT34), .ZN(n518) );
  XNOR2_X1 U473 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U474 ( .A(n617), .B(n399), .ZN(n664) );
  INV_X1 U475 ( .A(KEYINPUT105), .ZN(n399) );
  AND2_X1 U476 ( .A1(n619), .A2(n550), .ZN(n551) );
  XNOR2_X1 U477 ( .A(n487), .B(n388), .ZN(n661) );
  XNOR2_X1 U478 ( .A(n456), .B(n365), .ZN(n388) );
  XNOR2_X1 U479 ( .A(n618), .B(n387), .ZN(n763) );
  XNOR2_X1 U480 ( .A(KEYINPUT110), .B(KEYINPUT40), .ZN(n387) );
  NOR2_X1 U481 ( .A1(n383), .A2(n379), .ZN(n656) );
  NOR2_X1 U482 ( .A1(n357), .A2(n385), .ZN(n383) );
  NAND2_X1 U483 ( .A1(n429), .A2(n427), .ZN(n725) );
  NOR2_X1 U484 ( .A1(n724), .A2(n428), .ZN(n427) );
  AND2_X1 U485 ( .A1(n506), .A2(G210), .ZN(n360) );
  XOR2_X1 U486 ( .A(n528), .B(n527), .Z(n361) );
  AND2_X1 U487 ( .A1(G224), .A2(n759), .ZN(n362) );
  AND2_X1 U488 ( .A1(n590), .A2(n401), .ZN(n363) );
  AND2_X1 U489 ( .A1(n674), .A2(n602), .ZN(n364) );
  AND2_X1 U490 ( .A1(n535), .A2(G210), .ZN(n365) );
  AND2_X1 U491 ( .A1(n588), .A2(KEYINPUT83), .ZN(n366) );
  INV_X1 U492 ( .A(G134), .ZN(n458) );
  NOR2_X1 U493 ( .A1(n718), .A2(n431), .ZN(n368) );
  XOR2_X1 U494 ( .A(KEYINPUT103), .B(KEYINPUT33), .Z(n369) );
  XOR2_X1 U495 ( .A(KEYINPUT86), .B(KEYINPUT35), .Z(n370) );
  XOR2_X1 U496 ( .A(n729), .B(n728), .Z(n371) );
  XNOR2_X1 U497 ( .A(n734), .B(n733), .ZN(n372) );
  XOR2_X1 U498 ( .A(n659), .B(n658), .Z(n373) );
  XOR2_X1 U499 ( .A(n661), .B(KEYINPUT62), .Z(n374) );
  AND2_X1 U500 ( .A1(n385), .A2(G478), .ZN(n375) );
  XNOR2_X1 U501 ( .A(KEYINPUT119), .B(KEYINPUT56), .ZN(n376) );
  XOR2_X1 U502 ( .A(KEYINPUT60), .B(KEYINPUT66), .Z(n377) );
  INV_X1 U503 ( .A(n739), .ZN(n384) );
  NAND2_X1 U504 ( .A1(n382), .A2(n380), .ZN(n379) );
  XNOR2_X1 U505 ( .A(n444), .B(n600), .ZN(n443) );
  XNOR2_X1 U506 ( .A(n378), .B(n361), .ZN(n538) );
  XNOR2_X1 U507 ( .A(n534), .B(n531), .ZN(n378) );
  NAND2_X1 U508 ( .A1(n714), .A2(KEYINPUT47), .ZN(n590) );
  XNOR2_X2 U509 ( .A(n417), .B(KEYINPUT101), .ZN(n714) );
  NOR2_X1 U510 ( .A1(n664), .A2(n603), .ZN(n605) );
  XNOR2_X2 U511 ( .A(n645), .B(KEYINPUT80), .ZN(n687) );
  NOR2_X1 U512 ( .A1(n385), .A2(G478), .ZN(n381) );
  XNOR2_X1 U513 ( .A(n502), .B(n501), .ZN(n503) );
  NAND2_X1 U514 ( .A1(n627), .A2(n386), .ZN(n629) );
  XNOR2_X1 U515 ( .A(n626), .B(KEYINPUT46), .ZN(n386) );
  XNOR2_X1 U516 ( .A(n389), .B(KEYINPUT72), .ZN(n627) );
  AND2_X1 U517 ( .A1(n443), .A2(n445), .ZN(n389) );
  INV_X1 U518 ( .A(n358), .ZN(n571) );
  XNOR2_X1 U519 ( .A(n547), .B(n426), .ZN(n425) );
  NAND2_X1 U520 ( .A1(n425), .A2(n367), .ZN(n424) );
  XNOR2_X1 U521 ( .A(n390), .B(n376), .ZN(G51) );
  NAND2_X1 U522 ( .A1(n393), .A2(n384), .ZN(n390) );
  XNOR2_X1 U523 ( .A(n391), .B(KEYINPUT121), .ZN(G54) );
  NAND2_X1 U524 ( .A1(n398), .A2(n384), .ZN(n391) );
  XNOR2_X1 U525 ( .A(n392), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U526 ( .A1(n397), .A2(n384), .ZN(n392) );
  XNOR2_X1 U527 ( .A(n660), .B(n373), .ZN(n393) );
  XNOR2_X1 U528 ( .A(n493), .B(n522), .ZN(n394) );
  XNOR2_X1 U529 ( .A(n395), .B(n518), .ZN(n543) );
  NAND2_X1 U530 ( .A1(n396), .A2(n447), .ZN(n582) );
  XNOR2_X1 U531 ( .A(n424), .B(KEYINPUT76), .ZN(n396) );
  XNOR2_X1 U532 ( .A(n662), .B(n374), .ZN(n397) );
  XNOR2_X1 U533 ( .A(n730), .B(n371), .ZN(n398) );
  NAND2_X1 U534 ( .A1(n566), .A2(n565), .ZN(n617) );
  INV_X1 U535 ( .A(KEYINPUT83), .ZN(n401) );
  NAND2_X1 U536 ( .A1(n589), .A2(n588), .ZN(n436) );
  NAND2_X1 U537 ( .A1(n589), .A2(n366), .ZN(n403) );
  NAND2_X1 U538 ( .A1(n405), .A2(KEYINPUT83), .ZN(n404) );
  INV_X1 U539 ( .A(n590), .ZN(n405) );
  NAND2_X1 U540 ( .A1(n406), .A2(n599), .ZN(n444) );
  NAND2_X1 U541 ( .A1(n631), .A2(n617), .ZN(n417) );
  XNOR2_X1 U542 ( .A(n423), .B(G101), .ZN(n748) );
  XNOR2_X1 U543 ( .A(n538), .B(n537), .ZN(n734) );
  XNOR2_X2 U544 ( .A(n559), .B(KEYINPUT32), .ZN(n764) );
  NAND2_X1 U545 ( .A1(n430), .A2(n517), .ZN(n689) );
  INV_X1 U546 ( .A(n707), .ZN(n430) );
  INV_X1 U547 ( .A(n517), .ZN(n431) );
  XNOR2_X1 U548 ( .A(n432), .B(n377), .ZN(G60) );
  NAND2_X1 U549 ( .A1(n433), .A2(n384), .ZN(n432) );
  XNOR2_X1 U550 ( .A(n434), .B(n372), .ZN(n433) );
  NAND2_X1 U551 ( .A1(n357), .A2(G475), .ZN(n434) );
  XNOR2_X1 U552 ( .A(n436), .B(G143), .ZN(G45) );
  XNOR2_X2 U553 ( .A(n438), .B(G104), .ZN(n533) );
  INV_X1 U554 ( .A(n546), .ZN(n439) );
  XNOR2_X1 U555 ( .A(n359), .B(G122), .ZN(G24) );
  NAND2_X1 U556 ( .A1(n442), .A2(n612), .ZN(n587) );
  NAND2_X1 U557 ( .A1(n699), .A2(n709), .ZN(n441) );
  NOR2_X1 U558 ( .A1(n681), .A2(n364), .ZN(n445) );
  XNOR2_X1 U559 ( .A(n536), .B(n446), .ZN(n537) );
  XNOR2_X2 U560 ( .A(n490), .B(n489), .ZN(n622) );
  XNOR2_X2 U561 ( .A(n505), .B(n360), .ZN(n613) );
  AND2_X1 U562 ( .A1(n535), .A2(G214), .ZN(n446) );
  AND2_X1 U563 ( .A1(n580), .A2(n579), .ZN(n447) );
  INV_X1 U564 ( .A(KEYINPUT84), .ZN(n600) );
  XNOR2_X1 U565 ( .A(n448), .B(G116), .ZN(n455) );
  XNOR2_X1 U566 ( .A(n493), .B(n455), .ZN(n456) );
  XNOR2_X1 U567 ( .A(n500), .B(n362), .ZN(n501) );
  INV_X1 U568 ( .A(KEYINPUT48), .ZN(n628) );
  INV_X1 U569 ( .A(KEYINPUT45), .ZN(n581) );
  NOR2_X2 U570 ( .A1(n597), .A2(n515), .ZN(n516) );
  INV_X1 U571 ( .A(KEYINPUT19), .ZN(n509) );
  INV_X1 U572 ( .A(KEYINPUT36), .ZN(n608) );
  NOR2_X1 U573 ( .A1(n759), .A2(G952), .ZN(n739) );
  INV_X1 U574 ( .A(G119), .ZN(n449) );
  NAND2_X1 U575 ( .A1(G113), .A2(n449), .ZN(n452) );
  INV_X1 U576 ( .A(G113), .ZN(n450) );
  NAND2_X1 U577 ( .A1(n450), .A2(G119), .ZN(n451) );
  NAND2_X1 U578 ( .A1(n452), .A2(n451), .ZN(n454) );
  NOR2_X1 U579 ( .A1(G953), .A2(G237), .ZN(n535) );
  XNOR2_X2 U580 ( .A(G143), .B(G128), .ZN(n520) );
  XNOR2_X1 U581 ( .A(n497), .B(G146), .ZN(n459) );
  XNOR2_X2 U582 ( .A(n460), .B(G472), .ZN(n699) );
  XNOR2_X1 U583 ( .A(KEYINPUT102), .B(KEYINPUT6), .ZN(n461) );
  XNOR2_X1 U584 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n463) );
  NAND2_X1 U585 ( .A1(G234), .A2(n759), .ZN(n462) );
  XNOR2_X1 U586 ( .A(n463), .B(n462), .ZN(n524) );
  NAND2_X1 U587 ( .A1(n524), .A2(G221), .ZN(n471) );
  XNOR2_X1 U588 ( .A(n464), .B(G137), .ZN(n484) );
  XOR2_X1 U589 ( .A(KEYINPUT92), .B(KEYINPUT75), .Z(n466) );
  XNOR2_X1 U590 ( .A(G119), .B(G110), .ZN(n465) );
  XNOR2_X1 U591 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U592 ( .A(n469), .B(n468), .ZN(n470) );
  NOR2_X1 U593 ( .A1(G902), .A2(n736), .ZN(n476) );
  NAND2_X1 U594 ( .A1(n646), .A2(G234), .ZN(n472) );
  XNOR2_X1 U595 ( .A(n472), .B(KEYINPUT20), .ZN(n477) );
  NAND2_X1 U596 ( .A1(n477), .A2(G217), .ZN(n474) );
  INV_X1 U597 ( .A(KEYINPUT25), .ZN(n473) );
  NAND2_X1 U598 ( .A1(G221), .A2(n477), .ZN(n478) );
  XOR2_X1 U599 ( .A(KEYINPUT21), .B(n478), .Z(n695) );
  INV_X1 U600 ( .A(KEYINPUT94), .ZN(n479) );
  XNOR2_X1 U601 ( .A(n695), .B(n479), .ZN(n549) );
  NOR2_X1 U602 ( .A1(n603), .A2(n691), .ZN(n491) );
  NAND2_X1 U603 ( .A1(n759), .A2(G227), .ZN(n480) );
  XNOR2_X1 U604 ( .A(n481), .B(n480), .ZN(n483) );
  INV_X1 U605 ( .A(KEYINPUT90), .ZN(n482) );
  XNOR2_X1 U606 ( .A(n483), .B(n494), .ZN(n485) );
  XNOR2_X1 U607 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U608 ( .A(n487), .B(n486), .ZN(n729) );
  INV_X1 U609 ( .A(KEYINPUT73), .ZN(n488) );
  XNOR2_X1 U610 ( .A(n488), .B(G469), .ZN(n489) );
  NAND2_X1 U611 ( .A1(n491), .A2(n633), .ZN(n492) );
  XNOR2_X1 U612 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U613 ( .A(n499), .B(n498), .ZN(n502) );
  NAND2_X1 U614 ( .A1(n659), .A2(n646), .ZN(n505) );
  NOR2_X1 U615 ( .A1(G902), .A2(G237), .ZN(n504) );
  XOR2_X1 U616 ( .A(KEYINPUT78), .B(n504), .Z(n506) );
  NAND2_X1 U617 ( .A1(n506), .A2(G214), .ZN(n709) );
  NAND2_X1 U618 ( .A1(n613), .A2(n709), .ZN(n508) );
  XNOR2_X2 U619 ( .A(n508), .B(n507), .ZN(n607) );
  NAND2_X1 U620 ( .A1(G237), .A2(G234), .ZN(n510) );
  XNOR2_X1 U621 ( .A(n510), .B(KEYINPUT14), .ZN(n721) );
  OR2_X1 U622 ( .A1(n759), .A2(G902), .ZN(n511) );
  NAND2_X1 U623 ( .A1(n721), .A2(n511), .ZN(n513) );
  NOR2_X1 U624 ( .A1(G953), .A2(G952), .ZN(n512) );
  NOR2_X1 U625 ( .A1(n513), .A2(n512), .ZN(n584) );
  XNOR2_X1 U626 ( .A(n520), .B(n519), .ZN(n523) );
  NAND2_X1 U627 ( .A1(G217), .A2(n524), .ZN(n525) );
  NOR2_X1 U628 ( .A1(G902), .A2(n654), .ZN(n526) );
  XNOR2_X1 U629 ( .A(G478), .B(n526), .ZN(n565) );
  INV_X1 U630 ( .A(n565), .ZN(n548) );
  XNOR2_X1 U631 ( .A(KEYINPUT13), .B(G475), .ZN(n540) );
  XNOR2_X1 U632 ( .A(n533), .B(n532), .ZN(n534) );
  NOR2_X1 U633 ( .A1(G902), .A2(n734), .ZN(n539) );
  NAND2_X1 U634 ( .A1(n548), .A2(n566), .ZN(n542) );
  INV_X1 U635 ( .A(KEYINPUT104), .ZN(n541) );
  XNOR2_X1 U636 ( .A(n542), .B(n541), .ZN(n588) );
  NAND2_X1 U637 ( .A1(n543), .A2(n588), .ZN(n544) );
  INV_X1 U638 ( .A(KEYINPUT44), .ZN(n545) );
  NAND2_X1 U639 ( .A1(n546), .A2(n545), .ZN(n547) );
  INV_X1 U640 ( .A(KEYINPUT22), .ZN(n554) );
  NOR2_X1 U641 ( .A1(n566), .A2(n548), .ZN(n619) );
  INV_X1 U642 ( .A(n549), .ZN(n550) );
  NAND2_X1 U643 ( .A1(n358), .A2(n551), .ZN(n553) );
  XNOR2_X1 U644 ( .A(n554), .B(n553), .ZN(n577) );
  INV_X1 U645 ( .A(n555), .ZN(n696) );
  NAND2_X1 U646 ( .A1(n603), .A2(n555), .ZN(n556) );
  INV_X1 U647 ( .A(n633), .ZN(n690) );
  NOR2_X1 U648 ( .A1(n556), .A2(n690), .ZN(n557) );
  XNOR2_X1 U649 ( .A(n557), .B(KEYINPUT82), .ZN(n558) );
  NAND2_X1 U650 ( .A1(n577), .A2(n558), .ZN(n559) );
  INV_X1 U651 ( .A(n699), .ZN(n567) );
  NAND2_X1 U652 ( .A1(n555), .A2(n567), .ZN(n560) );
  NOR2_X1 U653 ( .A1(n560), .A2(n633), .ZN(n561) );
  NAND2_X1 U654 ( .A1(n577), .A2(n561), .ZN(n671) );
  INV_X1 U655 ( .A(n671), .ZN(n562) );
  NAND2_X1 U656 ( .A1(n563), .A2(n764), .ZN(n564) );
  NAND2_X1 U657 ( .A1(n564), .A2(KEYINPUT44), .ZN(n580) );
  NOR2_X1 U658 ( .A1(n691), .A2(n567), .ZN(n568) );
  NAND2_X1 U659 ( .A1(n568), .A2(n633), .ZN(n704) );
  NOR2_X1 U660 ( .A1(n571), .A2(n704), .ZN(n569) );
  XOR2_X1 U661 ( .A(KEYINPUT31), .B(n569), .Z(n679) );
  INV_X1 U662 ( .A(n622), .ZN(n596) );
  OR2_X1 U663 ( .A1(n691), .A2(n596), .ZN(n570) );
  NOR2_X1 U664 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U665 ( .A(n572), .B(KEYINPUT95), .ZN(n573) );
  NOR2_X1 U666 ( .A1(n699), .A2(n573), .ZN(n667) );
  NOR2_X1 U667 ( .A1(n679), .A2(n667), .ZN(n574) );
  NOR2_X1 U668 ( .A1(n714), .A2(n574), .ZN(n578) );
  NAND2_X1 U669 ( .A1(n603), .A2(n696), .ZN(n575) );
  NOR2_X1 U670 ( .A1(n575), .A2(n633), .ZN(n576) );
  AND2_X1 U671 ( .A1(n577), .A2(n576), .ZN(n663) );
  NOR2_X1 U672 ( .A1(n578), .A2(n663), .ZN(n579) );
  XNOR2_X2 U673 ( .A(n582), .B(n581), .ZN(n740) );
  NAND2_X1 U674 ( .A1(G953), .A2(G900), .ZN(n583) );
  NAND2_X1 U675 ( .A1(n584), .A2(n583), .ZN(n591) );
  INV_X1 U676 ( .A(n613), .ZN(n638) );
  INV_X1 U677 ( .A(KEYINPUT108), .ZN(n586) );
  XNOR2_X1 U678 ( .A(n587), .B(n586), .ZN(n589) );
  INV_X1 U679 ( .A(n591), .ZN(n592) );
  NAND2_X1 U680 ( .A1(n695), .A2(n592), .ZN(n593) );
  NOR2_X1 U681 ( .A1(n696), .A2(n593), .ZN(n604) );
  AND2_X1 U682 ( .A1(n699), .A2(n604), .ZN(n595) );
  XOR2_X1 U683 ( .A(KEYINPUT109), .B(KEYINPUT28), .Z(n594) );
  XNOR2_X1 U684 ( .A(n595), .B(n594), .ZN(n623) );
  NOR2_X1 U685 ( .A1(n597), .A2(n596), .ZN(n601) );
  NAND2_X1 U686 ( .A1(n623), .A2(n601), .ZN(n598) );
  NAND2_X1 U687 ( .A1(KEYINPUT47), .A2(n598), .ZN(n599) );
  AND2_X1 U688 ( .A1(n623), .A2(n601), .ZN(n674) );
  NOR2_X1 U689 ( .A1(KEYINPUT47), .A2(n714), .ZN(n602) );
  NAND2_X1 U690 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U691 ( .A1(n635), .A2(n607), .ZN(n609) );
  XNOR2_X1 U692 ( .A(n609), .B(n608), .ZN(n610) );
  NOR2_X1 U693 ( .A1(n610), .A2(n690), .ZN(n681) );
  NAND2_X1 U694 ( .A1(n612), .A2(n611), .ZN(n615) );
  INV_X1 U695 ( .A(n710), .ZN(n614) );
  XNOR2_X1 U696 ( .A(n616), .B(KEYINPUT39), .ZN(n630) );
  NOR2_X1 U697 ( .A1(n617), .A2(n630), .ZN(n618) );
  NAND2_X1 U698 ( .A1(n710), .A2(n709), .ZN(n713) );
  INV_X1 U699 ( .A(n619), .ZN(n712) );
  NOR2_X1 U700 ( .A1(n713), .A2(n712), .ZN(n621) );
  XOR2_X1 U701 ( .A(KEYINPUT111), .B(KEYINPUT41), .Z(n620) );
  XNOR2_X1 U702 ( .A(n621), .B(n620), .ZN(n707) );
  NAND2_X1 U703 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U704 ( .A1(n707), .A2(n624), .ZN(n625) );
  XNOR2_X1 U705 ( .A(KEYINPUT42), .B(n625), .ZN(n765) );
  NOR2_X1 U706 ( .A1(n763), .A2(n765), .ZN(n626) );
  NOR2_X1 U707 ( .A1(n631), .A2(n630), .ZN(n683) );
  INV_X1 U708 ( .A(n683), .ZN(n640) );
  INV_X1 U709 ( .A(n709), .ZN(n632) );
  OR2_X1 U710 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U711 ( .A1(n635), .A2(n634), .ZN(n637) );
  INV_X1 U712 ( .A(KEYINPUT43), .ZN(n636) );
  XNOR2_X1 U713 ( .A(n637), .B(n636), .ZN(n639) );
  NAND2_X1 U714 ( .A1(n639), .A2(n638), .ZN(n684) );
  AND2_X1 U715 ( .A1(n640), .A2(n684), .ZN(n641) );
  INV_X1 U716 ( .A(n757), .ZN(n643) );
  NAND2_X1 U717 ( .A1(n643), .A2(KEYINPUT2), .ZN(n644) );
  NOR2_X2 U718 ( .A1(n740), .A2(n644), .ZN(n645) );
  INV_X1 U719 ( .A(n646), .ZN(n649) );
  XNOR2_X1 U720 ( .A(n757), .B(KEYINPUT79), .ZN(n647) );
  NAND2_X1 U721 ( .A1(KEYINPUT2), .A2(n649), .ZN(n650) );
  XNOR2_X1 U722 ( .A(KEYINPUT65), .B(n650), .ZN(n651) );
  INV_X1 U723 ( .A(KEYINPUT123), .ZN(n655) );
  XNOR2_X1 U724 ( .A(n656), .B(n655), .ZN(G63) );
  NAND2_X1 U725 ( .A1(n356), .A2(G210), .ZN(n660) );
  XNOR2_X1 U726 ( .A(KEYINPUT88), .B(KEYINPUT54), .ZN(n657) );
  XNOR2_X1 U727 ( .A(n657), .B(KEYINPUT55), .ZN(n658) );
  NAND2_X1 U728 ( .A1(n735), .A2(G472), .ZN(n662) );
  XOR2_X1 U729 ( .A(G101), .B(n663), .Z(G3) );
  INV_X1 U730 ( .A(n664), .ZN(n676) );
  NAND2_X1 U731 ( .A1(n667), .A2(n676), .ZN(n665) );
  XNOR2_X1 U732 ( .A(n665), .B(KEYINPUT112), .ZN(n666) );
  XNOR2_X1 U733 ( .A(G104), .B(n666), .ZN(G6) );
  XOR2_X1 U734 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n669) );
  NAND2_X1 U735 ( .A1(n667), .A2(n678), .ZN(n668) );
  XNOR2_X1 U736 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U737 ( .A(G107), .B(n670), .ZN(G9) );
  XNOR2_X1 U738 ( .A(G110), .B(n671), .ZN(G12) );
  XOR2_X1 U739 ( .A(G128), .B(KEYINPUT29), .Z(n673) );
  NAND2_X1 U740 ( .A1(n674), .A2(n678), .ZN(n672) );
  XNOR2_X1 U741 ( .A(n673), .B(n672), .ZN(G30) );
  NAND2_X1 U742 ( .A1(n674), .A2(n676), .ZN(n675) );
  XNOR2_X1 U743 ( .A(n675), .B(G146), .ZN(G48) );
  NAND2_X1 U744 ( .A1(n679), .A2(n676), .ZN(n677) );
  XNOR2_X1 U745 ( .A(n677), .B(G113), .ZN(G15) );
  NAND2_X1 U746 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U747 ( .A(n680), .B(G116), .ZN(G18) );
  XNOR2_X1 U748 ( .A(n681), .B(G125), .ZN(n682) );
  XNOR2_X1 U749 ( .A(n682), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U750 ( .A(G134), .B(n683), .Z(G36) );
  XNOR2_X1 U751 ( .A(G140), .B(n684), .ZN(G42) );
  XOR2_X1 U752 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n726) );
  NOR2_X1 U753 ( .A1(n757), .A2(n740), .ZN(n685) );
  NOR2_X1 U754 ( .A1(n685), .A2(KEYINPUT2), .ZN(n686) );
  NOR2_X1 U755 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U756 ( .A1(n691), .A2(n690), .ZN(n694) );
  XOR2_X1 U757 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n692) );
  XNOR2_X1 U758 ( .A(KEYINPUT50), .B(n692), .ZN(n693) );
  XNOR2_X1 U759 ( .A(n694), .B(n693), .ZN(n702) );
  NOR2_X1 U760 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U761 ( .A(KEYINPUT49), .B(n697), .Z(n698) );
  NOR2_X1 U762 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U763 ( .A(KEYINPUT113), .B(n700), .Z(n701) );
  NAND2_X1 U764 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U765 ( .A(n703), .B(KEYINPUT116), .ZN(n705) );
  NAND2_X1 U766 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U767 ( .A(KEYINPUT51), .B(n706), .ZN(n708) );
  NOR2_X1 U768 ( .A1(n708), .A2(n707), .ZN(n719) );
  NOR2_X1 U769 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U770 ( .A1(n712), .A2(n711), .ZN(n716) );
  NOR2_X1 U771 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U772 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U773 ( .A(KEYINPUT117), .B(n717), .Z(n718) );
  NOR2_X1 U774 ( .A1(n719), .A2(n368), .ZN(n720) );
  XNOR2_X1 U775 ( .A(KEYINPUT52), .B(n720), .ZN(n723) );
  NAND2_X1 U776 ( .A1(n721), .A2(G952), .ZN(n722) );
  NOR2_X1 U777 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U778 ( .A(n726), .B(n725), .ZN(G75) );
  NAND2_X1 U779 ( .A1(n735), .A2(G469), .ZN(n730) );
  XOR2_X1 U780 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n727) );
  XNOR2_X1 U781 ( .A(n727), .B(KEYINPUT120), .ZN(n728) );
  XOR2_X1 U782 ( .A(KEYINPUT89), .B(KEYINPUT64), .Z(n732) );
  XNOR2_X1 U783 ( .A(KEYINPUT122), .B(KEYINPUT59), .ZN(n731) );
  XNOR2_X1 U784 ( .A(n732), .B(n731), .ZN(n733) );
  NAND2_X1 U785 ( .A1(n356), .A2(G217), .ZN(n737) );
  XNOR2_X1 U786 ( .A(n737), .B(n736), .ZN(n738) );
  NOR2_X1 U787 ( .A1(n739), .A2(n738), .ZN(G66) );
  NOR2_X1 U788 ( .A1(n740), .A2(G953), .ZN(n745) );
  NAND2_X1 U789 ( .A1(G953), .A2(G224), .ZN(n741) );
  XNOR2_X1 U790 ( .A(KEYINPUT61), .B(n741), .ZN(n742) );
  NAND2_X1 U791 ( .A1(n742), .A2(G898), .ZN(n743) );
  XOR2_X1 U792 ( .A(KEYINPUT124), .B(n743), .Z(n744) );
  NOR2_X1 U793 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U794 ( .A(n746), .B(KEYINPUT125), .ZN(n750) );
  NOR2_X1 U795 ( .A1(n759), .A2(G898), .ZN(n747) );
  NOR2_X1 U796 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U797 ( .A(n750), .B(n749), .ZN(G69) );
  XNOR2_X1 U798 ( .A(n751), .B(KEYINPUT126), .ZN(n752) );
  XNOR2_X1 U799 ( .A(n753), .B(n752), .ZN(n758) );
  XNOR2_X1 U800 ( .A(KEYINPUT127), .B(n758), .ZN(n754) );
  XNOR2_X1 U801 ( .A(G227), .B(n754), .ZN(n755) );
  NAND2_X1 U802 ( .A1(n755), .A2(G900), .ZN(n756) );
  NAND2_X1 U803 ( .A1(n756), .A2(G953), .ZN(n762) );
  XOR2_X1 U804 ( .A(n758), .B(n757), .Z(n760) );
  NAND2_X1 U805 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U806 ( .A1(n762), .A2(n761), .ZN(G72) );
  XOR2_X1 U807 ( .A(n763), .B(G131), .Z(G33) );
  XNOR2_X1 U808 ( .A(n764), .B(G119), .ZN(G21) );
  XOR2_X1 U809 ( .A(G137), .B(n765), .Z(G39) );
endmodule

