//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 0 0 0 1 1 0 0 1 1 0 0 1 0 1 1 0 0 0 0 1 1 0 0 1 0 1 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  OAI21_X1  g001(.A(G210), .B1(G237), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT6), .ZN(new_n189));
  INV_X1    g003(.A(G104), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT3), .B1(new_n190), .B2(G107), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT3), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G104), .ZN(new_n194));
  INV_X1    g008(.A(G101), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n190), .A2(G107), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n191), .A2(new_n194), .A3(new_n195), .A4(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n190), .A2(G107), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n193), .A2(G104), .ZN(new_n199));
  OAI21_X1  g013(.A(G101), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n197), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G119), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G116), .ZN(new_n204));
  INV_X1    g018(.A(G116), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G119), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT2), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(G113), .ZN(new_n208));
  INV_X1    g022(.A(G113), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(KEYINPUT2), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n204), .B(new_n206), .C1(new_n208), .C2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n204), .A2(new_n206), .A3(KEYINPUT5), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n212), .B(G113), .C1(KEYINPUT5), .C2(new_n204), .ZN(new_n213));
  AND3_X1   g027(.A1(new_n202), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n191), .A2(new_n194), .A3(new_n196), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G101), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(KEYINPUT4), .A3(new_n197), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT80), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n197), .A2(KEYINPUT4), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT80), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n220), .A3(new_n216), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT81), .B(KEYINPUT4), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n215), .A2(G101), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n204), .A2(new_n206), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT2), .B(G113), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n211), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n211), .A2(new_n228), .A3(KEYINPUT66), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n225), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n214), .B1(new_n222), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(G110), .B(G122), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n189), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n235), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n211), .A2(new_n228), .A3(KEYINPUT66), .ZN(new_n238));
  AOI21_X1  g052(.A(KEYINPUT66), .B1(new_n211), .B2(new_n228), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n224), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n240), .B1(new_n221), .B2(new_n218), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n237), .B1(new_n241), .B2(new_n214), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n236), .A2(new_n242), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n189), .B(new_n237), .C1(new_n241), .C2(new_n214), .ZN(new_n244));
  XNOR2_X1  g058(.A(G143), .B(G146), .ZN(new_n245));
  XNOR2_X1  g059(.A(KEYINPUT0), .B(G128), .ZN(new_n246));
  OAI21_X1  g060(.A(KEYINPUT64), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G146), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G143), .ZN(new_n249));
  INV_X1    g063(.A(G143), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G146), .ZN(new_n251));
  AND2_X1   g065(.A1(KEYINPUT0), .A2(G128), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n249), .A2(new_n251), .ZN(new_n255));
  NOR2_X1   g069(.A1(KEYINPUT0), .A2(G128), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT64), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n255), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n247), .A2(new_n254), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G125), .ZN(new_n261));
  OAI21_X1  g075(.A(KEYINPUT1), .B1(new_n250), .B2(G146), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n250), .A2(G146), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n248), .A2(G143), .ZN(new_n264));
  OAI211_X1 g078(.A(G128), .B(new_n262), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G128), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n249), .B(new_n251), .C1(KEYINPUT1), .C2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G125), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n268), .A2(KEYINPUT84), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT84), .B1(new_n268), .B2(new_n269), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n261), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G224), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n273), .A2(G953), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n272), .B(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n243), .A2(new_n244), .A3(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT85), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n243), .A2(new_n244), .A3(KEYINPUT85), .A4(new_n275), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G902), .ZN(new_n281));
  INV_X1    g095(.A(new_n274), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n261), .A2(KEYINPUT86), .B1(KEYINPUT7), .B2(new_n282), .ZN(new_n283));
  OR2_X1    g097(.A1(new_n283), .A2(new_n272), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n272), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n235), .B(KEYINPUT8), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n202), .B1(new_n211), .B2(new_n213), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n286), .B1(new_n214), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n284), .A2(new_n285), .A3(new_n288), .ZN(new_n289));
  NOR3_X1   g103(.A1(new_n241), .A2(new_n237), .A3(new_n214), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n281), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n188), .B1(new_n280), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n188), .ZN(new_n294));
  AOI211_X1 g108(.A(new_n294), .B(new_n291), .C1(new_n278), .C2(new_n279), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n187), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT16), .ZN(new_n297));
  INV_X1    g111(.A(G140), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n298), .A3(G125), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(G125), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n269), .A2(G140), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n299), .B1(new_n302), .B2(new_n297), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n248), .ZN(new_n304));
  OAI211_X1 g118(.A(G146), .B(new_n299), .C1(new_n302), .C2(new_n297), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G237), .ZN(new_n308));
  INV_X1    g122(.A(G953), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(new_n309), .A3(G214), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n310), .B(new_n250), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(KEYINPUT17), .A3(G131), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(G131), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n310), .B(G143), .ZN(new_n314));
  INV_X1    g128(.A(G131), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n307), .B(new_n312), .C1(new_n317), .C2(KEYINPUT17), .ZN(new_n318));
  XNOR2_X1  g132(.A(G113), .B(G122), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n319), .B(new_n190), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n302), .A2(KEYINPUT75), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT75), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n300), .A2(new_n301), .A3(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n321), .A2(new_n248), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n302), .A2(G146), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(KEYINPUT18), .A2(G131), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n311), .A2(KEYINPUT87), .A3(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT87), .ZN(new_n329));
  AOI22_X1  g143(.A1(new_n314), .A2(new_n329), .B1(KEYINPUT18), .B2(G131), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n326), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n318), .A2(new_n320), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n320), .B1(new_n318), .B2(new_n331), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n281), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G475), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n317), .A2(new_n305), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT19), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n321), .A2(new_n338), .A3(new_n323), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n302), .A2(KEYINPUT19), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n341), .A2(G146), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n331), .B1(new_n337), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n320), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n332), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT20), .ZN(new_n347));
  NOR2_X1   g161(.A1(G475), .A2(G902), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n347), .B1(new_n346), .B2(new_n348), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n336), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n309), .A2(G952), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n352), .B1(G234), .B2(G237), .ZN(new_n353));
  AOI211_X1 g167(.A(new_n281), .B(new_n309), .C1(G234), .C2(G237), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT21), .B(G898), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(KEYINPUT13), .B1(new_n266), .B2(G143), .ZN(new_n357));
  INV_X1    g171(.A(G134), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(G128), .B(G143), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n359), .B(new_n360), .ZN(new_n361));
  OR2_X1    g175(.A1(KEYINPUT88), .A2(G122), .ZN(new_n362));
  NAND2_X1  g176(.A1(KEYINPUT88), .A2(G122), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n205), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n205), .A2(G122), .ZN(new_n366));
  AND3_X1   g180(.A1(new_n365), .A2(new_n193), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n193), .B1(new_n365), .B2(new_n366), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n361), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n366), .B(KEYINPUT14), .ZN(new_n370));
  OAI21_X1  g184(.A(G107), .B1(new_n370), .B2(new_n364), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n365), .A2(new_n193), .A3(new_n366), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n360), .B(new_n358), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n369), .A2(new_n374), .ZN(new_n375));
  XOR2_X1   g189(.A(KEYINPUT9), .B(G234), .Z(new_n376));
  XNOR2_X1  g190(.A(new_n376), .B(KEYINPUT79), .ZN(new_n377));
  INV_X1    g191(.A(G217), .ZN(new_n378));
  NOR3_X1   g192(.A1(new_n377), .A2(new_n378), .A3(G953), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n375), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n379), .A2(new_n369), .A3(new_n374), .ZN(new_n382));
  AOI21_X1  g196(.A(G902), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G478), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n384), .A2(KEYINPUT15), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n383), .B(new_n386), .ZN(new_n387));
  NOR3_X1   g201(.A1(new_n351), .A2(new_n356), .A3(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(G221), .B1(new_n377), .B2(G902), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT11), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n390), .B1(new_n358), .B2(G137), .ZN(new_n391));
  INV_X1    g205(.A(G137), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(KEYINPUT11), .A3(G134), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n358), .A2(G137), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n391), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G131), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n391), .A2(new_n393), .A3(new_n315), .A4(new_n394), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n265), .A2(new_n197), .A3(new_n200), .A4(new_n267), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n399), .A2(KEYINPUT10), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n265), .A2(KEYINPUT67), .A3(new_n267), .ZN(new_n401));
  AOI21_X1  g215(.A(KEYINPUT67), .B1(new_n265), .B2(new_n267), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n202), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n400), .B1(new_n403), .B2(KEYINPUT10), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n224), .A2(new_n247), .A3(new_n254), .A4(new_n259), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n405), .B1(new_n218), .B2(new_n221), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n398), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n400), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT67), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n268), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n265), .A2(KEYINPUT67), .A3(new_n267), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n201), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT10), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n408), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n398), .ZN(new_n415));
  INV_X1    g229(.A(new_n405), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n217), .A2(KEYINPUT80), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n220), .B1(new_n219), .B2(new_n216), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n414), .A2(new_n415), .A3(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(G110), .B(G140), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n309), .A2(G227), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n421), .B(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n407), .A2(new_n420), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n268), .A2(new_n201), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n399), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT12), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n427), .A2(new_n428), .A3(new_n398), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n428), .B1(new_n427), .B2(new_n398), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n424), .B1(new_n420), .B2(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n425), .A2(new_n432), .ZN(new_n433));
  OAI211_X1 g247(.A(KEYINPUT82), .B(G469), .C1(new_n433), .C2(G902), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT82), .ZN(new_n435));
  INV_X1    g249(.A(G469), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n436), .A2(new_n281), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n407), .A2(new_n420), .A3(new_n424), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n420), .A2(new_n431), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n439), .B1(new_n440), .B2(new_n424), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n435), .B(new_n438), .C1(new_n441), .C2(new_n436), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n434), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n420), .A2(new_n431), .A3(new_n424), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n424), .B1(new_n407), .B2(new_n420), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n444), .B1(new_n445), .B2(KEYINPUT83), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT83), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n440), .A2(new_n447), .A3(new_n424), .ZN(new_n448));
  AOI211_X1 g262(.A(G469), .B(G902), .C1(new_n446), .C2(new_n448), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n388), .B(new_n389), .C1(new_n443), .C2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n296), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT70), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n238), .A2(new_n239), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n245), .A2(new_n246), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n253), .B1(new_n455), .B2(new_n258), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n456), .A2(new_n398), .A3(KEYINPUT65), .A4(new_n247), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n358), .A2(G137), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n392), .A2(G134), .ZN(new_n459));
  OAI21_X1  g273(.A(G131), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n397), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(new_n267), .A3(new_n265), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n457), .A2(new_n462), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n247), .A2(new_n254), .A3(new_n259), .ZN(new_n464));
  AOI21_X1  g278(.A(KEYINPUT65), .B1(new_n464), .B2(new_n398), .ZN(new_n465));
  OAI211_X1 g279(.A(KEYINPUT69), .B(new_n454), .C1(new_n463), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n464), .A2(new_n398), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n461), .B1(new_n401), .B2(new_n402), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(new_n468), .A3(new_n453), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT65), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n471), .B1(new_n415), .B2(new_n260), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(new_n462), .A3(new_n457), .ZN(new_n473));
  AOI21_X1  g287(.A(KEYINPUT69), .B1(new_n473), .B2(new_n454), .ZN(new_n474));
  OAI21_X1  g288(.A(KEYINPUT28), .B1(new_n470), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT28), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n469), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n308), .A2(new_n309), .A3(G210), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n479), .B(KEYINPUT27), .ZN(new_n480));
  XNOR2_X1  g294(.A(KEYINPUT26), .B(G101), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n480), .B(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n482), .B(KEYINPUT68), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT30), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n484), .B1(new_n463), .B2(new_n465), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n467), .A2(new_n468), .A3(KEYINPUT30), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(new_n454), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(new_n469), .A3(new_n482), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT31), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n487), .A2(KEYINPUT31), .A3(new_n469), .A4(new_n482), .ZN(new_n491));
  AOI22_X1  g305(.A1(new_n478), .A2(new_n483), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(G472), .A2(G902), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n452), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n490), .A2(new_n491), .ZN(new_n496));
  INV_X1    g310(.A(new_n483), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n497), .B1(new_n475), .B2(new_n477), .ZN(new_n498));
  OAI211_X1 g312(.A(KEYINPUT70), .B(new_n493), .C1(new_n496), .C2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT32), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n495), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT71), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n487), .A2(new_n469), .ZN(new_n503));
  INV_X1    g317(.A(new_n482), .ZN(new_n504));
  AOI21_X1  g318(.A(KEYINPUT29), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n483), .B1(new_n476), .B2(new_n469), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n475), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n469), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n453), .B1(new_n467), .B2(new_n468), .ZN(new_n510));
  OAI21_X1  g324(.A(KEYINPUT28), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n482), .A2(KEYINPUT29), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n511), .A2(new_n477), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n281), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n502), .B(G472), .C1(new_n508), .C2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n514), .B1(new_n505), .B2(new_n507), .ZN(new_n516));
  INV_X1    g330(.A(G472), .ZN(new_n517));
  OAI21_X1  g331(.A(KEYINPUT71), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n478), .A2(new_n483), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n490), .A2(new_n491), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n522), .A2(KEYINPUT32), .A3(new_n493), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n501), .A2(new_n519), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n378), .B1(G234), .B2(new_n281), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT78), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n527), .A2(KEYINPUT25), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT74), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n266), .B(G119), .C1(KEYINPUT73), .C2(KEYINPUT23), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT23), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n531), .B1(new_n203), .B2(G128), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT73), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n533), .B1(new_n203), .B2(G128), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n530), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n529), .B1(new_n535), .B2(G110), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n266), .A2(G119), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n203), .A2(G128), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(G110), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(KEYINPUT24), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT24), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(G110), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT72), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n541), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n544), .B1(new_n541), .B2(new_n543), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n539), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n266), .A2(G119), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n533), .B(new_n537), .C1(new_n548), .C2(new_n531), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n549), .A2(KEYINPUT74), .A3(new_n540), .A4(new_n530), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n536), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n324), .A2(new_n305), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NOR3_X1   g367(.A1(new_n545), .A2(new_n546), .A3(new_n539), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n540), .B1(new_n549), .B2(new_n530), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n306), .ZN(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT22), .B(G137), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n309), .A2(G221), .A3(G234), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n558), .B(new_n559), .ZN(new_n560));
  AND4_X1   g374(.A1(KEYINPUT77), .A2(new_n553), .A3(new_n557), .A4(new_n560), .ZN(new_n561));
  AOI22_X1  g375(.A1(new_n551), .A2(new_n552), .B1(new_n556), .B2(new_n306), .ZN(new_n562));
  AOI21_X1  g376(.A(KEYINPUT77), .B1(new_n562), .B2(new_n560), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n553), .A2(new_n557), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n560), .B(KEYINPUT76), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n561), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n528), .B1(new_n567), .B2(G902), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n562), .A2(KEYINPUT77), .A3(new_n560), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n553), .A2(new_n557), .A3(new_n560), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT77), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  XOR2_X1   g386(.A(new_n560), .B(KEYINPUT76), .Z(new_n573));
  NOR2_X1   g387(.A1(new_n562), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n569), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n528), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(new_n281), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n526), .B1(new_n568), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n525), .A2(G902), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n451), .A2(new_n524), .A3(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(G101), .ZN(G3));
  NOR3_X1   g398(.A1(new_n293), .A2(new_n295), .A3(KEYINPUT89), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n280), .A2(new_n188), .A3(new_n292), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT89), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n187), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(KEYINPUT90), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n356), .ZN(new_n590));
  INV_X1    g404(.A(new_n383), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n591), .A2(KEYINPUT93), .A3(new_n384), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT93), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n593), .B1(new_n383), .B2(G478), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n382), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n379), .B1(new_n369), .B2(new_n374), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT91), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n598), .A2(KEYINPUT92), .A3(KEYINPUT33), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT92), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n381), .A2(new_n382), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n600), .B1(new_n601), .B2(KEYINPUT91), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n603), .B1(new_n601), .B2(new_n600), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n599), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n281), .A2(G478), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n595), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n351), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n280), .A2(new_n292), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n294), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n611), .A2(new_n587), .A3(new_n586), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT90), .ZN(new_n613));
  INV_X1    g427(.A(new_n187), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n614), .B1(new_n295), .B2(KEYINPUT89), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n612), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n589), .A2(new_n590), .A3(new_n609), .A4(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n389), .B1(new_n443), .B2(new_n449), .ZN(new_n618));
  INV_X1    g432(.A(new_n582), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(G472), .B1(new_n492), .B2(G902), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n495), .A2(new_n621), .A3(new_n499), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n617), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT95), .B(G104), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT94), .B(KEYINPUT34), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G6));
  NOR3_X1   g442(.A1(new_n585), .A2(KEYINPUT90), .A3(new_n588), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n613), .B1(new_n612), .B2(new_n615), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n351), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n387), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n631), .A2(new_n590), .A3(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n635), .A2(new_n623), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT35), .B(G107), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G9));
  AOI21_X1  g452(.A(KEYINPUT70), .B1(new_n522), .B2(new_n493), .ZN(new_n639));
  AOI211_X1 g453(.A(new_n452), .B(new_n494), .C1(new_n520), .C2(new_n521), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n567), .A2(G902), .A3(new_n528), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n576), .B1(new_n575), .B2(new_n281), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n525), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n565), .A2(KEYINPUT36), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(new_n564), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n579), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n641), .A2(KEYINPUT96), .A3(new_n621), .A4(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n495), .A2(new_n621), .A3(new_n499), .A4(new_n648), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT96), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n649), .A2(new_n451), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT37), .B(G110), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G12));
  INV_X1    g469(.A(new_n648), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n494), .B1(new_n520), .B2(new_n521), .ZN(new_n657));
  AOI22_X1  g471(.A1(new_n515), .A2(new_n518), .B1(KEYINPUT32), .B2(new_n657), .ZN(new_n658));
  AOI211_X1 g472(.A(new_n656), .B(new_n618), .C1(new_n658), .C2(new_n501), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT97), .B(G900), .Z(new_n660));
  AOI21_X1  g474(.A(new_n353), .B1(new_n354), .B2(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n633), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n659), .A2(new_n616), .A3(new_n589), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT98), .B(G128), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G30));
  NOR2_X1   g479(.A1(new_n293), .A2(new_n295), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n667));
  XOR2_X1   g481(.A(new_n666), .B(new_n667), .Z(new_n668));
  OAI21_X1  g482(.A(new_n483), .B1(new_n509), .B2(new_n510), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n488), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n517), .B1(new_n670), .B2(new_n281), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n671), .B1(new_n657), .B2(KEYINPUT32), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n501), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n387), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n632), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n676), .A2(new_n656), .A3(new_n187), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n668), .A2(new_n674), .A3(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n618), .ZN(new_n679));
  XOR2_X1   g493(.A(new_n661), .B(KEYINPUT39), .Z(new_n680));
  AND2_X1   g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(KEYINPUT40), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G143), .ZN(G45));
  NOR2_X1   g498(.A1(new_n608), .A2(new_n661), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n659), .A2(new_n616), .A3(new_n589), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G146), .ZN(G48));
  AOI21_X1  g501(.A(new_n619), .B1(new_n658), .B2(new_n501), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n446), .A2(new_n448), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n436), .B1(new_n689), .B2(new_n281), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n689), .A2(new_n436), .A3(new_n281), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n691), .A2(new_n389), .A3(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n688), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n617), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT41), .B(G113), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G15));
  AOI211_X1 g512(.A(new_n619), .B(new_n693), .C1(new_n658), .C2(new_n501), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n631), .A2(new_n590), .A3(new_n634), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G116), .ZN(G18));
  AND3_X1   g515(.A1(new_n524), .A2(new_n388), .A3(new_n648), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n631), .A2(new_n694), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G119), .ZN(G21));
  OAI21_X1  g518(.A(KEYINPUT100), .B1(new_n578), .B2(new_n581), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT100), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n644), .A2(new_n706), .A3(new_n580), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n497), .B1(new_n511), .B2(new_n477), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n493), .B1(new_n496), .B2(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n708), .A2(new_n621), .A3(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n690), .A2(new_n449), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(new_n389), .A3(new_n590), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n589), .A2(new_n714), .A3(new_n616), .A4(new_n676), .ZN(new_n715));
  XNOR2_X1  g529(.A(KEYINPUT101), .B(G122), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G24));
  INV_X1    g531(.A(new_n685), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n621), .A2(new_n648), .A3(new_n710), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n589), .A2(new_n616), .A3(new_n694), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G125), .ZN(G27));
  NOR3_X1   g536(.A1(new_n293), .A2(new_n295), .A3(new_n614), .ZN(new_n723));
  INV_X1    g537(.A(new_n389), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT103), .ZN(new_n725));
  OAI21_X1  g539(.A(KEYINPUT102), .B1(new_n425), .B2(new_n432), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT102), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n439), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n726), .A2(G469), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n438), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n725), .B1(new_n730), .B2(new_n449), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n692), .A2(KEYINPUT103), .A3(new_n438), .A4(new_n729), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n724), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n688), .A2(new_n685), .A3(new_n723), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(KEYINPUT104), .B(KEYINPUT42), .ZN(new_n735));
  INV_X1    g549(.A(new_n708), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n500), .B1(new_n492), .B2(new_n494), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT105), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n523), .A3(new_n738), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n739), .A2(new_n519), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n737), .A2(new_n523), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT105), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n736), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n685), .A2(KEYINPUT42), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n744), .A2(new_n733), .A3(new_n723), .ZN(new_n745));
  AOI22_X1  g559(.A1(new_n734), .A2(new_n735), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(new_n315), .ZN(G33));
  NAND4_X1  g561(.A1(new_n688), .A2(new_n662), .A3(new_n723), .A4(new_n733), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G134), .ZN(G36));
  OAI21_X1  g563(.A(G469), .B1(new_n433), .B2(KEYINPUT45), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n726), .A2(new_n728), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n750), .B1(new_n751), .B2(KEYINPUT45), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n752), .A2(new_n437), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n753), .A2(KEYINPUT46), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(KEYINPUT46), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(new_n692), .A3(new_n755), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n756), .A2(new_n389), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n680), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n632), .A2(new_n607), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(KEYINPUT43), .ZN(new_n761));
  OR3_X1    g575(.A1(new_n761), .A2(new_n622), .A3(new_n656), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT44), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n759), .A2(new_n723), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  XOR2_X1   g580(.A(KEYINPUT106), .B(G137), .Z(new_n767));
  XNOR2_X1  g581(.A(new_n766), .B(new_n767), .ZN(G39));
  OR2_X1    g582(.A1(new_n757), .A2(KEYINPUT47), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n757), .A2(KEYINPUT47), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(new_n723), .ZN(new_n772));
  NOR4_X1   g586(.A1(new_n524), .A2(new_n772), .A3(new_n582), .A4(new_n718), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G140), .ZN(G42));
  NOR3_X1   g589(.A1(new_n760), .A2(new_n614), .A3(new_n724), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT49), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n776), .B(new_n708), .C1(new_n777), .C2(new_n712), .ZN(new_n778));
  XOR2_X1   g592(.A(new_n778), .B(KEYINPUT107), .Z(new_n779));
  NAND2_X1  g593(.A1(new_n712), .A2(new_n777), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n779), .A2(new_n674), .A3(new_n668), .A4(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n353), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n761), .A2(new_n711), .A3(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n631), .A2(new_n783), .A3(new_n694), .ZN(new_n784));
  XOR2_X1   g598(.A(new_n784), .B(KEYINPUT116), .Z(new_n785));
  NOR2_X1   g599(.A1(new_n761), .A2(new_n782), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n772), .A2(new_n693), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n743), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(KEYINPUT48), .ZN(new_n789));
  XOR2_X1   g603(.A(new_n352), .B(KEYINPUT115), .Z(new_n790));
  AND4_X1   g604(.A1(new_n582), .A2(new_n787), .A3(new_n353), .A4(new_n674), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n790), .B1(new_n791), .B2(new_n609), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n785), .A2(new_n789), .A3(new_n792), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n690), .A2(new_n449), .A3(new_n389), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n723), .B(new_n783), .C1(new_n771), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n787), .A2(new_n786), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n796), .A2(new_n719), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n668), .A2(new_n783), .A3(new_n614), .A4(new_n694), .ZN(new_n798));
  NOR2_X1   g612(.A1(KEYINPUT112), .A2(KEYINPUT50), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n797), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n607), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n791), .A2(new_n632), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT113), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n795), .A2(new_n802), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n793), .B1(new_n807), .B2(KEYINPUT51), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n809));
  XNOR2_X1  g623(.A(KEYINPUT111), .B(KEYINPUT51), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n806), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n809), .B1(new_n806), .B2(new_n810), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n808), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n648), .A2(new_n661), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n673), .A2(new_n733), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n631), .A2(new_n676), .A3(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n816), .A2(new_n663), .A3(new_n686), .A4(new_n721), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT52), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n631), .B(new_n659), .C1(new_n662), .C2(new_n685), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT52), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n819), .A2(new_n820), .A3(new_n721), .A4(new_n816), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n296), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n356), .B1(new_n633), .B2(new_n608), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n823), .A2(new_n620), .A3(new_n622), .A4(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n653), .A2(new_n583), .A3(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT108), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n653), .A2(new_n583), .A3(KEYINPUT108), .A4(new_n825), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n631), .A2(new_n590), .A3(new_n609), .A4(new_n699), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(new_n700), .A3(new_n703), .A4(new_n715), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n656), .B1(new_n658), .B2(new_n501), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n351), .A2(new_n387), .A3(new_n661), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n611), .A2(new_n187), .A3(new_n586), .A4(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT109), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n666), .A2(KEYINPUT109), .A3(new_n187), .A4(new_n834), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n833), .A2(new_n679), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n720), .A2(new_n723), .A3(new_n733), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n748), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n524), .A2(new_n582), .A3(new_n733), .A4(new_n723), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n735), .B1(new_n842), .B2(new_n718), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n733), .A2(new_n723), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n742), .A2(new_n519), .A3(new_n739), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n844), .A2(new_n708), .A3(new_n845), .A4(new_n744), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n841), .A2(new_n847), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n830), .A2(new_n832), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n822), .A2(new_n849), .A3(KEYINPUT53), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n818), .A2(new_n821), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n748), .A2(new_n839), .A3(new_n840), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n746), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n828), .A2(new_n829), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n589), .A2(new_n616), .A3(new_n694), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n833), .A2(new_n388), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n715), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n858), .A2(new_n696), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n854), .A2(new_n855), .A3(new_n859), .A4(new_n700), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n851), .B1(new_n852), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n850), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n862), .A2(KEYINPUT54), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT110), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n862), .A2(KEYINPUT54), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n863), .A2(KEYINPUT110), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n813), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(G952), .A2(G953), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n781), .B1(new_n869), .B2(new_n870), .ZN(G75));
  NOR2_X1   g685(.A1(new_n309), .A2(G952), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(G210), .A2(G902), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n874), .B1(new_n850), .B2(new_n861), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n275), .B(KEYINPUT55), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT118), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n243), .A2(new_n244), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT117), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n877), .B(new_n879), .ZN(new_n880));
  OR2_X1    g694(.A1(new_n880), .A2(KEYINPUT56), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n873), .B1(new_n875), .B2(new_n881), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n875), .A2(KEYINPUT119), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT56), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n884), .B1(new_n875), .B2(KEYINPUT119), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n880), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT120), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI211_X1 g702(.A(KEYINPUT120), .B(new_n880), .C1(new_n883), .C2(new_n885), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n882), .B1(new_n888), .B2(new_n889), .ZN(G51));
  XNOR2_X1  g704(.A(new_n437), .B(KEYINPUT57), .ZN(new_n891));
  INV_X1    g705(.A(new_n866), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n891), .B1(new_n892), .B2(new_n863), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n689), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n862), .A2(G902), .A3(new_n752), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n872), .B1(new_n894), .B2(new_n895), .ZN(G54));
  NAND4_X1  g710(.A1(new_n862), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT121), .ZN(new_n898));
  INV_X1    g712(.A(new_n346), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n873), .B1(new_n897), .B2(new_n899), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n898), .B1(new_n897), .B2(new_n899), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(G60));
  INV_X1    g717(.A(new_n605), .ZN(new_n904));
  NAND2_X1  g718(.A1(G478), .A2(G902), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT59), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n904), .B(new_n906), .C1(new_n892), .C2(new_n863), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n873), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n867), .A2(new_n868), .A3(new_n906), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n908), .B1(new_n605), .B2(new_n909), .ZN(G63));
  INV_X1    g724(.A(KEYINPUT123), .ZN(new_n911));
  XNOR2_X1  g725(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n378), .A2(new_n281), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n912), .B(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n911), .B1(new_n862), .B2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(new_n914), .ZN(new_n916));
  AOI211_X1 g730(.A(KEYINPUT123), .B(new_n916), .C1(new_n850), .C2(new_n861), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n646), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT53), .B1(new_n822), .B2(new_n849), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n852), .A2(new_n860), .A3(new_n851), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n914), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(KEYINPUT123), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n862), .A2(new_n911), .A3(new_n914), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n922), .A2(new_n567), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n918), .A2(new_n924), .A3(new_n873), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT61), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n918), .A2(new_n924), .A3(KEYINPUT61), .A4(new_n873), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(G66));
  OAI21_X1  g743(.A(G953), .B1(new_n355), .B2(new_n273), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n830), .A2(new_n832), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n930), .B1(new_n931), .B2(G953), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n879), .B1(G898), .B2(new_n309), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT124), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n932), .B(new_n934), .ZN(G69));
  AOI21_X1  g749(.A(new_n309), .B1(G227), .B2(G900), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n759), .A2(new_n631), .A3(new_n676), .A4(new_n743), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n774), .A2(new_n748), .A3(new_n766), .A4(new_n937), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n819), .A2(new_n721), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n847), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n938), .A2(G953), .A3(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n485), .A2(new_n486), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT125), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(new_n341), .ZN(new_n945));
  NAND2_X1  g759(.A1(G900), .A2(G953), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n942), .A2(KEYINPUT127), .A3(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT127), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(new_n941), .B2(new_n947), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n633), .A2(new_n608), .ZN(new_n953));
  AND4_X1   g767(.A1(new_n688), .A2(new_n681), .A3(new_n723), .A4(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n774), .A2(new_n766), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n939), .A2(new_n683), .ZN(new_n957));
  OR2_X1    g771(.A1(new_n957), .A2(KEYINPUT62), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(KEYINPUT62), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n956), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n945), .B1(new_n960), .B2(new_n309), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n936), .B1(new_n952), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n936), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n963), .B1(new_n941), .B2(new_n947), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n964), .A2(new_n961), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n965), .A2(KEYINPUT126), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT126), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n964), .A2(new_n961), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n962), .B1(new_n966), .B2(new_n968), .ZN(G72));
  NAND2_X1  g783(.A1(new_n503), .A2(new_n482), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n956), .A2(new_n931), .A3(new_n958), .A4(new_n959), .ZN(new_n971));
  NAND2_X1  g785(.A1(G472), .A2(G902), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT63), .Z(new_n973));
  AOI21_X1  g787(.A(new_n970), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n973), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n938), .A2(new_n940), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n975), .B1(new_n976), .B2(new_n931), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n487), .A2(new_n469), .A3(new_n504), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n873), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n503), .A2(new_n504), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n975), .B1(new_n980), .B2(new_n488), .ZN(new_n981));
  AOI211_X1 g795(.A(new_n974), .B(new_n979), .C1(new_n862), .C2(new_n981), .ZN(G57));
endmodule


