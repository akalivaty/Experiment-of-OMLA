

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770;

  INV_X2 U377 ( .A(G953), .ZN(n763) );
  INV_X2 U378 ( .A(n503), .ZN(n516) );
  XNOR2_X2 U379 ( .A(n578), .B(KEYINPUT0), .ZN(n605) );
  XNOR2_X2 U380 ( .A(n502), .B(KEYINPUT42), .ZN(n770) );
  NOR2_X2 U381 ( .A1(n662), .A2(n529), .ZN(n502) );
  XNOR2_X2 U382 ( .A(n483), .B(n386), .ZN(n756) );
  XNOR2_X2 U383 ( .A(n443), .B(n442), .ZN(n483) );
  AND2_X2 U384 ( .A1(n713), .A2(n624), .ZN(n419) );
  INV_X1 U385 ( .A(KEYINPUT74), .ZN(n359) );
  NAND2_X1 U386 ( .A1(n394), .A2(n392), .ZN(n699) );
  AND2_X1 U387 ( .A1(n397), .A2(n395), .ZN(n394) );
  NAND2_X1 U388 ( .A1(n393), .A2(KEYINPUT118), .ZN(n392) );
  AND2_X1 U389 ( .A1(n402), .A2(n387), .ZN(n631) );
  XNOR2_X1 U390 ( .A(n360), .B(n359), .ZN(n558) );
  NOR2_X1 U391 ( .A1(n597), .A2(n654), .ZN(n600) );
  XNOR2_X1 U392 ( .A(n596), .B(KEYINPUT35), .ZN(n654) );
  AND2_X1 U393 ( .A1(n553), .A2(n727), .ZN(n557) );
  XNOR2_X1 U394 ( .A(n581), .B(n582), .ZN(n373) );
  XNOR2_X1 U395 ( .A(n531), .B(KEYINPUT38), .ZN(n510) );
  XNOR2_X1 U396 ( .A(n470), .B(n469), .ZN(n503) );
  OR2_X1 U397 ( .A1(n742), .A2(G902), .ZN(n501) );
  XNOR2_X1 U398 ( .A(n500), .B(n389), .ZN(n640) );
  XNOR2_X1 U399 ( .A(n756), .B(G146), .ZN(n500) );
  XNOR2_X1 U400 ( .A(n411), .B(G122), .ZN(n441) );
  XNOR2_X1 U401 ( .A(n372), .B(KEYINPUT3), .ZN(n487) );
  XOR2_X1 U402 ( .A(G119), .B(G110), .Z(n462) );
  XNOR2_X1 U403 ( .A(G113), .B(G101), .ZN(n372) );
  BUF_X1 U404 ( .A(n606), .Z(n355) );
  INV_X1 U405 ( .A(n695), .ZN(n356) );
  INV_X1 U406 ( .A(n687), .ZN(n357) );
  XNOR2_X1 U407 ( .A(n592), .B(KEYINPUT33), .ZN(n686) );
  XNOR2_X1 U408 ( .A(n358), .B(n415), .ZN(n404) );
  XOR2_X1 U409 ( .A(n430), .B(n443), .Z(n358) );
  NAND2_X1 U410 ( .A1(n557), .A2(n556), .ZN(n360) );
  XNOR2_X1 U411 ( .A(n374), .B(n391), .ZN(n535) );
  NAND2_X1 U412 ( .A1(n362), .A2(n375), .ZN(n374) );
  NOR2_X2 U413 ( .A1(n682), .A2(n680), .ZN(n451) );
  XNOR2_X2 U414 ( .A(n422), .B(n421), .ZN(n682) );
  XNOR2_X1 U415 ( .A(n482), .B(KEYINPUT70), .ZN(n386) );
  NOR2_X1 U416 ( .A1(n550), .A2(n530), .ZN(n380) );
  XNOR2_X1 U417 ( .A(n493), .B(n492), .ZN(n375) );
  AND2_X1 U418 ( .A1(n503), .A2(n520), .ZN(n491) );
  AND2_X1 U419 ( .A1(n534), .A2(n369), .ZN(n578) );
  NAND2_X1 U420 ( .A1(n410), .A2(n409), .ZN(n411) );
  XNOR2_X1 U421 ( .A(KEYINPUT94), .B(G110), .ZN(n497) );
  XNOR2_X1 U422 ( .A(G107), .B(G101), .ZN(n495) );
  NOR2_X1 U423 ( .A1(n399), .A2(KEYINPUT118), .ZN(n398) );
  NAND2_X1 U424 ( .A1(n403), .A2(n402), .ZN(n401) );
  NOR2_X1 U425 ( .A1(n522), .A2(n521), .ZN(n523) );
  INV_X1 U426 ( .A(n668), .ZN(n381) );
  NAND2_X1 U427 ( .A1(n524), .A2(n378), .ZN(n377) );
  NOR2_X1 U428 ( .A1(n379), .A2(KEYINPUT36), .ZN(n378) );
  INV_X1 U429 ( .A(n380), .ZN(n379) );
  XNOR2_X1 U430 ( .A(n561), .B(n560), .ZN(n627) );
  XNOR2_X1 U431 ( .A(n453), .B(n452), .ZN(n757) );
  XNOR2_X1 U432 ( .A(G140), .B(G143), .ZN(n423) );
  INV_X1 U433 ( .A(KEYINPUT113), .ZN(n421) );
  XNOR2_X1 U434 ( .A(n390), .B(n487), .ZN(n389) );
  XNOR2_X1 U435 ( .A(n486), .B(n366), .ZN(n390) );
  NAND2_X1 U436 ( .A1(n524), .A2(n679), .ZN(n566) );
  XNOR2_X1 U437 ( .A(n506), .B(n505), .ZN(n508) );
  INV_X1 U438 ( .A(KEYINPUT30), .ZN(n505) );
  INV_X1 U439 ( .A(KEYINPUT112), .ZN(n391) );
  AND2_X1 U440 ( .A1(n373), .A2(n668), .ZN(n604) );
  XNOR2_X1 U441 ( .A(n413), .B(n412), .ZN(n748) );
  XNOR2_X1 U442 ( .A(n500), .B(n383), .ZN(n742) );
  XNOR2_X1 U443 ( .A(n385), .B(n384), .ZN(n383) );
  XNOR2_X1 U444 ( .A(n499), .B(n494), .ZN(n385) );
  NOR2_X1 U445 ( .A1(n396), .A2(G953), .ZN(n395) );
  NOR2_X1 U446 ( .A1(n363), .A2(n400), .ZN(n396) );
  NOR2_X1 U447 ( .A1(n376), .A2(n365), .ZN(n734) );
  NAND2_X1 U448 ( .A1(n377), .A2(n368), .ZN(n376) );
  XNOR2_X1 U449 ( .A(n388), .B(n370), .ZN(n595) );
  XOR2_X1 U450 ( .A(n404), .B(n416), .Z(n361) );
  XOR2_X1 U451 ( .A(n525), .B(KEYINPUT111), .Z(n362) );
  AND2_X1 U452 ( .A1(n697), .A2(n696), .ZN(n363) );
  OR2_X1 U453 ( .A1(n572), .A2(n737), .ZN(n364) );
  NOR2_X1 U454 ( .A1(n524), .A2(n382), .ZN(n365) );
  AND2_X1 U455 ( .A1(n488), .A2(G210), .ZN(n366) );
  OR2_X1 U456 ( .A1(n380), .A2(n382), .ZN(n367) );
  AND2_X1 U457 ( .A1(n381), .A2(n367), .ZN(n368) );
  AND2_X1 U458 ( .A1(n577), .A2(n576), .ZN(n369) );
  XOR2_X1 U459 ( .A(KEYINPUT78), .B(KEYINPUT34), .Z(n370) );
  XOR2_X1 U460 ( .A(n532), .B(KEYINPUT19), .Z(n371) );
  INV_X1 U461 ( .A(KEYINPUT36), .ZN(n382) );
  XNOR2_X1 U462 ( .A(n361), .B(n748), .ZN(n713) );
  INV_X1 U463 ( .A(KEYINPUT118), .ZN(n400) );
  XNOR2_X1 U464 ( .A(n533), .B(n371), .ZN(n534) );
  NAND2_X1 U465 ( .A1(n373), .A2(n585), .ZN(n587) );
  NAND2_X1 U466 ( .A1(n535), .A2(n534), .ZN(n537) );
  XNOR2_X2 U467 ( .A(n430), .B(n429), .ZN(n453) );
  NOR2_X1 U468 ( .A1(n770), .A2(n769), .ZN(n515) );
  INV_X1 U469 ( .A(n667), .ZN(n589) );
  NOR2_X1 U470 ( .A1(n528), .A2(n527), .ZN(n559) );
  XNOR2_X1 U471 ( .A(n496), .B(n495), .ZN(n384) );
  INV_X1 U472 ( .A(n624), .ZN(n387) );
  NAND2_X1 U473 ( .A1(n623), .A2(n657), .ZN(n402) );
  NAND2_X1 U474 ( .A1(n686), .A2(n605), .ZN(n388) );
  INV_X1 U475 ( .A(n535), .ZN(n529) );
  INV_X1 U476 ( .A(n401), .ZN(n393) );
  NAND2_X1 U477 ( .A1(n401), .A2(n398), .ZN(n397) );
  INV_X1 U478 ( .A(n363), .ZN(n399) );
  INV_X1 U479 ( .A(n661), .ZN(n403) );
  XNOR2_X1 U480 ( .A(n734), .B(n526), .ZN(n527) );
  NOR2_X2 U481 ( .A1(n606), .A2(n509), .ZN(n552) );
  INV_X1 U482 ( .A(KEYINPUT89), .ZN(n526) );
  XNOR2_X1 U483 ( .A(n414), .B(KEYINPUT17), .ZN(n415) );
  INV_X1 U484 ( .A(KEYINPUT28), .ZN(n492) );
  BUF_X1 U485 ( .A(n700), .Z(n701) );
  NAND2_X1 U486 ( .A1(n508), .A2(n507), .ZN(n509) );
  INV_X1 U487 ( .A(KEYINPUT63), .ZN(n644) );
  INV_X1 U488 ( .A(KEYINPUT91), .ZN(n405) );
  XNOR2_X1 U489 ( .A(n405), .B(G104), .ZN(n496) );
  XNOR2_X1 U490 ( .A(n462), .B(n496), .ZN(n406) );
  XNOR2_X1 U491 ( .A(n406), .B(n487), .ZN(n413) );
  INV_X1 U492 ( .A(G107), .ZN(n407) );
  NAND2_X1 U493 ( .A1(G116), .A2(n407), .ZN(n410) );
  INV_X1 U494 ( .A(G116), .ZN(n408) );
  NAND2_X1 U495 ( .A1(n408), .A2(G107), .ZN(n409) );
  XNOR2_X1 U496 ( .A(KEYINPUT16), .B(n441), .ZN(n412) );
  XNOR2_X2 U497 ( .A(G146), .B(G125), .ZN(n430) );
  XNOR2_X2 U498 ( .A(G143), .B(G128), .ZN(n443) );
  XOR2_X1 U499 ( .A(KEYINPUT18), .B(KEYINPUT4), .Z(n414) );
  NAND2_X1 U500 ( .A1(G224), .A2(n763), .ZN(n416) );
  XNOR2_X1 U501 ( .A(G902), .B(KEYINPUT90), .ZN(n417) );
  XNOR2_X1 U502 ( .A(n417), .B(KEYINPUT15), .ZN(n624) );
  OR2_X1 U503 ( .A1(G902), .A2(G237), .ZN(n420) );
  AND2_X1 U504 ( .A1(G210), .A2(n420), .ZN(n418) );
  XNOR2_X2 U505 ( .A(n419), .B(n418), .ZN(n531) );
  NAND2_X1 U506 ( .A1(G214), .A2(n420), .ZN(n679) );
  NAND2_X1 U507 ( .A1(n510), .A2(n679), .ZN(n422) );
  XOR2_X1 U508 ( .A(G113), .B(G131), .Z(n424) );
  XNOR2_X1 U509 ( .A(n424), .B(n423), .ZN(n428) );
  XOR2_X1 U510 ( .A(KEYINPUT11), .B(KEYINPUT101), .Z(n426) );
  XNOR2_X1 U511 ( .A(G104), .B(G122), .ZN(n425) );
  XNOR2_X1 U512 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U513 ( .A(n428), .B(n427), .Z(n435) );
  XNOR2_X2 U514 ( .A(KEYINPUT69), .B(KEYINPUT10), .ZN(n429) );
  XOR2_X1 U515 ( .A(KEYINPUT12), .B(KEYINPUT100), .Z(n432) );
  NOR2_X1 U516 ( .A1(G953), .A2(G237), .ZN(n488) );
  NAND2_X1 U517 ( .A1(G214), .A2(n488), .ZN(n431) );
  XNOR2_X1 U518 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U519 ( .A(n453), .B(n433), .ZN(n434) );
  XNOR2_X1 U520 ( .A(n435), .B(n434), .ZN(n706) );
  INV_X1 U521 ( .A(G902), .ZN(n489) );
  NAND2_X1 U522 ( .A1(n706), .A2(n489), .ZN(n437) );
  XNOR2_X1 U523 ( .A(KEYINPUT13), .B(G475), .ZN(n436) );
  XNOR2_X1 U524 ( .A(n437), .B(n436), .ZN(n549) );
  NAND2_X1 U525 ( .A1(G234), .A2(n763), .ZN(n439) );
  XOR2_X1 U526 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n438) );
  XNOR2_X1 U527 ( .A(n439), .B(n438), .ZN(n454) );
  NAND2_X1 U528 ( .A1(n454), .A2(G217), .ZN(n440) );
  XNOR2_X1 U529 ( .A(n441), .B(n440), .ZN(n448) );
  INV_X1 U530 ( .A(G134), .ZN(n442) );
  XOR2_X1 U531 ( .A(KEYINPUT102), .B(KEYINPUT7), .Z(n445) );
  XNOR2_X1 U532 ( .A(KEYINPUT103), .B(KEYINPUT9), .ZN(n444) );
  XNOR2_X1 U533 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U534 ( .A(n483), .B(n446), .ZN(n447) );
  XNOR2_X1 U535 ( .A(n448), .B(n447), .ZN(n634) );
  NOR2_X1 U536 ( .A1(n634), .A2(G902), .ZN(n450) );
  XNOR2_X1 U537 ( .A(KEYINPUT104), .B(G478), .ZN(n449) );
  XNOR2_X1 U538 ( .A(n450), .B(n449), .ZN(n548) );
  NAND2_X1 U539 ( .A1(n549), .A2(n548), .ZN(n680) );
  XNOR2_X1 U540 ( .A(n451), .B(KEYINPUT41), .ZN(n662) );
  XNOR2_X1 U541 ( .A(G140), .B(G137), .ZN(n498) );
  INV_X1 U542 ( .A(n498), .ZN(n452) );
  NAND2_X1 U543 ( .A1(n454), .A2(G221), .ZN(n455) );
  XNOR2_X1 U544 ( .A(n757), .B(n455), .ZN(n464) );
  XNOR2_X1 U545 ( .A(KEYINPUT24), .B(KEYINPUT96), .ZN(n457) );
  XNOR2_X1 U546 ( .A(KEYINPUT97), .B(KEYINPUT77), .ZN(n456) );
  XNOR2_X1 U547 ( .A(n457), .B(n456), .ZN(n460) );
  XNOR2_X1 U548 ( .A(G128), .B(KEYINPUT23), .ZN(n458) );
  XNOR2_X1 U549 ( .A(n458), .B(KEYINPUT95), .ZN(n459) );
  XNOR2_X1 U550 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U551 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U552 ( .A(n464), .B(n463), .ZN(n700) );
  OR2_X2 U553 ( .A1(n700), .A2(G902), .ZN(n470) );
  NAND2_X1 U554 ( .A1(n624), .A2(G234), .ZN(n466) );
  INV_X1 U555 ( .A(KEYINPUT20), .ZN(n465) );
  XNOR2_X1 U556 ( .A(n466), .B(n465), .ZN(n479) );
  INV_X1 U557 ( .A(G217), .ZN(n467) );
  OR2_X1 U558 ( .A1(n479), .A2(n467), .ZN(n468) );
  XNOR2_X1 U559 ( .A(n468), .B(KEYINPUT25), .ZN(n469) );
  XOR2_X1 U560 ( .A(KEYINPUT92), .B(KEYINPUT14), .Z(n472) );
  NAND2_X1 U561 ( .A1(G237), .A2(G234), .ZN(n471) );
  XNOR2_X1 U562 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U563 ( .A(KEYINPUT76), .B(n473), .ZN(n693) );
  INV_X1 U564 ( .A(n693), .ZN(n577) );
  NOR2_X1 U565 ( .A1(G900), .A2(n763), .ZN(n474) );
  NAND2_X1 U566 ( .A1(n474), .A2(G902), .ZN(n475) );
  NAND2_X1 U567 ( .A1(G952), .A2(n763), .ZN(n574) );
  NAND2_X1 U568 ( .A1(n475), .A2(n574), .ZN(n476) );
  NAND2_X1 U569 ( .A1(n577), .A2(n476), .ZN(n477) );
  XNOR2_X1 U570 ( .A(n477), .B(KEYINPUT81), .ZN(n507) );
  INV_X1 U571 ( .A(G221), .ZN(n478) );
  OR2_X1 U572 ( .A1(n479), .A2(n478), .ZN(n481) );
  INV_X1 U573 ( .A(KEYINPUT21), .ZN(n480) );
  XNOR2_X1 U574 ( .A(n481), .B(n480), .ZN(n664) );
  AND2_X1 U575 ( .A1(n507), .A2(n664), .ZN(n520) );
  XNOR2_X1 U576 ( .A(KEYINPUT4), .B(G131), .ZN(n482) );
  XOR2_X1 U577 ( .A(G116), .B(KEYINPUT5), .Z(n485) );
  XNOR2_X1 U578 ( .A(G137), .B(G119), .ZN(n484) );
  XNOR2_X1 U579 ( .A(n485), .B(n484), .ZN(n486) );
  NAND2_X1 U580 ( .A1(n640), .A2(n489), .ZN(n490) );
  XNOR2_X2 U581 ( .A(n490), .B(G472), .ZN(n519) );
  NAND2_X1 U582 ( .A1(n491), .A2(n519), .ZN(n493) );
  NAND2_X1 U583 ( .A1(n763), .A2(G227), .ZN(n494) );
  XNOR2_X1 U584 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X2 U585 ( .A(n501), .B(G469), .ZN(n525) );
  INV_X1 U586 ( .A(n548), .ZN(n538) );
  OR2_X1 U587 ( .A1(n549), .A2(n538), .ZN(n728) );
  INV_X1 U588 ( .A(n728), .ZN(n646) );
  NAND2_X1 U589 ( .A1(n516), .A2(n664), .ZN(n667) );
  NAND2_X1 U590 ( .A1(n589), .A2(n525), .ZN(n504) );
  XNOR2_X1 U591 ( .A(n504), .B(KEYINPUT98), .ZN(n606) );
  NAND2_X1 U592 ( .A1(n519), .A2(n679), .ZN(n506) );
  NAND2_X1 U593 ( .A1(n552), .A2(n510), .ZN(n512) );
  XOR2_X1 U594 ( .A(KEYINPUT73), .B(KEYINPUT39), .Z(n511) );
  XNOR2_X1 U595 ( .A(n512), .B(n511), .ZN(n564) );
  NAND2_X1 U596 ( .A1(n646), .A2(n564), .ZN(n513) );
  XOR2_X1 U597 ( .A(KEYINPUT40), .B(n513), .Z(n769) );
  INV_X1 U598 ( .A(KEYINPUT46), .ZN(n514) );
  XNOR2_X1 U599 ( .A(n515), .B(n514), .ZN(n528) );
  INV_X1 U600 ( .A(n516), .ZN(n601) );
  INV_X1 U601 ( .A(n601), .ZN(n665) );
  INV_X1 U602 ( .A(KEYINPUT106), .ZN(n517) );
  XNOR2_X1 U603 ( .A(n517), .B(KEYINPUT6), .ZN(n518) );
  XNOR2_X1 U604 ( .A(n519), .B(n518), .ZN(n602) );
  NAND2_X1 U605 ( .A1(n601), .A2(n602), .ZN(n522) );
  NAND2_X1 U606 ( .A1(n646), .A2(n520), .ZN(n521) );
  XNOR2_X1 U607 ( .A(n523), .B(KEYINPUT108), .ZN(n524) );
  INV_X1 U608 ( .A(n531), .ZN(n570) );
  INV_X1 U609 ( .A(n570), .ZN(n550) );
  XNOR2_X1 U610 ( .A(n525), .B(KEYINPUT1), .ZN(n590) );
  INV_X1 U611 ( .A(n590), .ZN(n668) );
  INV_X1 U612 ( .A(n679), .ZN(n530) );
  NOR2_X1 U613 ( .A1(n531), .A2(n530), .ZN(n533) );
  INV_X1 U614 ( .A(KEYINPUT67), .ZN(n532) );
  INV_X1 U615 ( .A(KEYINPUT80), .ZN(n536) );
  XNOR2_X2 U616 ( .A(n537), .B(n536), .ZN(n649) );
  NAND2_X1 U617 ( .A1(n549), .A2(n538), .ZN(n732) );
  INV_X1 U618 ( .A(KEYINPUT105), .ZN(n539) );
  XNOR2_X1 U619 ( .A(n732), .B(n539), .ZN(n562) );
  AND2_X1 U620 ( .A1(n562), .A2(n728), .ZN(n683) );
  INV_X1 U621 ( .A(n683), .ZN(n612) );
  INV_X1 U622 ( .A(KEYINPUT85), .ZN(n540) );
  AND2_X1 U623 ( .A1(n612), .A2(n540), .ZN(n541) );
  NAND2_X1 U624 ( .A1(n649), .A2(n541), .ZN(n543) );
  OR2_X1 U625 ( .A1(KEYINPUT85), .A2(KEYINPUT47), .ZN(n542) );
  AND2_X1 U626 ( .A1(n543), .A2(n542), .ZN(n547) );
  NAND2_X1 U627 ( .A1(KEYINPUT85), .A2(KEYINPUT47), .ZN(n544) );
  NOR2_X1 U628 ( .A1(n612), .A2(n544), .ZN(n545) );
  NAND2_X1 U629 ( .A1(n649), .A2(n545), .ZN(n546) );
  NAND2_X1 U630 ( .A1(n547), .A2(n546), .ZN(n553) );
  OR2_X1 U631 ( .A1(n549), .A2(n548), .ZN(n593) );
  NOR2_X1 U632 ( .A1(n550), .A2(n593), .ZN(n551) );
  NAND2_X1 U633 ( .A1(n552), .A2(n551), .ZN(n727) );
  NOR2_X1 U634 ( .A1(n683), .A2(KEYINPUT47), .ZN(n554) );
  AND2_X1 U635 ( .A1(n649), .A2(n554), .ZN(n555) );
  XNOR2_X1 U636 ( .A(KEYINPUT75), .B(n555), .ZN(n556) );
  NAND2_X1 U637 ( .A1(n559), .A2(n558), .ZN(n561) );
  XOR2_X1 U638 ( .A(KEYINPUT71), .B(KEYINPUT48), .Z(n560) );
  INV_X1 U639 ( .A(n562), .ZN(n563) );
  NAND2_X1 U640 ( .A1(n564), .A2(n563), .ZN(n736) );
  NAND2_X1 U641 ( .A1(n736), .A2(KEYINPUT2), .ZN(n565) );
  XNOR2_X1 U642 ( .A(n565), .B(KEYINPUT82), .ZN(n572) );
  XNOR2_X1 U643 ( .A(n566), .B(KEYINPUT109), .ZN(n567) );
  NAND2_X1 U644 ( .A1(n567), .A2(n668), .ZN(n569) );
  XOR2_X1 U645 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n568) );
  XNOR2_X1 U646 ( .A(n569), .B(n568), .ZN(n571) );
  NOR2_X1 U647 ( .A1(n571), .A2(n570), .ZN(n737) );
  NOR2_X1 U648 ( .A1(n627), .A2(n364), .ZN(n623) );
  XOR2_X1 U649 ( .A(KEYINPUT66), .B(KEYINPUT22), .Z(n582) );
  NOR2_X1 U650 ( .A1(G898), .A2(n763), .ZN(n573) );
  XOR2_X1 U651 ( .A(KEYINPUT93), .B(n573), .Z(n747) );
  NAND2_X1 U652 ( .A1(n747), .A2(G902), .ZN(n575) );
  NAND2_X1 U653 ( .A1(n575), .A2(n574), .ZN(n576) );
  INV_X1 U654 ( .A(n680), .ZN(n579) );
  AND2_X1 U655 ( .A1(n664), .A2(n579), .ZN(n580) );
  NAND2_X1 U656 ( .A1(n605), .A2(n580), .ZN(n581) );
  XNOR2_X1 U657 ( .A(KEYINPUT79), .B(n602), .ZN(n584) );
  AND2_X1 U658 ( .A1(n590), .A2(n601), .ZN(n583) );
  AND2_X1 U659 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U660 ( .A(KEYINPUT65), .B(KEYINPUT32), .Z(n586) );
  XNOR2_X1 U661 ( .A(n587), .B(n586), .ZN(n768) );
  NOR2_X1 U662 ( .A1(n519), .A2(n665), .ZN(n588) );
  NAND2_X1 U663 ( .A1(n604), .A2(n588), .ZN(n653) );
  NAND2_X1 U664 ( .A1(n768), .A2(n653), .ZN(n597) );
  NAND2_X1 U665 ( .A1(n590), .A2(n589), .ZN(n609) );
  XNOR2_X1 U666 ( .A(n609), .B(KEYINPUT107), .ZN(n591) );
  NAND2_X1 U667 ( .A1(n591), .A2(n602), .ZN(n592) );
  INV_X1 U668 ( .A(n593), .ZN(n594) );
  NAND2_X1 U669 ( .A1(n595), .A2(n594), .ZN(n596) );
  INV_X1 U670 ( .A(KEYINPUT44), .ZN(n598) );
  NAND2_X1 U671 ( .A1(n598), .A2(KEYINPUT72), .ZN(n599) );
  XNOR2_X1 U672 ( .A(n600), .B(n599), .ZN(n619) );
  NOR2_X1 U673 ( .A1(n602), .A2(n601), .ZN(n603) );
  NAND2_X1 U674 ( .A1(n604), .A2(n603), .ZN(n652) );
  INV_X1 U675 ( .A(n605), .ZN(n610) );
  NOR2_X1 U676 ( .A1(n355), .A2(n610), .ZN(n607) );
  INV_X1 U677 ( .A(n519), .ZN(n670) );
  AND2_X1 U678 ( .A1(n607), .A2(n670), .ZN(n608) );
  XNOR2_X1 U679 ( .A(n608), .B(KEYINPUT99), .ZN(n724) );
  OR2_X1 U680 ( .A1(n609), .A2(n670), .ZN(n663) );
  NOR2_X1 U681 ( .A1(n610), .A2(n663), .ZN(n611) );
  XNOR2_X1 U682 ( .A(KEYINPUT31), .B(n611), .ZN(n731) );
  NAND2_X1 U683 ( .A1(n724), .A2(n731), .ZN(n613) );
  NAND2_X1 U684 ( .A1(n613), .A2(n612), .ZN(n616) );
  INV_X1 U685 ( .A(KEYINPUT72), .ZN(n614) );
  NAND2_X1 U686 ( .A1(n614), .A2(KEYINPUT44), .ZN(n615) );
  AND2_X1 U687 ( .A1(n616), .A2(n615), .ZN(n617) );
  AND2_X1 U688 ( .A1(n652), .A2(n617), .ZN(n618) );
  NAND2_X1 U689 ( .A1(n619), .A2(n618), .ZN(n622) );
  INV_X1 U690 ( .A(KEYINPUT87), .ZN(n620) );
  XNOR2_X1 U691 ( .A(n620), .B(KEYINPUT45), .ZN(n621) );
  XNOR2_X2 U692 ( .A(n622), .B(n621), .ZN(n657) );
  INV_X1 U693 ( .A(n737), .ZN(n625) );
  NAND2_X1 U694 ( .A1(n625), .A2(n736), .ZN(n626) );
  NOR2_X2 U695 ( .A1(n627), .A2(n626), .ZN(n655) );
  BUF_X2 U696 ( .A(n655), .Z(n762) );
  NAND2_X1 U697 ( .A1(n762), .A2(n657), .ZN(n629) );
  INV_X1 U698 ( .A(KEYINPUT2), .ZN(n628) );
  NAND2_X1 U699 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U700 ( .A1(n630), .A2(n631), .ZN(n633) );
  INV_X1 U701 ( .A(KEYINPUT64), .ZN(n632) );
  XNOR2_X2 U702 ( .A(n633), .B(n632), .ZN(n712) );
  NAND2_X1 U703 ( .A1(n712), .A2(G478), .ZN(n635) );
  XNOR2_X1 U704 ( .A(n635), .B(n634), .ZN(n637) );
  INV_X1 U705 ( .A(G952), .ZN(n636) );
  AND2_X1 U706 ( .A1(n636), .A2(G953), .ZN(n746) );
  NOR2_X2 U707 ( .A1(n637), .A2(n746), .ZN(n639) );
  INV_X1 U708 ( .A(KEYINPUT123), .ZN(n638) );
  XNOR2_X1 U709 ( .A(n639), .B(n638), .ZN(G63) );
  NAND2_X1 U710 ( .A1(n712), .A2(G472), .ZN(n642) );
  XOR2_X1 U711 ( .A(KEYINPUT62), .B(n640), .Z(n641) );
  XNOR2_X1 U712 ( .A(n642), .B(n641), .ZN(n643) );
  NOR2_X2 U713 ( .A1(n643), .A2(n746), .ZN(n645) );
  XNOR2_X1 U714 ( .A(n645), .B(n644), .ZN(G57) );
  NAND2_X1 U715 ( .A1(n649), .A2(n646), .ZN(n647) );
  XNOR2_X1 U716 ( .A(n647), .B(G146), .ZN(G48) );
  INV_X1 U717 ( .A(n732), .ZN(n648) );
  NAND2_X1 U718 ( .A1(n649), .A2(n648), .ZN(n651) );
  XOR2_X1 U719 ( .A(G128), .B(KEYINPUT29), .Z(n650) );
  XNOR2_X1 U720 ( .A(n651), .B(n650), .ZN(G30) );
  XNOR2_X1 U721 ( .A(n652), .B(G101), .ZN(G3) );
  XNOR2_X1 U722 ( .A(n653), .B(G110), .ZN(G12) );
  XOR2_X1 U723 ( .A(G122), .B(n654), .Z(G24) );
  NOR2_X1 U724 ( .A1(n655), .A2(KEYINPUT2), .ZN(n656) );
  XNOR2_X1 U725 ( .A(n656), .B(KEYINPUT86), .ZN(n659) );
  NOR2_X1 U726 ( .A1(n657), .A2(KEYINPUT2), .ZN(n658) );
  NOR2_X1 U727 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U728 ( .A(n660), .B(KEYINPUT83), .ZN(n661) );
  INV_X1 U729 ( .A(n663), .ZN(n675) );
  NOR2_X1 U730 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U731 ( .A(KEYINPUT49), .B(n666), .Z(n673) );
  NAND2_X1 U732 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U733 ( .A(KEYINPUT50), .B(n669), .ZN(n671) );
  NAND2_X1 U734 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U735 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U736 ( .A1(n675), .A2(n674), .ZN(n676) );
  XOR2_X1 U737 ( .A(KEYINPUT51), .B(n676), .Z(n677) );
  NOR2_X1 U738 ( .A1(n356), .A2(n677), .ZN(n678) );
  XOR2_X1 U739 ( .A(KEYINPUT117), .B(n678), .Z(n690) );
  NOR2_X1 U740 ( .A1(n510), .A2(n679), .ZN(n681) );
  NOR2_X1 U741 ( .A1(n681), .A2(n680), .ZN(n685) );
  NOR2_X1 U742 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U743 ( .A1(n685), .A2(n684), .ZN(n688) );
  INV_X1 U744 ( .A(n686), .ZN(n687) );
  NOR2_X1 U745 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U746 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U747 ( .A(n691), .B(KEYINPUT52), .ZN(n692) );
  NOR2_X1 U748 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U749 ( .A1(n694), .A2(G952), .ZN(n697) );
  INV_X1 U750 ( .A(n662), .ZN(n695) );
  NAND2_X1 U751 ( .A1(n695), .A2(n357), .ZN(n696) );
  XNOR2_X1 U752 ( .A(KEYINPUT119), .B(KEYINPUT53), .ZN(n698) );
  XNOR2_X1 U753 ( .A(n699), .B(n698), .ZN(G75) );
  BUF_X1 U754 ( .A(n712), .Z(n739) );
  NAND2_X1 U755 ( .A1(n739), .A2(G217), .ZN(n703) );
  XNOR2_X1 U756 ( .A(n701), .B(KEYINPUT124), .ZN(n702) );
  XNOR2_X1 U757 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X1 U758 ( .A1(n704), .A2(n746), .ZN(G66) );
  NAND2_X1 U759 ( .A1(n712), .A2(G475), .ZN(n708) );
  XOR2_X1 U760 ( .A(KEYINPUT121), .B(KEYINPUT59), .Z(n705) );
  XNOR2_X1 U761 ( .A(n706), .B(n705), .ZN(n707) );
  XNOR2_X1 U762 ( .A(n708), .B(n707), .ZN(n709) );
  NOR2_X2 U763 ( .A1(n709), .A2(n746), .ZN(n711) );
  XNOR2_X1 U764 ( .A(KEYINPUT122), .B(KEYINPUT60), .ZN(n710) );
  XNOR2_X1 U765 ( .A(n711), .B(n710), .ZN(G60) );
  NAND2_X1 U766 ( .A1(n712), .A2(G210), .ZN(n717) );
  XNOR2_X1 U767 ( .A(KEYINPUT84), .B(KEYINPUT54), .ZN(n714) );
  XNOR2_X1 U768 ( .A(n714), .B(KEYINPUT55), .ZN(n715) );
  XNOR2_X1 U769 ( .A(n713), .B(n715), .ZN(n716) );
  XNOR2_X1 U770 ( .A(n717), .B(n716), .ZN(n718) );
  NOR2_X2 U771 ( .A1(n718), .A2(n746), .ZN(n720) );
  XNOR2_X1 U772 ( .A(KEYINPUT88), .B(KEYINPUT56), .ZN(n719) );
  XNOR2_X1 U773 ( .A(n720), .B(n719), .ZN(G51) );
  NOR2_X1 U774 ( .A1(n728), .A2(n724), .ZN(n721) );
  XOR2_X1 U775 ( .A(G104), .B(n721), .Z(G6) );
  XOR2_X1 U776 ( .A(KEYINPUT114), .B(KEYINPUT26), .Z(n723) );
  XNOR2_X1 U777 ( .A(G107), .B(KEYINPUT27), .ZN(n722) );
  XNOR2_X1 U778 ( .A(n723), .B(n722), .ZN(n726) );
  NOR2_X1 U779 ( .A1(n732), .A2(n724), .ZN(n725) );
  XOR2_X1 U780 ( .A(n726), .B(n725), .Z(G9) );
  XNOR2_X1 U781 ( .A(G143), .B(n727), .ZN(G45) );
  NOR2_X1 U782 ( .A1(n728), .A2(n731), .ZN(n730) );
  XNOR2_X1 U783 ( .A(G113), .B(KEYINPUT115), .ZN(n729) );
  XNOR2_X1 U784 ( .A(n730), .B(n729), .ZN(G15) );
  NOR2_X1 U785 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U786 ( .A(G116), .B(n733), .Z(G18) );
  XNOR2_X1 U787 ( .A(n734), .B(G125), .ZN(n735) );
  XNOR2_X1 U788 ( .A(n735), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U789 ( .A(G134), .B(n736), .ZN(G36) );
  XOR2_X1 U790 ( .A(G140), .B(n737), .Z(n738) );
  XNOR2_X1 U791 ( .A(KEYINPUT116), .B(n738), .ZN(G42) );
  NAND2_X1 U792 ( .A1(n739), .A2(G469), .ZN(n744) );
  XOR2_X1 U793 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n740) );
  XNOR2_X1 U794 ( .A(n740), .B(KEYINPUT120), .ZN(n741) );
  XNOR2_X1 U795 ( .A(n742), .B(n741), .ZN(n743) );
  XNOR2_X1 U796 ( .A(n744), .B(n743), .ZN(n745) );
  NOR2_X1 U797 ( .A1(n746), .A2(n745), .ZN(G54) );
  NOR2_X1 U798 ( .A1(n748), .A2(n747), .ZN(n755) );
  NAND2_X1 U799 ( .A1(n657), .A2(n763), .ZN(n749) );
  XOR2_X1 U800 ( .A(KEYINPUT125), .B(n749), .Z(n753) );
  NAND2_X1 U801 ( .A1(G953), .A2(G224), .ZN(n750) );
  XNOR2_X1 U802 ( .A(KEYINPUT61), .B(n750), .ZN(n751) );
  NAND2_X1 U803 ( .A1(n751), .A2(G898), .ZN(n752) );
  NAND2_X1 U804 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U805 ( .A(n755), .B(n754), .ZN(G69) );
  XNOR2_X1 U806 ( .A(n756), .B(n757), .ZN(n760) );
  XOR2_X1 U807 ( .A(G227), .B(n760), .Z(n758) );
  NOR2_X1 U808 ( .A1(n763), .A2(n758), .ZN(n759) );
  NAND2_X1 U809 ( .A1(n759), .A2(G900), .ZN(n766) );
  XNOR2_X1 U810 ( .A(n760), .B(KEYINPUT126), .ZN(n761) );
  XNOR2_X1 U811 ( .A(n762), .B(n761), .ZN(n764) );
  NAND2_X1 U812 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U813 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U814 ( .A(n767), .B(KEYINPUT127), .ZN(G72) );
  XNOR2_X1 U815 ( .A(n768), .B(G119), .ZN(G21) );
  XOR2_X1 U816 ( .A(G131), .B(n769), .Z(G33) );
  XOR2_X1 U817 ( .A(G137), .B(n770), .Z(G39) );
endmodule

