//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 0 0 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n772,
    new_n773, new_n774, new_n775, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981,
    new_n982;
  XOR2_X1   g000(.A(KEYINPUT89), .B(KEYINPUT38), .Z(new_n202));
  XNOR2_X1  g001(.A(G8gat), .B(G36gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  NAND2_X1  g004(.A1(G226gat), .A2(G233gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT75), .ZN(new_n207));
  INV_X1    g006(.A(G169gat), .ZN(new_n208));
  INV_X1    g007(.A(G176gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AND2_X1   g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n210), .B(KEYINPUT67), .C1(new_n211), .C2(KEYINPUT26), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT67), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n212), .B(new_n216), .C1(KEYINPUT26), .C2(new_n210), .ZN(new_n217));
  INV_X1    g016(.A(G183gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT27), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT27), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G183gat), .ZN(new_n221));
  INV_X1    g020(.A(G190gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n219), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  OR2_X1    g022(.A1(new_n223), .A2(KEYINPUT28), .ZN(new_n224));
  AOI22_X1  g023(.A1(new_n223), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n225));
  AND3_X1   g024(.A1(new_n217), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n208), .A2(new_n209), .A3(KEYINPUT23), .ZN(new_n228));
  OAI22_X1  g027(.A1(KEYINPUT64), .A2(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n227), .B(new_n228), .C1(new_n229), .C2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT65), .ZN(new_n233));
  OR2_X1    g032(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n234), .A2(new_n210), .A3(new_n230), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT65), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n235), .A2(new_n236), .A3(new_n227), .A4(new_n228), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT24), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n218), .A2(G190gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n222), .A2(G183gat), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n238), .A2(G183gat), .A3(G190gat), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n233), .A2(new_n237), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT25), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT66), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n248), .B1(new_n241), .B2(new_n243), .ZN(new_n249));
  XNOR2_X1  g048(.A(G183gat), .B(G190gat), .ZN(new_n250));
  OAI211_X1 g049(.A(KEYINPUT66), .B(new_n242), .C1(new_n250), .C2(new_n238), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n232), .A2(new_n246), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n226), .B1(new_n247), .B2(new_n254), .ZN(new_n255));
  OAI211_X1 g054(.A(KEYINPUT77), .B(new_n207), .C1(new_n255), .C2(KEYINPUT29), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n247), .A2(new_n254), .ZN(new_n257));
  INV_X1    g056(.A(new_n226), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n207), .B(KEYINPUT76), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G197gat), .B(G204gat), .ZN(new_n263));
  INV_X1    g062(.A(G211gat), .ZN(new_n264));
  INV_X1    g063(.A(G218gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n263), .B1(KEYINPUT22), .B2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G211gat), .B(G218gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT29), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n245), .A2(new_n246), .B1(new_n252), .B2(new_n253), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n270), .B1(new_n271), .B2(new_n226), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT77), .B1(new_n272), .B2(new_n207), .ZN(new_n273));
  NOR3_X1   g072(.A1(new_n262), .A2(new_n269), .A3(new_n273), .ZN(new_n274));
  XOR2_X1   g073(.A(new_n269), .B(KEYINPUT74), .Z(new_n275));
  OR2_X1    g074(.A1(new_n255), .A2(new_n207), .ZN(new_n276));
  INV_X1    g075(.A(new_n260), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n272), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n275), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT37), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n205), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n272), .A2(new_n207), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT77), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n269), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n285), .A2(new_n286), .A3(new_n261), .A4(new_n256), .ZN(new_n287));
  INV_X1    g086(.A(new_n279), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT37), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n202), .B1(new_n282), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n287), .A2(new_n288), .A3(new_n205), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n285), .A2(new_n261), .A3(new_n256), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  AOI22_X1  g094(.A1(new_n293), .A2(new_n269), .B1(new_n295), .B2(new_n275), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n202), .B1(new_n296), .B2(new_n281), .ZN(new_n297));
  INV_X1    g096(.A(new_n205), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n298), .B1(new_n289), .B2(KEYINPUT37), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n292), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n291), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT70), .ZN(new_n302));
  INV_X1    g101(.A(G120gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G113gat), .ZN(new_n304));
  INV_X1    g103(.A(G113gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G120gat), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT1), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G127gat), .B(G134gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT69), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT69), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n307), .A2(new_n311), .A3(new_n308), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n304), .A2(new_n306), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT1), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n308), .A2(KEYINPUT68), .ZN(new_n317));
  INV_X1    g116(.A(G127gat), .ZN(new_n318));
  OR3_X1    g117(.A1(new_n318), .A2(KEYINPUT68), .A3(G134gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n316), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n302), .B1(new_n313), .B2(new_n320), .ZN(new_n321));
  AND4_X1   g120(.A1(new_n311), .A2(new_n314), .A3(new_n308), .A4(new_n315), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n311), .B1(new_n307), .B2(new_n308), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n302), .B(new_n320), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G148gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT79), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT79), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(G148gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n328), .A2(new_n330), .A3(G141gat), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n327), .A2(G141gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT78), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT78), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n334), .B1(new_n327), .B2(G141gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n331), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(G155gat), .A2(G162gat), .ZN(new_n337));
  INV_X1    g136(.A(G155gat), .ZN(new_n338));
  INV_X1    g137(.A(G162gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n337), .B1(new_n340), .B2(KEYINPUT2), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT2), .ZN(new_n342));
  INV_X1    g141(.A(G141gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n343), .A2(G148gat), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n342), .B1(new_n332), .B2(new_n344), .ZN(new_n345));
  AND2_X1   g144(.A1(new_n340), .A2(new_n337), .ZN(new_n346));
  AOI22_X1  g145(.A1(new_n336), .A2(new_n341), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n326), .A2(KEYINPUT4), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n336), .A2(new_n341), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n345), .A2(new_n346), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT3), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n320), .B1(new_n322), .B2(new_n323), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT3), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n347), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(G225gat), .A2(G233gat), .ZN(new_n357));
  AND2_X1   g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n313), .A2(new_n347), .A3(new_n320), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT4), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n348), .A2(new_n358), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT5), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n353), .A2(new_n351), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n359), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n357), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n363), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n362), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT80), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n326), .A2(new_n369), .A3(new_n360), .A4(new_n347), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n353), .A2(KEYINPUT70), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n371), .A2(new_n360), .A3(new_n347), .A4(new_n324), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(KEYINPUT80), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n359), .A2(KEYINPUT4), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT81), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n359), .A2(KEYINPUT81), .A3(KEYINPUT4), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n370), .A2(new_n373), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT82), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n358), .A2(new_n363), .ZN(new_n380));
  NOR3_X1   g179(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n376), .A2(new_n377), .ZN(new_n382));
  AND2_X1   g181(.A1(new_n372), .A2(KEYINPUT80), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n372), .A2(KEYINPUT80), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n380), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT82), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n368), .B1(new_n381), .B2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G1gat), .B(G29gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n389), .B(KEYINPUT0), .ZN(new_n390));
  XNOR2_X1  g189(.A(G57gat), .B(G85gat), .ZN(new_n391));
  XOR2_X1   g190(.A(new_n390), .B(new_n391), .Z(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n388), .A2(KEYINPUT6), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT83), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n379), .B1(new_n378), .B2(new_n380), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n385), .A2(new_n386), .A3(KEYINPUT82), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n392), .B1(new_n399), .B2(new_n368), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n400), .A2(KEYINPUT83), .A3(KEYINPUT6), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT6), .B1(new_n388), .B2(new_n393), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n397), .A2(new_n398), .B1(new_n362), .B2(new_n367), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n392), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n301), .A2(new_n402), .A3(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT88), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n357), .B1(new_n385), .B2(new_n356), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT39), .B1(new_n365), .B2(new_n366), .ZN(new_n410));
  OR2_X1    g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT87), .B(KEYINPUT39), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n393), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n408), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT40), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n400), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n409), .A2(new_n412), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(new_n392), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n409), .A2(new_n410), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT88), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT40), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n298), .B1(new_n274), .B2(new_n279), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n422), .A2(KEYINPUT30), .A3(new_n292), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT30), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n280), .A2(new_n424), .A3(new_n205), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n423), .A2(KEYINPUT86), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n423), .A2(new_n425), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT86), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n416), .A2(new_n421), .A3(new_n426), .A4(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(G22gat), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n354), .B1(new_n269), .B2(KEYINPUT29), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n351), .ZN(new_n433));
  NAND2_X1  g232(.A1(G228gat), .A2(G233gat), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT29), .B1(new_n347), .B2(new_n354), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n433), .B(new_n435), .C1(new_n275), .C2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n433), .B1(new_n286), .B2(new_n436), .ZN(new_n438));
  XOR2_X1   g237(.A(new_n434), .B(KEYINPUT84), .Z(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n431), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n437), .A2(new_n440), .A3(new_n431), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(KEYINPUT85), .A3(new_n443), .ZN(new_n444));
  XOR2_X1   g243(.A(KEYINPUT31), .B(G50gat), .Z(new_n445));
  XNOR2_X1  g244(.A(G78gat), .B(G106gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  OR2_X1    g247(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT85), .ZN(new_n450));
  INV_X1    g249(.A(new_n443), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n450), .B1(new_n451), .B2(new_n441), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n444), .A2(new_n452), .A3(new_n448), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n407), .A2(new_n430), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT83), .B1(new_n400), .B2(KEYINPUT6), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT6), .ZN(new_n458));
  NOR4_X1   g257(.A1(new_n404), .A2(new_n395), .A3(new_n458), .A4(new_n392), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n406), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(new_n427), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n454), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT71), .B1(new_n321), .B2(new_n325), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT71), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n371), .A2(new_n464), .A3(new_n324), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n463), .A2(new_n259), .A3(new_n465), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n255), .B(KEYINPUT71), .C1(new_n321), .C2(new_n325), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(G227gat), .ZN(new_n469));
  INV_X1    g268(.A(G233gat), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT34), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n471), .B(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(G15gat), .B(G43gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(G71gat), .B(G99gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n474), .B(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n469), .A2(new_n470), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n466), .A2(new_n467), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n476), .B1(new_n478), .B2(KEYINPUT32), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT33), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(KEYINPUT72), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT72), .B1(new_n478), .B2(new_n480), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n479), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n478), .B(KEYINPUT32), .C1(new_n480), .C2(new_n476), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n473), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n473), .B1(new_n485), .B2(new_n484), .ZN(new_n488));
  NOR3_X1   g287(.A1(new_n487), .A2(new_n488), .A3(KEYINPUT36), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n484), .A2(new_n485), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n471), .B(KEYINPUT34), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT73), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT73), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n478), .A2(KEYINPUT32), .ZN(new_n495));
  INV_X1    g294(.A(new_n476), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n483), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n497), .B1(new_n498), .B2(new_n481), .ZN(new_n499));
  INV_X1    g298(.A(new_n485), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n494), .B(new_n491), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n493), .A2(new_n501), .A3(new_n486), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n489), .B1(new_n502), .B2(KEYINPUT36), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n456), .A2(new_n462), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT35), .ZN(new_n505));
  AOI22_X1  g304(.A1(new_n402), .A2(new_n406), .B1(new_n425), .B2(new_n423), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n501), .A2(new_n486), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n494), .B1(new_n490), .B2(new_n491), .ZN(new_n508));
  NOR3_X1   g307(.A1(new_n507), .A2(new_n454), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n505), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT90), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n396), .A2(new_n401), .B1(new_n405), .B2(new_n403), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n423), .A2(KEYINPUT86), .A3(new_n425), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT86), .B1(new_n423), .B2(new_n425), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n511), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n429), .A2(new_n426), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n460), .A2(KEYINPUT90), .A3(new_n517), .ZN(new_n518));
  NOR4_X1   g317(.A1(new_n454), .A2(new_n487), .A3(new_n488), .A4(KEYINPUT35), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n516), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT91), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n510), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n516), .A2(new_n518), .A3(KEYINPUT91), .A4(new_n519), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n504), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(G64gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(G57gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(KEYINPUT97), .B(G57gat), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n526), .B1(new_n527), .B2(new_n525), .ZN(new_n528));
  OR2_X1    g327(.A1(G71gat), .A2(G78gat), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT98), .ZN(new_n530));
  NAND2_X1  g329(.A1(G71gat), .A2(G78gat), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT9), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n529), .A2(new_n531), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT98), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n528), .A2(new_n532), .A3(new_n534), .A4(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G57gat), .B(G64gat), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n531), .B(new_n529), .C1(new_n538), .C2(new_n533), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  XOR2_X1   g340(.A(KEYINPUT99), .B(KEYINPUT21), .Z(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AND2_X1   g342(.A1(G231gat), .A2(G233gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(G127gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(G15gat), .B(G22gat), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT16), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n547), .B1(new_n548), .B2(G1gat), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n549), .B1(G1gat), .B2(new_n547), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(G8gat), .ZN(new_n551));
  INV_X1    g350(.A(G8gat), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n549), .B(new_n552), .C1(G1gat), .C2(new_n547), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n554), .B1(new_n541), .B2(KEYINPUT21), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n546), .B(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(new_n338), .ZN(new_n559));
  XOR2_X1   g358(.A(G183gat), .B(G211gat), .Z(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n557), .B(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT41), .ZN(new_n563));
  INV_X1    g362(.A(G232gat), .ZN(new_n564));
  NOR3_X1   g363(.A1(new_n563), .A2(new_n564), .A3(new_n470), .ZN(new_n565));
  XOR2_X1   g364(.A(G43gat), .B(G50gat), .Z(new_n566));
  INV_X1    g365(.A(KEYINPUT15), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT14), .ZN(new_n570));
  INV_X1    g369(.A(G29gat), .ZN(new_n571));
  INV_X1    g370(.A(G36gat), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n574));
  AOI22_X1  g373(.A1(new_n573), .A2(new_n574), .B1(G29gat), .B2(G36gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n566), .A2(new_n567), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n569), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NOR3_X1   g376(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n574), .B1(new_n578), .B2(KEYINPUT92), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT92), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n573), .A2(new_n580), .ZN(new_n581));
  OAI22_X1  g380(.A1(new_n579), .A2(new_n581), .B1(new_n571), .B2(new_n572), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT93), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n582), .A2(new_n583), .A3(new_n568), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n583), .B1(new_n582), .B2(new_n568), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n577), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(G85gat), .ZN(new_n588));
  INV_X1    g387(.A(G92gat), .ZN(new_n589));
  OAI21_X1  g388(.A(KEYINPUT7), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT7), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n591), .A2(G85gat), .A3(G92gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G99gat), .B(G106gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(G99gat), .A2(G106gat), .ZN(new_n595));
  AOI22_X1  g394(.A1(KEYINPUT8), .A2(new_n595), .B1(new_n588), .B2(new_n589), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n593), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n594), .B1(new_n593), .B2(new_n596), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n565), .B1(new_n587), .B2(new_n600), .ZN(new_n601));
  OAI211_X1 g400(.A(KEYINPUT17), .B(new_n577), .C1(new_n585), .C2(new_n586), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n593), .A2(new_n596), .ZN(new_n603));
  INV_X1    g402(.A(new_n594), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n597), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n586), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(new_n584), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT17), .B1(new_n609), .B2(new_n577), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n601), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G190gat), .B(G218gat), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT101), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(KEYINPUT100), .B(G134gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(G162gat), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n563), .B1(new_n564), .B2(new_n470), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n611), .A2(new_n612), .ZN(new_n620));
  AOI22_X1  g419(.A1(new_n615), .A2(new_n619), .B1(new_n620), .B2(new_n613), .ZN(new_n621));
  AND4_X1   g420(.A1(KEYINPUT101), .A2(new_n613), .A3(new_n620), .A4(new_n619), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n562), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G229gat), .A2(G233gat), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n587), .A2(new_n554), .ZN(new_n627));
  INV_X1    g426(.A(new_n554), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n602), .A2(new_n628), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n626), .B(new_n627), .C1(new_n629), .C2(new_n610), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT94), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT18), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT17), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n587), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n635), .A2(new_n628), .A3(new_n602), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n636), .A2(KEYINPUT94), .A3(new_n626), .A4(new_n627), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n632), .A2(new_n633), .A3(new_n637), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n636), .A2(KEYINPUT18), .A3(new_n626), .A4(new_n627), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n609), .A2(new_n577), .A3(new_n628), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n627), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n626), .B(KEYINPUT13), .Z(new_n642));
  AOI21_X1  g441(.A(KEYINPUT95), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT95), .ZN(new_n644));
  INV_X1    g443(.A(new_n642), .ZN(new_n645));
  AOI211_X1 g444(.A(new_n644), .B(new_n645), .C1(new_n627), .C2(new_n640), .ZN(new_n646));
  OAI211_X1 g445(.A(new_n638), .B(new_n639), .C1(new_n643), .C2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(G113gat), .B(G141gat), .ZN(new_n648));
  INV_X1    g447(.A(G197gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT11), .B(G169gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT12), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n647), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT96), .ZN(new_n656));
  OAI211_X1 g455(.A(new_n639), .B(new_n653), .C1(new_n643), .C2(new_n646), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n656), .B1(new_n658), .B2(new_n638), .ZN(new_n659));
  AND3_X1   g458(.A1(new_n632), .A2(new_n633), .A3(new_n637), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n660), .A2(new_n657), .A3(KEYINPUT96), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n655), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(G230gat), .A2(G233gat), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n597), .A2(KEYINPUT102), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n600), .B1(new_n540), .B2(new_n665), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n606), .A2(new_n539), .A3(new_n537), .A4(new_n664), .ZN(new_n667));
  AOI21_X1  g466(.A(KEYINPUT10), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT10), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n540), .A2(new_n606), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n663), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n663), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n666), .A2(new_n672), .A3(new_n667), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(G120gat), .B(G148gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(G176gat), .B(G204gat), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n675), .B(new_n676), .Z(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n671), .A2(new_n673), .A3(new_n677), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n625), .A2(new_n662), .A3(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n524), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(new_n512), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g485(.A(new_n552), .B1(new_n684), .B2(new_n515), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n520), .A2(new_n521), .ZN(new_n688));
  INV_X1    g487(.A(new_n510), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n688), .A2(new_n523), .A3(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n504), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n683), .ZN(new_n693));
  XOR2_X1   g492(.A(KEYINPUT16), .B(G8gat), .Z(new_n694));
  AND4_X1   g493(.A1(new_n515), .A2(new_n692), .A3(new_n693), .A4(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(KEYINPUT42), .B1(new_n687), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT103), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n684), .A2(new_n515), .A3(new_n694), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT42), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AND3_X1   g499(.A1(new_n696), .A2(new_n697), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n697), .B1(new_n696), .B2(new_n700), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(G1325gat));
  INV_X1    g502(.A(new_n684), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n487), .A2(new_n488), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  OR3_X1    g505(.A1(new_n704), .A2(G15gat), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(G15gat), .B1(new_n704), .B2(new_n503), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(G1326gat));
  NAND2_X1  g508(.A1(new_n684), .A2(new_n454), .ZN(new_n710));
  XNOR2_X1  g509(.A(KEYINPUT43), .B(G22gat), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(G1327gat));
  AOI21_X1  g511(.A(new_n623), .B1(new_n690), .B2(new_n691), .ZN(new_n713));
  INV_X1    g512(.A(new_n562), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n658), .A2(new_n656), .A3(new_n638), .ZN(new_n715));
  OAI21_X1  g514(.A(KEYINPUT96), .B1(new_n660), .B2(new_n657), .ZN(new_n716));
  AOI22_X1  g515(.A1(new_n715), .A2(new_n716), .B1(new_n647), .B2(new_n654), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n714), .A2(new_n717), .A3(new_n681), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n713), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n719), .A2(new_n571), .A3(new_n512), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT45), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n692), .A2(KEYINPUT44), .A3(new_n624), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n723), .B1(new_n524), .B2(new_n623), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n725), .A2(new_n512), .A3(new_n718), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(G29gat), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n721), .A2(new_n727), .ZN(G1328gat));
  NAND3_X1  g527(.A1(new_n719), .A2(new_n572), .A3(new_n515), .ZN(new_n729));
  OR2_X1    g528(.A1(new_n729), .A2(KEYINPUT46), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(KEYINPUT46), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n725), .A2(new_n515), .A3(new_n718), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n730), .B(new_n731), .C1(new_n572), .C2(new_n732), .ZN(G1329gat));
  INV_X1    g532(.A(G43gat), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n503), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n722), .A2(new_n724), .A3(new_n718), .A4(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n713), .A2(new_n705), .A3(new_n718), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n734), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT47), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n736), .A2(new_n738), .A3(KEYINPUT104), .A4(new_n739), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n736), .A2(new_n738), .A3(KEYINPUT104), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n741), .B2(new_n739), .ZN(G1330gat));
  INV_X1    g541(.A(G50gat), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n455), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n722), .A2(new_n724), .A3(new_n718), .A4(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n713), .A2(new_n454), .A3(new_n718), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n743), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g548(.A1(new_n625), .A2(new_n717), .A3(new_n681), .ZN(new_n750));
  XOR2_X1   g549(.A(new_n750), .B(KEYINPUT105), .Z(new_n751));
  NAND2_X1  g550(.A1(new_n692), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n512), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(new_n527), .ZN(G1332gat));
  AOI21_X1  g554(.A(new_n517), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT106), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n759));
  XOR2_X1   g558(.A(new_n758), .B(new_n759), .Z(G1333gat));
  INV_X1    g559(.A(G71gat), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n752), .B2(new_n706), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT107), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n503), .A2(new_n761), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n763), .B1(new_n753), .B2(new_n764), .ZN(new_n765));
  NOR4_X1   g564(.A1(new_n752), .A2(KEYINPUT107), .A3(new_n761), .A4(new_n503), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n762), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(KEYINPUT50), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT50), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n769), .B(new_n762), .C1(new_n765), .C2(new_n766), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n768), .A2(new_n770), .ZN(G1334gat));
  OR3_X1    g570(.A1(new_n752), .A2(KEYINPUT109), .A3(new_n455), .ZN(new_n772));
  OAI21_X1  g571(.A(KEYINPUT109), .B1(new_n752), .B2(new_n455), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(KEYINPUT108), .B(G78gat), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n774), .B(new_n775), .ZN(G1335gat));
  NOR2_X1   g575(.A1(new_n714), .A2(new_n662), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n778), .A2(new_n682), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n725), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(G85gat), .B1(new_n780), .B2(new_n460), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT51), .B1(new_n713), .B2(new_n777), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT51), .ZN(new_n783));
  NOR4_X1   g582(.A1(new_n524), .A2(new_n783), .A3(new_n623), .A4(new_n778), .ZN(new_n784));
  OR2_X1    g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n785), .A2(new_n588), .A3(new_n512), .A4(new_n681), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n781), .A2(new_n786), .ZN(G1336gat));
  NAND4_X1  g586(.A1(new_n722), .A2(new_n724), .A3(new_n515), .A4(new_n779), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(G92gat), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT110), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n517), .A2(G92gat), .A3(new_n682), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n791), .B1(new_n782), .B2(new_n784), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n789), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(KEYINPUT52), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n789), .A2(new_n790), .A3(new_n792), .A4(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(G1337gat));
  OAI21_X1  g596(.A(G99gat), .B1(new_n780), .B2(new_n503), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n706), .A2(G99gat), .A3(new_n682), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n785), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(G1338gat));
  NAND4_X1  g600(.A1(new_n722), .A2(new_n724), .A3(new_n454), .A4(new_n779), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(G106gat), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n455), .A2(G106gat), .A3(new_n682), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n804), .B1(new_n782), .B2(new_n784), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT53), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n803), .A2(new_n808), .A3(new_n805), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n809), .ZN(G1339gat));
  NAND3_X1  g609(.A1(new_n627), .A2(new_n640), .A3(new_n645), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(KEYINPUT113), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n636), .A2(new_n627), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n812), .B1(new_n626), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n652), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n681), .B(new_n815), .C1(new_n659), .C2(new_n661), .ZN(new_n816));
  OR3_X1    g615(.A1(new_n668), .A2(new_n663), .A3(new_n670), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n817), .A2(KEYINPUT54), .A3(new_n671), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n819), .B(new_n663), .C1(new_n668), .C2(new_n670), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n820), .A2(KEYINPUT111), .A3(new_n678), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT111), .B1(new_n820), .B2(new_n678), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n818), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI211_X1 g624(.A(KEYINPUT55), .B(new_n818), .C1(new_n821), .C2(new_n822), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n826), .A2(KEYINPUT112), .A3(new_n680), .ZN(new_n827));
  AOI21_X1  g626(.A(KEYINPUT112), .B1(new_n826), .B2(new_n680), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n825), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n816), .B1(new_n829), .B2(new_n717), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n623), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n829), .A2(new_n623), .ZN(new_n832));
  AOI22_X1  g631(.A1(new_n715), .A2(new_n716), .B1(new_n652), .B2(new_n814), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n714), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  NOR4_X1   g634(.A1(new_n562), .A2(new_n662), .A3(new_n624), .A4(new_n681), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT114), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n836), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT114), .ZN(new_n839));
  AOI22_X1  g638(.A1(new_n830), .A2(new_n623), .B1(new_n832), .B2(new_n833), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n838), .B(new_n839), .C1(new_n840), .C2(new_n714), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n837), .A2(new_n512), .A3(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n705), .A2(new_n455), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n842), .A2(new_n843), .A3(new_n517), .A4(new_n845), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n837), .A2(new_n841), .A3(new_n512), .A4(new_n517), .ZN(new_n847));
  OAI21_X1  g646(.A(KEYINPUT115), .B1(new_n847), .B2(new_n844), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n846), .A2(G113gat), .A3(new_n848), .A4(new_n662), .ZN(new_n849));
  INV_X1    g648(.A(new_n847), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n509), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n305), .B1(new_n851), .B2(new_n717), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n849), .A2(new_n852), .ZN(G1340gat));
  NAND4_X1  g652(.A1(new_n846), .A2(G120gat), .A3(new_n848), .A4(new_n681), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n303), .B1(new_n851), .B2(new_n682), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n854), .A2(new_n855), .ZN(G1341gat));
  AND3_X1   g655(.A1(new_n846), .A2(new_n714), .A3(new_n848), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n714), .A2(new_n318), .ZN(new_n858));
  OAI22_X1  g657(.A1(new_n857), .A2(new_n318), .B1(new_n851), .B2(new_n858), .ZN(G1342gat));
  NAND3_X1  g658(.A1(new_n846), .A2(new_n624), .A3(new_n848), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(G134gat), .ZN(new_n861));
  INV_X1    g660(.A(new_n509), .ZN(new_n862));
  NOR4_X1   g661(.A1(new_n862), .A2(G134gat), .A3(new_n515), .A4(new_n623), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n837), .A2(new_n841), .A3(new_n512), .A4(new_n863), .ZN(new_n864));
  OR3_X1    g663(.A1(new_n864), .A2(KEYINPUT116), .A3(KEYINPUT56), .ZN(new_n865));
  OAI21_X1  g664(.A(KEYINPUT116), .B1(new_n864), .B2(KEYINPUT56), .ZN(new_n866));
  AOI22_X1  g665(.A1(new_n865), .A2(new_n866), .B1(KEYINPUT56), .B2(new_n864), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n861), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(KEYINPUT117), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT117), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n861), .A2(new_n870), .A3(new_n867), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n871), .ZN(G1343gat));
  INV_X1    g671(.A(new_n503), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n873), .A2(new_n455), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n850), .A2(new_n343), .A3(new_n662), .A4(new_n874), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n825), .A2(new_n680), .A3(new_n826), .ZN(new_n876));
  AOI22_X1  g675(.A1(new_n662), .A2(new_n876), .B1(new_n833), .B2(new_n681), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n834), .B1(new_n877), .B2(new_n624), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n836), .B1(new_n878), .B2(new_n562), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n455), .A2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n837), .A2(new_n454), .A3(new_n841), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n883), .B1(new_n884), .B2(new_n880), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n503), .A2(new_n512), .A3(new_n517), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n885), .A2(new_n717), .A3(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n875), .B1(new_n887), .B2(new_n343), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT118), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n889), .B1(new_n887), .B2(new_n343), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n888), .A2(new_n890), .A3(KEYINPUT58), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT58), .ZN(new_n892));
  OAI221_X1 g691(.A(new_n875), .B1(new_n889), .B2(new_n892), .C1(new_n887), .C2(new_n343), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(new_n893), .ZN(G1344gat));
  NOR4_X1   g693(.A1(new_n847), .A2(new_n455), .A3(new_n873), .A4(new_n682), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n328), .B(new_n330), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n885), .A2(new_n886), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n896), .A3(new_n681), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n837), .A2(new_n841), .A3(new_n881), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n880), .B1(new_n879), .B2(new_n455), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n886), .A2(new_n682), .ZN(new_n903));
  OAI211_X1 g702(.A(KEYINPUT59), .B(G148gat), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n897), .A2(new_n899), .A3(new_n904), .ZN(G1345gat));
  NAND2_X1  g704(.A1(new_n714), .A2(G155gat), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT119), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n850), .A2(new_n714), .A3(new_n874), .ZN(new_n908));
  AOI22_X1  g707(.A1(new_n898), .A2(new_n907), .B1(new_n908), .B2(new_n338), .ZN(G1346gat));
  NOR3_X1   g708(.A1(new_n885), .A2(new_n623), .A3(new_n886), .ZN(new_n910));
  INV_X1    g709(.A(new_n842), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n874), .A2(new_n339), .A3(new_n517), .A4(new_n624), .ZN(new_n912));
  OAI22_X1  g711(.A1(new_n910), .A2(new_n339), .B1(new_n911), .B2(new_n912), .ZN(G1347gat));
  NOR2_X1   g712(.A1(new_n512), .A2(new_n517), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n837), .A2(new_n841), .A3(new_n509), .A4(new_n914), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n915), .A2(KEYINPUT120), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(KEYINPUT120), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n916), .A2(new_n662), .A3(new_n917), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n837), .A2(new_n841), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n914), .B(new_n920), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n921), .A2(new_n844), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n919), .A2(KEYINPUT122), .A3(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n922), .A2(new_n841), .A3(new_n837), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT122), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n717), .A2(new_n208), .ZN(new_n928));
  AOI22_X1  g727(.A1(new_n208), .A2(new_n918), .B1(new_n927), .B2(new_n928), .ZN(G1348gat));
  NAND3_X1  g728(.A1(new_n923), .A2(new_n926), .A3(new_n681), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(G176gat), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n916), .A2(new_n209), .A3(new_n681), .A4(new_n917), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(KEYINPUT123), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT123), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n931), .A2(new_n935), .A3(new_n932), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(G1349gat));
  NAND3_X1  g736(.A1(new_n923), .A2(new_n926), .A3(new_n714), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(G183gat), .ZN(new_n939));
  INV_X1    g738(.A(new_n915), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n940), .A2(new_n219), .A3(new_n221), .A4(new_n714), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n942), .A2(KEYINPUT124), .A3(KEYINPUT60), .ZN(new_n943));
  NAND2_X1  g742(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n939), .A2(new_n944), .A3(new_n941), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(new_n945), .ZN(G1350gat));
  NAND4_X1  g745(.A1(new_n916), .A2(new_n222), .A3(new_n624), .A4(new_n917), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n923), .A2(new_n926), .A3(new_n624), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT61), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n948), .A2(new_n949), .A3(G190gat), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n949), .B1(new_n948), .B2(G190gat), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n947), .B1(new_n950), .B2(new_n951), .ZN(G1351gat));
  AND2_X1   g751(.A1(new_n919), .A2(new_n914), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(new_n874), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(G197gat), .B1(new_n955), .B2(new_n662), .ZN(new_n956));
  OR2_X1    g755(.A1(new_n921), .A2(new_n873), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n957), .B1(new_n900), .B2(new_n901), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n717), .A2(new_n649), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(G1352gat));
  INV_X1    g759(.A(G204gat), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n681), .A2(new_n961), .ZN(new_n962));
  XOR2_X1   g761(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n963));
  INV_X1    g762(.A(new_n963), .ZN(new_n964));
  OR3_X1    g763(.A1(new_n954), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n954), .B2(new_n962), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n958), .A2(new_n681), .ZN(new_n967));
  OAI211_X1 g766(.A(new_n965), .B(new_n966), .C1(new_n961), .C2(new_n967), .ZN(G1353gat));
  NAND3_X1  g767(.A1(new_n955), .A2(new_n264), .A3(new_n714), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT126), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n958), .A2(new_n970), .A3(new_n714), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n971), .A2(G211gat), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n970), .B1(new_n958), .B2(new_n714), .ZN(new_n973));
  INV_X1    g772(.A(new_n973), .ZN(new_n974));
  AOI21_X1  g773(.A(KEYINPUT63), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n971), .A2(G211gat), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT63), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n976), .A2(new_n977), .A3(new_n973), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n969), .B1(new_n975), .B2(new_n978), .ZN(G1354gat));
  AOI21_X1  g778(.A(G218gat), .B1(new_n955), .B2(new_n624), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n624), .A2(G218gat), .ZN(new_n981));
  XNOR2_X1  g780(.A(new_n981), .B(KEYINPUT127), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n980), .B1(new_n958), .B2(new_n982), .ZN(G1355gat));
endmodule


