//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 0 1 0 1 0 0 0 1 1 0 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 1 1 0 1 0 0 0 0 0 0 0 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1263, new_n1264, new_n1265, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n206), .A2(new_n207), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(KEYINPUT65), .B(G77), .ZN(new_n220));
  AND2_X1   g0020(.A1(new_n220), .A2(G244), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G50), .A2(G226), .ZN(new_n225));
  NAND4_X1  g0025(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n211), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n214), .B(new_n219), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G226), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  XNOR2_X1  g0038(.A(G68), .B(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT66), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G50), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G58), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  AND2_X1   g0047(.A1(new_n247), .A2(new_n216), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n208), .A2(G20), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT8), .B(G58), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n217), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  AOI22_X1  g0054(.A1(new_n251), .A2(new_n253), .B1(G150), .B2(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n248), .B1(new_n249), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G13), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(G1), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G20), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n247), .A2(new_n216), .ZN(new_n261));
  INV_X1    g0061(.A(G1), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n261), .B1(new_n262), .B2(G20), .ZN(new_n263));
  MUX2_X1   g0063(.A(new_n260), .B(new_n263), .S(G50), .Z(new_n264));
  NOR2_X1   g0064(.A1(new_n256), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT9), .ZN(new_n266));
  XNOR2_X1  g0066(.A(new_n265), .B(new_n266), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT3), .B(G33), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(G223), .A3(G1698), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT3), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n220), .ZN(new_n275));
  INV_X1    g0075(.A(G1698), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n268), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G222), .ZN(new_n278));
  OAI211_X1 g0078(.A(new_n269), .B(new_n275), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n262), .B1(G41), .B2(G45), .ZN(new_n282));
  INV_X1    g0082(.A(G274), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G41), .ZN(new_n285));
  OAI211_X1 g0085(.A(G1), .B(G13), .C1(new_n270), .C2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n282), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n284), .B1(new_n288), .B2(G226), .ZN(new_n289));
  AOI21_X1  g0089(.A(KEYINPUT67), .B1(new_n281), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n281), .A2(KEYINPUT67), .A3(new_n289), .ZN(new_n292));
  AOI21_X1  g0092(.A(G190), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n292), .ZN(new_n294));
  NOR3_X1   g0094(.A1(new_n294), .A2(G200), .A3(new_n290), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n267), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT69), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT10), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n297), .A2(KEYINPUT10), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n296), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G190), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n301), .B1(new_n294), .B2(new_n290), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n291), .A2(new_n292), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n302), .B1(new_n303), .B2(G200), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n304), .A2(new_n297), .A3(KEYINPUT10), .A4(new_n267), .ZN(new_n305));
  INV_X1    g0105(.A(new_n265), .ZN(new_n306));
  INV_X1    g0106(.A(G169), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G179), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n309), .B1(new_n291), .B2(new_n292), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n306), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n300), .A2(new_n305), .A3(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n258), .A2(G20), .A3(new_n203), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n313), .B(KEYINPUT12), .ZN(new_n314));
  INV_X1    g0114(.A(new_n263), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n314), .B1(new_n203), .B2(new_n315), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n254), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n317));
  INV_X1    g0117(.A(G77), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n317), .B1(new_n318), .B2(new_n252), .ZN(new_n319));
  AND3_X1   g0119(.A1(new_n319), .A2(KEYINPUT11), .A3(new_n261), .ZN(new_n320));
  AOI21_X1  g0120(.A(KEYINPUT11), .B1(new_n319), .B2(new_n261), .ZN(new_n321));
  NOR3_X1   g0121(.A1(new_n316), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n271), .A2(new_n273), .A3(G226), .A4(new_n276), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n271), .A2(new_n273), .A3(G232), .A4(G1698), .ZN(new_n325));
  NAND2_X1  g0125(.A1(G33), .A2(G97), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT70), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT70), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n324), .A2(new_n325), .A3(new_n329), .A4(new_n326), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n328), .A2(new_n330), .A3(new_n280), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n284), .B1(new_n288), .B2(G238), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT13), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT13), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n331), .A2(new_n335), .A3(new_n332), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n334), .A2(G179), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n307), .B1(new_n334), .B2(new_n336), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT14), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n336), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n335), .B1(new_n331), .B2(new_n332), .ZN(new_n342));
  OAI21_X1  g0142(.A(G169), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n343), .A2(KEYINPUT14), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n323), .B1(new_n340), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G200), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(new_n341), .B2(new_n342), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n334), .A2(new_n301), .A3(new_n336), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n323), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n345), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(G58), .A2(G68), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n204), .A2(new_n205), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(G20), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n254), .A2(G159), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT71), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT71), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n354), .A2(new_n358), .A3(new_n355), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT7), .ZN(new_n360));
  NOR3_X1   g0160(.A1(new_n268), .A2(new_n360), .A3(G20), .ZN(new_n361));
  AOI21_X1  g0161(.A(KEYINPUT7), .B1(new_n274), .B2(new_n217), .ZN(new_n362));
  OAI21_X1  g0162(.A(G68), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n357), .A2(KEYINPUT16), .A3(new_n359), .A4(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT16), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT73), .B1(new_n270), .B2(KEYINPUT3), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT72), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n272), .B2(G33), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT73), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n369), .A2(new_n272), .A3(G33), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n270), .A2(KEYINPUT72), .A3(KEYINPUT3), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n366), .A2(new_n368), .A3(new_n370), .A4(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n360), .A2(G20), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n360), .B1(new_n268), .B2(G20), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n203), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n365), .B1(new_n376), .B2(new_n356), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n364), .A2(new_n377), .A3(new_n261), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n259), .A2(new_n250), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(new_n263), .B2(new_n250), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n271), .A2(new_n273), .A3(G223), .A4(new_n276), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n271), .A2(new_n273), .A3(G226), .A4(G1698), .ZN(new_n383));
  INV_X1    g0183(.A(G87), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n382), .B(new_n383), .C1(new_n270), .C2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n280), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n284), .B1(new_n288), .B2(G232), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n386), .A2(new_n387), .A3(new_n309), .ZN(new_n388));
  INV_X1    g0188(.A(new_n284), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n287), .B2(new_n233), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(new_n280), .B2(new_n385), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n388), .B1(new_n391), .B2(G169), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n381), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT18), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT18), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n381), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n386), .A2(new_n387), .A3(new_n301), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n398), .B1(new_n391), .B2(G200), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n378), .A2(new_n380), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT17), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n378), .A2(KEYINPUT17), .A3(new_n380), .A4(new_n399), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n395), .A2(new_n397), .A3(new_n402), .A4(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(G244), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n389), .B1(new_n287), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n268), .A2(G238), .A3(G1698), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n274), .A2(G107), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n407), .B(new_n408), .C1(new_n277), .C2(new_n233), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n406), .B1(new_n409), .B2(new_n280), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT68), .B1(new_n410), .B2(new_n346), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(G190), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n251), .A2(new_n254), .B1(new_n220), .B2(G20), .ZN(new_n414));
  XNOR2_X1  g0214(.A(KEYINPUT15), .B(G87), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n253), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n248), .B1(new_n414), .B2(new_n417), .ZN(new_n418));
  OAI22_X1  g0218(.A1(new_n315), .A2(new_n318), .B1(new_n220), .B2(new_n259), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT68), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n413), .B(new_n420), .C1(new_n421), .C2(new_n412), .ZN(new_n422));
  OR2_X1    g0222(.A1(new_n418), .A2(new_n419), .ZN(new_n423));
  AND2_X1   g0223(.A1(new_n410), .A2(G179), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n410), .A2(new_n307), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  NOR4_X1   g0227(.A1(new_n312), .A2(new_n351), .A3(new_n404), .A4(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  OR2_X1    g0229(.A1(KEYINPUT5), .A2(G41), .ZN(new_n430));
  NAND2_X1  g0230(.A1(KEYINPUT5), .A2(G41), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(G45), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n433), .A2(G1), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n435), .A2(G270), .A3(new_n286), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT74), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n262), .A2(G45), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n438), .B1(new_n430), .B2(new_n431), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n437), .B1(new_n439), .B2(G274), .ZN(new_n440));
  NOR2_X1   g0240(.A1(KEYINPUT5), .A2(G41), .ZN(new_n441));
  AND2_X1   g0241(.A1(KEYINPUT5), .A2(G41), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n434), .B(G274), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(KEYINPUT74), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n436), .B1(new_n440), .B2(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n272), .A2(G33), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n270), .A2(KEYINPUT3), .ZN(new_n447));
  NOR2_X1   g0247(.A1(KEYINPUT77), .A2(G303), .ZN(new_n448));
  AND2_X1   g0248(.A1(KEYINPUT77), .A2(G303), .ZN(new_n449));
  OAI22_X1  g0249(.A1(new_n446), .A2(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT78), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n271), .A2(new_n273), .A3(G264), .A4(G1698), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n271), .A2(new_n273), .A3(G257), .A4(new_n276), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n450), .A2(new_n451), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n454), .A2(new_n280), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n450), .A2(new_n452), .A3(new_n453), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT78), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n445), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT20), .ZN(new_n459));
  INV_X1    g0259(.A(G116), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n217), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G283), .ZN(new_n462));
  INV_X1    g0262(.A(G97), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n462), .B1(new_n463), .B2(G33), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n461), .B1(new_n464), .B2(new_n217), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n459), .B1(new_n465), .B2(new_n248), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n270), .A2(G97), .ZN(new_n467));
  AOI21_X1  g0267(.A(G20), .B1(new_n467), .B2(new_n462), .ZN(new_n468));
  OAI211_X1 g0268(.A(KEYINPUT20), .B(new_n261), .C1(new_n468), .C2(new_n461), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n262), .A2(G33), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n248), .A2(new_n259), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G116), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n259), .A2(new_n460), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n458), .A2(G179), .A3(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT79), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n432), .A2(new_n437), .A3(G274), .A4(new_n434), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n443), .A2(KEYINPUT74), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n280), .B1(new_n434), .B2(new_n432), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n479), .A2(new_n480), .B1(new_n481), .B2(G270), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n456), .A2(KEYINPUT78), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n454), .A2(new_n280), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n307), .B1(new_n470), .B2(new_n475), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n478), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT21), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n477), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AOI211_X1 g0289(.A(new_n478), .B(KEYINPUT21), .C1(new_n485), .C2(new_n486), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n485), .A2(new_n346), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n457), .A2(new_n280), .A3(new_n454), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n492), .A2(new_n301), .A3(new_n482), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n476), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NOR3_X1   g0294(.A1(new_n489), .A2(new_n490), .A3(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n271), .A2(new_n273), .A3(G250), .A4(new_n276), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n271), .A2(new_n273), .A3(G257), .A4(G1698), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G294), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n280), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n480), .A2(new_n479), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n435), .A2(G264), .A3(new_n286), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n504), .A2(new_n309), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n280), .A2(new_n500), .B1(new_n481), .B2(G264), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n307), .B1(new_n506), .B2(new_n502), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n271), .A2(new_n273), .A3(new_n217), .A4(G87), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT22), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT22), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n268), .A2(new_n511), .A3(new_n217), .A4(G87), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT24), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G33), .A2(G116), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n515), .A2(G20), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT23), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(new_n217), .B2(G107), .ZN(new_n518));
  INV_X1    g0318(.A(G107), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n519), .A2(KEYINPUT23), .A3(G20), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n516), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n513), .A2(new_n514), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT80), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT80), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n513), .A2(new_n524), .A3(new_n514), .A4(new_n521), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n513), .A2(new_n521), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(KEYINPUT24), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n523), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n261), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n258), .A2(G20), .A3(new_n519), .ZN(new_n530));
  OR2_X1    g0330(.A1(new_n530), .A2(KEYINPUT25), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(KEYINPUT25), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n531), .B(new_n532), .C1(new_n519), .C2(new_n472), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n508), .B1(new_n529), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n533), .B1(new_n528), .B2(new_n261), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n501), .A2(new_n502), .A3(new_n301), .A4(new_n503), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT81), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n504), .A2(new_n346), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n504), .A2(KEYINPUT81), .A3(new_n346), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n536), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n519), .B1(new_n374), .B2(new_n375), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT6), .ZN(new_n545));
  AND2_X1   g0345(.A1(G97), .A2(G107), .ZN(new_n546));
  NOR2_X1   g0346(.A1(G97), .A2(G107), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n519), .A2(KEYINPUT6), .A3(G97), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(G20), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n254), .A2(G77), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n261), .B1(new_n544), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n260), .A2(G97), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n555), .B1(new_n472), .B2(G97), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n271), .A2(new_n273), .A3(G244), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT4), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n560), .A2(G1698), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n562), .A2(new_n271), .A3(new_n273), .A4(G244), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n561), .A2(new_n462), .A3(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n271), .A2(new_n273), .A3(G250), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n276), .B1(new_n565), .B2(KEYINPUT4), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n280), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n479), .A2(new_n480), .B1(new_n481), .B2(G257), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n567), .A2(G179), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n307), .B1(new_n567), .B2(new_n568), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n558), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT19), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n217), .B1(new_n326), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(G87), .A2(G97), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n519), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n217), .A2(G33), .A3(G97), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n573), .A2(new_n575), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n268), .A2(new_n217), .A3(G68), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n248), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n416), .A2(new_n259), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g0381(.A(new_n415), .B(KEYINPUT76), .ZN(new_n582));
  INV_X1    g0382(.A(new_n472), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n271), .A2(new_n273), .A3(G238), .A4(new_n276), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n271), .A2(new_n273), .A3(G244), .A4(G1698), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n586), .A2(new_n587), .A3(new_n515), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n280), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT75), .ZN(new_n590));
  INV_X1    g0390(.A(G250), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n283), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n434), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n438), .A2(new_n590), .A3(G250), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n286), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n589), .A2(G179), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n280), .B1(new_n593), .B2(new_n594), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n598), .B1(new_n280), .B2(new_n588), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n597), .B1(new_n599), .B2(new_n307), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n589), .A2(new_n301), .A3(new_n596), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n599), .B2(G200), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n472), .A2(new_n384), .ZN(new_n603));
  NOR3_X1   g0403(.A1(new_n579), .A2(new_n603), .A3(new_n580), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n585), .A2(new_n600), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n550), .A2(G20), .B1(G77), .B2(new_n254), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n274), .A2(new_n217), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n372), .A2(new_n373), .B1(new_n607), .B2(new_n360), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n606), .B1(new_n608), .B2(new_n519), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n556), .B1(new_n609), .B2(new_n261), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n567), .A2(new_n301), .A3(new_n568), .ZN(new_n611));
  AOI21_X1  g0411(.A(G200), .B1(new_n567), .B2(new_n568), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n543), .A2(new_n571), .A3(new_n605), .A4(new_n613), .ZN(new_n614));
  NOR4_X1   g0414(.A1(new_n429), .A2(new_n496), .A3(new_n535), .A4(new_n614), .ZN(G372));
  NOR3_X1   g0415(.A1(new_n535), .A2(new_n489), .A3(new_n490), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n616), .A2(new_n614), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n600), .A2(new_n585), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n602), .A2(new_n604), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(KEYINPUT26), .B1(new_n620), .B2(new_n571), .ZN(new_n621));
  INV_X1    g0421(.A(new_n570), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n567), .A2(G179), .A3(new_n568), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n610), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT26), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n624), .A2(new_n605), .A3(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n621), .A2(new_n626), .A3(new_n618), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n428), .B1(new_n617), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n311), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n345), .A2(new_n426), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n402), .A2(new_n403), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(new_n350), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n396), .B1(new_n381), .B2(new_n393), .ZN(new_n633));
  AOI211_X1 g0433(.A(KEYINPUT18), .B(new_n392), .C1(new_n378), .C2(new_n380), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n300), .A2(new_n305), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n629), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n628), .A2(new_n638), .ZN(G369));
  INV_X1    g0439(.A(new_n476), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n262), .A2(G13), .ZN(new_n641));
  OR3_X1    g0441(.A1(new_n641), .A2(KEYINPUT27), .A3(G20), .ZN(new_n642));
  OAI21_X1  g0442(.A(KEYINPUT27), .B1(new_n641), .B2(G20), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(G213), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT82), .ZN(new_n645));
  XNOR2_X1  g0445(.A(new_n644), .B(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(G343), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n496), .B1(new_n640), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n489), .A2(new_n490), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n651), .A2(new_n476), .A3(new_n648), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n650), .A2(G330), .A3(new_n652), .ZN(new_n653));
  NOR3_X1   g0453(.A1(new_n536), .A2(new_n508), .A3(new_n648), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n543), .B1(new_n536), .B2(new_n649), .ZN(new_n655));
  INV_X1    g0455(.A(new_n535), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n653), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT83), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(new_n651), .B2(new_n648), .ZN(new_n662));
  OAI211_X1 g0462(.A(KEYINPUT83), .B(new_n649), .C1(new_n489), .C2(new_n490), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n654), .B1(new_n664), .B2(new_n657), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n660), .A2(new_n665), .ZN(G399));
  NAND3_X1  g0466(.A1(new_n574), .A2(new_n519), .A3(new_n460), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n212), .A2(new_n285), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(new_n669), .A3(G1), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT84), .ZN(new_n671));
  INV_X1    g0471(.A(new_n669), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n215), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n670), .A2(KEYINPUT84), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n671), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT28), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n536), .A2(new_n542), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n605), .A2(new_n571), .A3(new_n613), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n679), .A2(new_n495), .A3(new_n656), .A4(new_n649), .ZN(new_n680));
  XNOR2_X1  g0480(.A(KEYINPUT86), .B(KEYINPUT30), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n492), .A2(KEYINPUT85), .A3(G179), .A4(new_n482), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n567), .A2(new_n568), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n599), .A2(new_n506), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n683), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  OAI211_X1 g0487(.A(G179), .B(new_n482), .C1(new_n483), .C2(new_n484), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT85), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n682), .B1(new_n687), .B2(new_n690), .ZN(new_n691));
  AND4_X1   g0491(.A1(new_n506), .A2(new_n567), .A3(new_n568), .A4(new_n599), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n690), .A2(new_n692), .A3(KEYINPUT30), .A4(new_n683), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n599), .A2(G179), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n485), .A2(new_n694), .A3(new_n684), .A4(new_n504), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n648), .B1(new_n691), .B2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT31), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n683), .A2(new_n685), .A3(new_n686), .ZN(new_n700));
  AOI21_X1  g0500(.A(KEYINPUT85), .B1(new_n458), .B2(G179), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n681), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n702), .A2(new_n693), .A3(new_n695), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n703), .A2(KEYINPUT31), .A3(new_n648), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n680), .A2(new_n699), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G330), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT29), .ZN(new_n707));
  AND3_X1   g0507(.A1(new_n605), .A2(new_n571), .A3(new_n613), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n476), .A2(G169), .ZN(new_n709));
  OAI21_X1  g0509(.A(KEYINPUT79), .B1(new_n709), .B2(new_n458), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(KEYINPUT21), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n487), .A2(new_n488), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(new_n712), .A3(new_n477), .ZN(new_n713));
  OAI211_X1 g0513(.A(new_n543), .B(new_n708), .C1(new_n713), .C2(new_n535), .ZN(new_n714));
  AND3_X1   g0514(.A1(new_n621), .A2(new_n626), .A3(new_n618), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n648), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT87), .ZN(new_n717));
  OAI211_X1 g0517(.A(KEYINPUT88), .B(new_n707), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT88), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n649), .B1(new_n617), .B2(new_n627), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n719), .B1(new_n720), .B2(KEYINPUT87), .ZN(new_n721));
  OAI21_X1  g0521(.A(KEYINPUT29), .B1(new_n716), .B2(KEYINPUT88), .ZN(new_n722));
  OAI211_X1 g0522(.A(new_n706), .B(new_n718), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n676), .B1(new_n724), .B2(G1), .ZN(G364));
  NOR2_X1   g0525(.A1(new_n257), .A2(G20), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n262), .B1(new_n726), .B2(G45), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(new_n672), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n653), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n650), .A2(new_n652), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n731), .B1(G330), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(G13), .A2(G33), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G20), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n733), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n217), .A2(G190), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(new_n309), .A3(G200), .ZN(new_n741));
  OR2_X1    g0541(.A1(new_n741), .A2(KEYINPUT90), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(KEYINPUT90), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n309), .A2(new_n346), .ZN(new_n746));
  NAND2_X1  g0546(.A1(G20), .A2(G190), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT92), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI22_X1  g0551(.A1(G283), .A2(new_n745), .B1(new_n751), .B2(G326), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT91), .ZN(new_n753));
  AND3_X1   g0553(.A1(new_n746), .A2(new_n753), .A3(new_n740), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n753), .B1(new_n746), .B2(new_n740), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XOR2_X1   g0556(.A(KEYINPUT33), .B(G317), .Z(new_n757));
  OAI21_X1  g0557(.A(new_n752), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n309), .A2(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n740), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n747), .A2(new_n346), .A3(G179), .ZN(new_n762));
  AOI22_X1  g0562(.A1(new_n761), .A2(G311), .B1(new_n762), .B2(G303), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n759), .A2(new_n748), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n268), .B1(new_n765), .B2(G322), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G179), .A2(G200), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n740), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G329), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n217), .B1(new_n767), .B2(G190), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G294), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n763), .A2(new_n766), .A3(new_n770), .A4(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n749), .ZN(new_n775));
  AOI22_X1  g0575(.A1(G50), .A2(new_n775), .B1(new_n765), .B2(G58), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n762), .A2(G87), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n771), .A2(new_n463), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n274), .B1(new_n761), .B2(new_n220), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n776), .A2(new_n777), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G159), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n768), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT32), .ZN(new_n784));
  OAI221_X1 g0584(.A(new_n784), .B1(new_n203), .B2(new_n756), .C1(new_n519), .C2(new_n744), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n758), .A2(new_n774), .B1(new_n781), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n216), .B1(G20), .B2(new_n307), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n730), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n268), .A2(new_n212), .ZN(new_n789));
  INV_X1    g0589(.A(G355), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n789), .A2(new_n790), .B1(G116), .B2(new_n212), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n242), .A2(G45), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n274), .A2(new_n212), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n793), .B1(new_n215), .B2(new_n433), .ZN(new_n794));
  XOR2_X1   g0594(.A(new_n794), .B(KEYINPUT89), .Z(new_n795));
  AOI21_X1  g0595(.A(new_n791), .B1(new_n792), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n737), .A2(new_n787), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n788), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n734), .B1(new_n739), .B2(new_n799), .ZN(G396));
  NAND2_X1  g0600(.A1(new_n648), .A2(new_n423), .ZN(new_n801));
  AND2_X1   g0601(.A1(new_n411), .A2(new_n412), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n420), .B1(new_n412), .B2(new_n421), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n426), .B(new_n801), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(KEYINPUT93), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT93), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n422), .A2(new_n807), .A3(new_n426), .A4(new_n801), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n716), .A2(new_n810), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n426), .A2(new_n649), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(new_n805), .B2(new_n808), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT94), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n814), .B(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n811), .B1(new_n816), .B2(new_n716), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n706), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n729), .B1(new_n818), .B2(new_n819), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n814), .A2(new_n735), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n744), .A2(new_n203), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n274), .B1(new_n769), .B2(G132), .ZN(new_n825));
  INV_X1    g0625(.A(new_n762), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n825), .B1(new_n207), .B2(new_n826), .C1(new_n202), .C2(new_n771), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n775), .A2(G137), .B1(new_n761), .B2(G159), .ZN(new_n828));
  INV_X1    g0628(.A(G143), .ZN(new_n829));
  INV_X1    g0629(.A(G150), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n828), .B1(new_n829), .B2(new_n764), .C1(new_n830), .C2(new_n756), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT34), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n824), .B(new_n827), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n832), .B2(new_n831), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n760), .A2(new_n460), .ZN(new_n835));
  INV_X1    g0635(.A(G294), .ZN(new_n836));
  INV_X1    g0636(.A(G311), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n764), .A2(new_n836), .B1(new_n768), .B2(new_n837), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n835), .B(new_n838), .C1(G303), .C2(new_n775), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n745), .A2(G87), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n268), .B(new_n778), .C1(G107), .C2(new_n762), .ZN(new_n841));
  INV_X1    g0641(.A(new_n756), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(G283), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n839), .A2(new_n840), .A3(new_n841), .A4(new_n843), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n834), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n787), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n787), .A2(new_n735), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n730), .B(new_n847), .C1(new_n318), .C2(new_n848), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n821), .A2(new_n822), .B1(new_n823), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(G384));
  OAI211_X1 g0651(.A(G116), .B(new_n218), .C1(new_n550), .C2(KEYINPUT35), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(KEYINPUT35), .B2(new_n550), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n853), .B(KEYINPUT36), .ZN(new_n854));
  INV_X1    g0654(.A(new_n353), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n855), .A2(G50), .A3(new_n220), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n207), .A2(G68), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n262), .B(G13), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n699), .A2(KEYINPUT97), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT31), .B1(new_n703), .B2(new_n648), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT97), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n860), .A2(new_n863), .A3(new_n680), .A4(new_n704), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n649), .A2(new_n322), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n345), .A2(new_n350), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n343), .A2(KEYINPUT14), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n338), .A2(new_n339), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n868), .A2(new_n869), .A3(new_n337), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n323), .B(new_n648), .C1(new_n870), .C2(new_n349), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n814), .B1(new_n867), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n864), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n357), .A2(new_n359), .A3(new_n363), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n365), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n875), .A2(new_n261), .A3(new_n364), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n646), .B1(new_n876), .B2(new_n380), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n878), .B1(new_n631), .B2(new_n635), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n644), .B(KEYINPUT82), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n381), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT37), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n394), .A2(new_n881), .A3(new_n882), .A4(new_n400), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n386), .A2(new_n387), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n307), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n880), .B1(new_n885), .B2(new_n388), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n886), .B1(new_n876), .B2(new_n380), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n378), .A2(new_n380), .A3(new_n399), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT37), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n883), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT38), .ZN(new_n891));
  NOR3_X1   g0691(.A1(new_n879), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n404), .A2(new_n877), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n883), .A2(new_n889), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT38), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT95), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n891), .B1(new_n879), .B2(new_n890), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n893), .A2(KEYINPUT38), .A3(new_n894), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT95), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n873), .B1(new_n896), .B2(new_n900), .ZN(new_n901));
  OR2_X1    g0701(.A1(new_n901), .A2(KEYINPUT40), .ZN(new_n902));
  INV_X1    g0702(.A(new_n873), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n394), .A2(new_n881), .A3(new_n400), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT37), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n905), .A2(KEYINPUT96), .A3(new_n883), .ZN(new_n906));
  INV_X1    g0706(.A(new_n881), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n404), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT96), .B1(new_n905), .B2(new_n883), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n891), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n898), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n903), .A2(KEYINPUT40), .A3(new_n912), .ZN(new_n913));
  AND2_X1   g0713(.A1(new_n902), .A2(new_n913), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n428), .A2(new_n864), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n913), .B(G330), .C1(new_n901), .C2(KEYINPUT40), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n428), .A2(new_n864), .A3(G330), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n914), .A2(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OR2_X1    g0718(.A1(new_n426), .A2(new_n648), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n920), .B1(new_n716), .B2(new_n810), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n867), .A2(new_n871), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n897), .A2(new_n899), .A3(new_n898), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n899), .B1(new_n897), .B2(new_n898), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n635), .A2(new_n880), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n870), .A2(new_n323), .A3(new_n649), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT39), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n911), .A2(new_n932), .A3(new_n898), .ZN(new_n933));
  OAI21_X1  g0733(.A(KEYINPUT39), .B1(new_n892), .B2(new_n895), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n930), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n718), .B1(new_n721), .B2(new_n722), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n428), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n638), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n936), .B(new_n939), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n918), .A2(new_n940), .B1(new_n262), .B2(new_n726), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n918), .A2(new_n940), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n859), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n943), .B(KEYINPUT98), .Z(G367));
  OAI211_X1 g0744(.A(new_n571), .B(new_n613), .C1(new_n610), .C2(new_n649), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n624), .A2(new_n648), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(KEYINPUT83), .B1(new_n713), .B2(new_n649), .ZN(new_n948));
  INV_X1    g0748(.A(new_n663), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n657), .B(new_n947), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(KEYINPUT100), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT100), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n664), .A2(new_n952), .A3(new_n657), .A4(new_n947), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(KEYINPUT42), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT42), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n951), .A2(new_n956), .A3(new_n953), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n571), .B1(new_n656), .B2(new_n945), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n649), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n649), .A2(new_n604), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n960), .A2(new_n605), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(new_n618), .B2(new_n960), .ZN(new_n962));
  XOR2_X1   g0762(.A(KEYINPUT99), .B(KEYINPUT43), .Z(new_n963));
  NOR2_X1   g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n955), .A2(new_n957), .A3(new_n959), .A4(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(KEYINPUT101), .ZN(new_n966));
  AND2_X1   g0766(.A1(new_n957), .A2(new_n959), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT101), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n967), .A2(new_n968), .A3(new_n955), .A4(new_n964), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n964), .B1(KEYINPUT43), .B2(new_n962), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n957), .A2(new_n959), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n956), .B1(new_n951), .B2(new_n953), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n966), .A2(new_n969), .A3(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n947), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n660), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n966), .A2(new_n969), .A3(new_n976), .A4(new_n973), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n669), .B(KEYINPUT41), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n657), .B1(new_n948), .B2(new_n949), .ZN(new_n981));
  INV_X1    g0781(.A(new_n654), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n981), .A2(new_n982), .A3(new_n947), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT45), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(KEYINPUT45), .B1(new_n665), .B2(new_n947), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(KEYINPUT44), .B1(new_n665), .B2(new_n947), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n981), .A2(new_n982), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT44), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n989), .A2(new_n990), .A3(new_n975), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n988), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n659), .B1(new_n987), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n658), .A2(new_n662), .A3(new_n663), .ZN(new_n994));
  AND3_X1   g0794(.A1(new_n994), .A2(new_n653), .A3(new_n981), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n653), .B1(new_n994), .B2(new_n981), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n997), .A2(new_n723), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n983), .A2(new_n984), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n665), .A2(KEYINPUT45), .A3(new_n947), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n1001), .A2(new_n660), .A3(new_n988), .A4(new_n991), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n993), .A2(new_n998), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n980), .B1(new_n1003), .B2(new_n724), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n978), .B(new_n979), .C1(new_n1004), .C2(new_n728), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n237), .A2(new_n793), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n797), .B1(new_n212), .B2(new_n415), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n729), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n826), .A2(new_n202), .B1(new_n760), .B2(new_n207), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n772), .A2(G68), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1010), .B(new_n268), .C1(new_n830), .C2(new_n764), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n1009), .B(new_n1011), .C1(G137), .C2(new_n769), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n745), .A2(new_n220), .B1(G159), .B2(new_n842), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1012), .B(new_n1013), .C1(new_n829), .C2(new_n750), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n449), .A2(new_n448), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n750), .A2(new_n837), .B1(new_n1015), .B2(new_n764), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT102), .Z(new_n1017));
  NOR2_X1   g0817(.A1(new_n826), .A2(new_n460), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n1018), .A2(KEYINPUT46), .B1(new_n519), .B2(new_n771), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(KEYINPUT46), .B2(new_n1018), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n842), .A2(G294), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n745), .A2(G97), .ZN(new_n1022));
  INV_X1    g0822(.A(G317), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n274), .B1(new_n768), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(G283), .B2(new_n761), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .A4(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1014), .B1(new_n1017), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT47), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  AND2_X1   g0829(.A1(new_n1029), .A2(new_n787), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1008), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n738), .B2(new_n962), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1005), .A2(new_n1033), .ZN(G387));
  INV_X1    g0834(.A(new_n998), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n997), .A2(new_n723), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1035), .A2(new_n672), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n997), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n789), .A2(new_n668), .B1(G107), .B2(new_n212), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n234), .A2(G45), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n250), .A2(G50), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT50), .ZN(new_n1042));
  AOI211_X1 g0842(.A(G45), .B(new_n667), .C1(G68), .C2(G77), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n793), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1039), .B1(new_n1040), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n729), .B1(new_n1045), .B2(new_n798), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT103), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n268), .B1(new_n760), .B2(new_n203), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n764), .A2(new_n207), .B1(new_n768), .B2(new_n830), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n1048), .B(new_n1049), .C1(new_n220), .C2(new_n762), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n842), .A2(new_n251), .B1(new_n582), .B2(new_n772), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n749), .A2(new_n782), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT104), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1050), .A2(new_n1022), .A3(new_n1051), .A4(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n268), .B1(new_n769), .B2(G326), .ZN(new_n1055));
  INV_X1    g0855(.A(G283), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n826), .A2(new_n836), .B1(new_n771), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1015), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n761), .A2(new_n1058), .B1(new_n765), .B2(G317), .ZN(new_n1059));
  INV_X1    g0859(.A(G322), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1059), .B1(new_n756), .B2(new_n837), .C1(new_n750), .C2(new_n1060), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT105), .Z(new_n1062));
  AOI21_X1  g0862(.A(new_n1057), .B1(new_n1062), .B2(KEYINPUT48), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(KEYINPUT48), .B2(new_n1062), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT49), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1055), .B1(new_n460), .B2(new_n744), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1054), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1047), .B1(new_n1068), .B2(new_n787), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n658), .A2(new_n737), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n1038), .A2(new_n728), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1037), .A2(new_n1071), .ZN(G393));
  NAND2_X1  g0872(.A1(new_n1003), .A2(new_n672), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n998), .B1(new_n993), .B2(new_n1002), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n993), .A2(new_n728), .A3(new_n1002), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n245), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n797), .B1(new_n463), .B2(new_n212), .C1(new_n1077), .C2(new_n793), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n729), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G294), .A2(new_n761), .B1(new_n772), .B2(G116), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n756), .B2(new_n1015), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT106), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n744), .A2(new_n519), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n749), .A2(new_n1023), .B1(new_n764), .B2(new_n837), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT52), .Z(new_n1085));
  OAI221_X1 g0885(.A(new_n274), .B1(new_n768), .B2(new_n1060), .C1(new_n826), .C2(new_n1056), .ZN(new_n1086));
  NOR4_X1   g0886(.A1(new_n1082), .A2(new_n1083), .A3(new_n1085), .A4(new_n1086), .ZN(new_n1087));
  OR2_X1    g0887(.A1(new_n1087), .A2(KEYINPUT107), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(KEYINPUT107), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n749), .A2(new_n830), .B1(new_n764), .B2(new_n782), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT51), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n826), .A2(new_n203), .B1(new_n760), .B2(new_n250), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n771), .A2(new_n318), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n268), .B1(new_n768), .B2(new_n829), .ZN(new_n1094));
  NOR3_X1   g0894(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n842), .A2(G50), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n840), .A2(new_n1091), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1088), .A2(new_n1089), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1079), .B1(new_n1098), .B2(new_n787), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n738), .B2(new_n947), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1076), .A2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(KEYINPUT108), .B1(new_n1075), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1101), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT108), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1103), .B(new_n1104), .C1(new_n1074), .C2(new_n1073), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1102), .A2(new_n1105), .ZN(G390));
  OAI211_X1 g0906(.A(new_n912), .B(new_n931), .C1(new_n923), .C2(new_n921), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n931), .B1(new_n921), .B2(new_n923), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n933), .A2(new_n1108), .A3(new_n934), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n819), .A2(new_n872), .ZN(new_n1110));
  AND3_X1   g0910(.A1(new_n1107), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n680), .B(new_n704), .C1(new_n862), .C2(new_n861), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n863), .ZN(new_n1113));
  OAI211_X1 g0913(.A(G330), .B(new_n872), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1111), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n728), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n730), .B1(new_n250), .B2(new_n848), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n268), .B(new_n1093), .C1(G87), .C2(new_n762), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n775), .A2(G283), .B1(new_n761), .B2(G97), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(G116), .A2(new_n765), .B1(new_n769), .B2(G294), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n824), .B(new_n1122), .C1(G107), .C2(new_n842), .ZN(new_n1123));
  INV_X1    g0923(.A(G125), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n268), .B1(new_n1124), .B2(new_n768), .C1(new_n744), .C2(new_n207), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT113), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1128));
  NOR3_X1   g0928(.A1(new_n826), .A2(KEYINPUT53), .A3(new_n830), .ZN(new_n1129));
  OAI21_X1  g0929(.A(KEYINPUT53), .B1(new_n826), .B2(new_n830), .ZN(new_n1130));
  INV_X1    g0930(.A(G128), .ZN(new_n1131));
  INV_X1    g0931(.A(G132), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n1130), .B1(new_n1131), .B2(new_n749), .C1(new_n1132), .C2(new_n764), .ZN(new_n1133));
  NOR4_X1   g0933(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .A4(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(KEYINPUT54), .B(G143), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n760), .A2(new_n1135), .B1(new_n771), .B2(new_n782), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(new_n842), .B2(G137), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT112), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1123), .B1(new_n1134), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n933), .A2(new_n934), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n1118), .B1(new_n846), .B2(new_n1139), .C1(new_n1140), .C2(new_n736), .ZN(new_n1141));
  AND2_X1   g0941(.A1(new_n1117), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT109), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n917), .A2(new_n1143), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n428), .A2(new_n864), .A3(KEYINPUT109), .A4(G330), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n938), .A2(new_n638), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n864), .A2(new_n816), .A3(G330), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n921), .B(new_n1110), .C1(new_n1148), .C2(new_n922), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT110), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n814), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n705), .A2(G330), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n923), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n1114), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n811), .A2(new_n919), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1150), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  AOI211_X1 g0956(.A(KEYINPUT110), .B(new_n921), .C1(new_n1153), .C2(new_n1114), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1149), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1116), .A2(new_n1147), .A3(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1159), .A2(KEYINPUT111), .A3(new_n672), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1158), .A2(new_n1147), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1107), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1162), .B1(new_n1163), .B2(new_n1114), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1161), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1160), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(KEYINPUT111), .B1(new_n1159), .B2(new_n672), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1142), .B1(new_n1166), .B2(new_n1167), .ZN(G378));
  INV_X1    g0968(.A(KEYINPUT115), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT57), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n265), .A2(new_n646), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n312), .B(new_n1171), .ZN(new_n1172));
  XOR2_X1   g0972(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1173));
  XNOR2_X1  g0973(.A(new_n1172), .B(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n930), .B2(new_n935), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n931), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1140), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n896), .A2(new_n900), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n928), .B1(new_n1178), .B2(new_n924), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1174), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1177), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  AND3_X1   g0981(.A1(new_n1175), .A2(new_n1181), .A3(new_n916), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n916), .B1(new_n1175), .B2(new_n1181), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1146), .B1(new_n1116), .B2(new_n1158), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1169), .B(new_n1170), .C1(new_n1184), .C2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1147), .B1(new_n1161), .B2(new_n1164), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1187), .B(KEYINPUT57), .C1(new_n1183), .C2(new_n1182), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1186), .A2(new_n672), .A3(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1187), .B1(new_n1183), .B2(new_n1182), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1169), .B1(new_n1190), .B2(new_n1170), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n582), .A2(new_n761), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1193), .B1(new_n463), .B2(new_n756), .C1(new_n202), .C2(new_n744), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(G107), .A2(new_n765), .B1(new_n769), .B2(G283), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n775), .A2(G116), .B1(new_n220), .B2(new_n762), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n268), .A2(G41), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1195), .A2(new_n1196), .A3(new_n1010), .A4(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1194), .A2(new_n1198), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT114), .Z(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(KEYINPUT58), .ZN(new_n1201));
  AOI211_X1 g1001(.A(G50), .B(new_n1197), .C1(new_n270), .C2(new_n285), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n826), .A2(new_n1135), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n749), .A2(new_n1124), .B1(new_n764), .B2(new_n1131), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1203), .B(new_n1204), .C1(G137), .C2(new_n761), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1205), .B1(new_n1132), .B2(new_n756), .C1(new_n830), .C2(new_n771), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1207));
  AOI211_X1 g1007(.A(G33), .B(G41), .C1(new_n769), .C2(G124), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n744), .B2(new_n782), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n1206), .B2(KEYINPUT59), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1202), .B1(new_n1207), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1201), .A2(new_n1211), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1200), .A2(KEYINPUT58), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n787), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n848), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1214), .B(new_n729), .C1(G50), .C2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n1180), .B2(new_n735), .ZN(new_n1217));
  OR2_X1    g1017(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1217), .B1(new_n1218), .B2(new_n728), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1192), .A2(new_n1219), .ZN(G375));
  NAND2_X1  g1020(.A1(new_n923), .A2(new_n735), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n729), .B1(new_n1215), .B2(G68), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n274), .B1(new_n744), .B2(new_n318), .ZN(new_n1223));
  XOR2_X1   g1023(.A(new_n1223), .B(KEYINPUT117), .Z(new_n1224));
  NAND2_X1  g1024(.A1(new_n842), .A2(G116), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n749), .A2(new_n836), .B1(new_n760), .B2(new_n519), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(G303), .B2(new_n769), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n582), .A2(new_n772), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n765), .A2(G283), .B1(G97), .B2(new_n762), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1225), .A2(new_n1227), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  OR3_X1    g1030(.A1(new_n1224), .A2(KEYINPUT118), .A3(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(KEYINPUT118), .B1(new_n1224), .B2(new_n1230), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n274), .B1(new_n745), .B2(G58), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1233), .A2(KEYINPUT119), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(KEYINPUT119), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(G132), .A2(new_n775), .B1(new_n765), .B2(G137), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n782), .B2(new_n826), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(G150), .A2(new_n761), .B1(new_n769), .B2(G128), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n207), .B2(new_n771), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1235), .B(new_n1240), .C1(new_n756), .C2(new_n1135), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1231), .B(new_n1232), .C1(new_n1234), .C2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1222), .B1(new_n1242), .B2(new_n787), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n1158), .A2(new_n728), .B1(new_n1221), .B2(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(KEYINPUT116), .B1(new_n1158), .B2(new_n1147), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n921), .B1(new_n1153), .B2(new_n1114), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1246), .B(new_n1150), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT116), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1247), .A2(new_n1248), .A3(new_n1146), .A4(new_n1149), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1245), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n980), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1161), .A2(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1244), .B1(new_n1250), .B2(new_n1252), .ZN(G381));
  INV_X1    g1053(.A(new_n1167), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1254), .A2(new_n1160), .A3(new_n1165), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1192), .A2(new_n1255), .A3(new_n1142), .A4(new_n1219), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(G393), .A2(G396), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1257), .A2(new_n850), .A3(new_n1258), .ZN(new_n1259));
  OR3_X1    g1059(.A1(new_n1259), .A2(G387), .A3(G381), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1256), .A2(new_n1260), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(new_n1261), .B(KEYINPUT120), .ZN(G407));
  NAND2_X1  g1062(.A1(new_n647), .A2(G213), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1256), .A2(new_n1263), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(new_n1264), .B(KEYINPUT121), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(G407), .A2(new_n1265), .A3(G213), .ZN(G409));
  INV_X1    g1066(.A(KEYINPUT63), .ZN(new_n1267));
  OAI211_X1 g1067(.A(G378), .B(new_n1219), .C1(new_n1189), .C2(new_n1191), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1219), .B1(new_n980), .B2(new_n1190), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1269), .A2(new_n1255), .A3(new_n1142), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1268), .A2(new_n1270), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1158), .A2(new_n1147), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n669), .B1(new_n1272), .B2(KEYINPUT60), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT60), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1274), .B1(new_n1158), .B2(new_n1147), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1273), .B1(new_n1250), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1244), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n850), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1276), .A2(G384), .A3(new_n1244), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1271), .A2(new_n1263), .A3(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1267), .B1(new_n1282), .B2(KEYINPUT122), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT124), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT123), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(G387), .A2(new_n1285), .A3(new_n1105), .A4(new_n1102), .ZN(new_n1286));
  AND2_X1   g1086(.A1(G393), .A2(G396), .ZN(new_n1287));
  OR2_X1    g1087(.A1(new_n1287), .A2(new_n1258), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT123), .B1(new_n1005), .B2(new_n1033), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1257), .A2(new_n1290), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1284), .B1(new_n1289), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1290), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(G390), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1294), .A2(KEYINPUT124), .A3(new_n1286), .A4(new_n1288), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1288), .B1(G390), .B2(G387), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1296), .B1(G387), .B2(G390), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1292), .A2(new_n1295), .A3(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT61), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1263), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1300), .B1(new_n1268), .B2(new_n1270), .ZN(new_n1301));
  AND3_X1   g1101(.A1(new_n1276), .A2(G384), .A3(new_n1244), .ZN(new_n1302));
  AOI21_X1  g1102(.A(G384), .B1(new_n1276), .B2(new_n1244), .ZN(new_n1303));
  OAI211_X1 g1103(.A(G2897), .B(new_n1300), .C1(new_n1302), .C2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1300), .A2(G2897), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1278), .A2(new_n1279), .A3(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1304), .A2(new_n1306), .ZN(new_n1307));
  OAI211_X1 g1107(.A(new_n1298), .B(new_n1299), .C1(new_n1301), .C2(new_n1307), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1283), .A2(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1282), .A2(KEYINPUT122), .A3(new_n1267), .ZN(new_n1310));
  AOI21_X1  g1110(.A(KEYINPUT125), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1308), .ZN(new_n1312));
  AOI211_X1 g1112(.A(new_n1300), .B(new_n1280), .C1(new_n1268), .C2(new_n1270), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT122), .ZN(new_n1314));
  OAI21_X1  g1114(.A(KEYINPUT63), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  AND4_X1   g1115(.A1(KEYINPUT125), .A2(new_n1312), .A3(new_n1315), .A4(new_n1310), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT126), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1299), .B1(new_n1301), .B2(new_n1307), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT62), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1319), .B1(new_n1301), .B2(new_n1281), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1318), .A2(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1301), .A2(new_n1319), .A3(new_n1281), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1317), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1271), .A2(new_n1263), .ZN(new_n1324));
  AND2_X1   g1124(.A1(new_n1304), .A2(new_n1306), .ZN(new_n1325));
  AOI21_X1  g1125(.A(KEYINPUT61), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1282), .A2(KEYINPUT62), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1326), .A2(new_n1327), .A3(new_n1317), .A4(new_n1322), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1298), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  OAI22_X1  g1130(.A1(new_n1311), .A2(new_n1316), .B1(new_n1323), .B2(new_n1330), .ZN(G405));
  NAND2_X1  g1131(.A1(G375), .A2(G378), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(new_n1256), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1333), .A2(new_n1281), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1332), .A2(new_n1256), .A3(new_n1280), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1334), .A2(new_n1298), .A3(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT127), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1334), .A2(KEYINPUT127), .A3(new_n1298), .A4(new_n1335), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1340), .A2(new_n1329), .ZN(new_n1341));
  AND3_X1   g1141(.A1(new_n1338), .A2(new_n1339), .A3(new_n1341), .ZN(G402));
endmodule


