//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 0 1 0 1 0 0 1 0 0 1 1 0 1 0 1 0 0 1 0 1 1 0 0 0 0 0 0 1 1 1 1 0 0 1 0 1 1 0 0 0 0 0 0 1 0 1 0 1 0 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1250, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  OAI21_X1  g0011(.A(G50), .B1(G58), .B2(G68), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G68), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n208), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n211), .B(new_n217), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT64), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  INV_X1    g0046(.A(G1698), .ZN(new_n247));
  OR2_X1    g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  AOI21_X1  g0049(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  AND2_X1   g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  NOR2_X1   g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI22_X1  g0053(.A1(new_n250), .A2(G223), .B1(new_n253), .B2(G77), .ZN(new_n254));
  AOI21_X1  g0054(.A(G1698), .B1(new_n248), .B2(new_n249), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G222), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G274), .ZN(new_n260));
  AND2_X1   g0060(.A1(G1), .A2(G13), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G33), .A2(G41), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G41), .ZN(new_n264));
  INV_X1    g0064(.A(G45), .ZN(new_n265));
  AOI21_X1  g0065(.A(G1), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n264), .A2(new_n265), .ZN(new_n268));
  INV_X1    g0068(.A(G1), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT66), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT66), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G1), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n268), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n261), .A2(new_n262), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  XOR2_X1   g0076(.A(KEYINPUT65), .B(G226), .Z(new_n277));
  AOI21_X1  g0077(.A(new_n267), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n259), .A2(G190), .A3(new_n278), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n259), .A2(new_n278), .ZN(new_n280));
  INV_X1    g0080(.A(G200), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G20), .A2(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G150), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT8), .B(G58), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n215), .A2(G33), .ZN(new_n286));
  OAI221_X1 g0086(.A(new_n284), .B1(new_n201), .B2(new_n215), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(KEYINPUT67), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT67), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n290), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n289), .A2(new_n214), .A3(new_n291), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n270), .A2(new_n272), .A3(G13), .A4(G20), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G50), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n287), .A2(new_n292), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT70), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n270), .A2(new_n272), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n292), .B1(G20), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G50), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n296), .A2(new_n297), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n297), .B1(new_n296), .B2(new_n300), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT9), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n296), .A2(new_n300), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT70), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT9), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n306), .A2(new_n307), .A3(new_n301), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n282), .B1(new_n304), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT10), .ZN(new_n310));
  OAI21_X1  g0110(.A(KEYINPUT72), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n281), .B1(new_n259), .B2(new_n278), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n312), .B1(G190), .B2(new_n280), .ZN(new_n313));
  NOR3_X1   g0113(.A1(new_n302), .A2(KEYINPUT9), .A3(new_n303), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n307), .B1(new_n306), .B2(new_n301), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT72), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT10), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n311), .A2(new_n318), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n310), .B(new_n313), .C1(new_n314), .C2(new_n315), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT71), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n309), .A2(KEYINPUT71), .A3(new_n310), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G179), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n280), .A2(new_n326), .ZN(new_n327));
  XOR2_X1   g0127(.A(new_n327), .B(KEYINPUT68), .Z(new_n328));
  OAI211_X1 g0128(.A(new_n328), .B(new_n305), .C1(G169), .C2(new_n280), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n293), .A2(new_n285), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n330), .B1(new_n299), .B2(new_n285), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  AND3_X1   g0132(.A1(new_n289), .A2(new_n214), .A3(new_n291), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n248), .A2(KEYINPUT7), .A3(new_n215), .A4(new_n249), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT77), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n253), .A2(KEYINPUT77), .A3(KEYINPUT7), .A4(new_n215), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT7), .ZN(new_n338));
  XNOR2_X1  g0138(.A(KEYINPUT3), .B(G33), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n338), .B1(new_n339), .B2(G20), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n336), .A2(new_n337), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(G68), .ZN(new_n342));
  INV_X1    g0142(.A(G58), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n343), .A2(new_n219), .ZN(new_n344));
  NOR2_X1   g0144(.A1(G58), .A2(G68), .ZN(new_n345));
  OAI21_X1  g0145(.A(G20), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G159), .ZN(new_n347));
  INV_X1    g0147(.A(new_n283), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT16), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n333), .B1(new_n342), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n219), .B1(new_n340), .B2(new_n334), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n350), .B1(new_n353), .B2(new_n349), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n332), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT78), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(new_n275), .B2(new_n231), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n273), .A2(KEYINPUT78), .A3(G232), .A4(new_n274), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI211_X1 g0159(.A(G223), .B(new_n247), .C1(new_n251), .C2(new_n252), .ZN(new_n360));
  OAI211_X1 g0160(.A(G226), .B(G1698), .C1(new_n251), .C2(new_n252), .ZN(new_n361));
  INV_X1    g0161(.A(G33), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n360), .B(new_n361), .C1(new_n362), .C2(new_n221), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n267), .B1(new_n363), .B2(new_n258), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n359), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n281), .ZN(new_n366));
  INV_X1    g0166(.A(G190), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n359), .A2(new_n364), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n355), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT17), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n359), .A2(new_n364), .A3(G179), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(G169), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n375), .B1(new_n359), .B2(new_n364), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT18), .B1(new_n377), .B2(new_n355), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n365), .A2(G169), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n373), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT18), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n342), .A2(new_n351), .ZN(new_n382));
  AND3_X1   g0182(.A1(new_n382), .A2(new_n292), .A3(new_n354), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n380), .B(new_n381), .C1(new_n383), .C2(new_n332), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n355), .A2(new_n369), .A3(KEYINPUT17), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n372), .A2(new_n378), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n299), .A2(G77), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n294), .A2(new_n202), .ZN(new_n388));
  NAND2_X1  g0188(.A1(G20), .A2(G77), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n285), .B2(new_n348), .ZN(new_n390));
  INV_X1    g0190(.A(new_n286), .ZN(new_n391));
  XNOR2_X1  g0191(.A(KEYINPUT15), .B(G87), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n390), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n387), .B(new_n388), .C1(new_n333), .C2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT69), .ZN(new_n396));
  OR2_X1    g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n395), .A2(new_n396), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n250), .A2(G238), .B1(new_n253), .B2(G107), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n255), .A2(G232), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n258), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n267), .B1(new_n276), .B2(G244), .ZN(new_n404));
  AOI21_X1  g0204(.A(G169), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AND2_X1   g0205(.A1(new_n403), .A2(new_n404), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n405), .B1(new_n326), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n399), .A2(new_n407), .ZN(new_n408));
  OR2_X1    g0208(.A1(new_n406), .A2(new_n281), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n406), .A2(G190), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n408), .B1(new_n411), .B2(new_n399), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n386), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n325), .A2(new_n329), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n299), .A2(G68), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT11), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n348), .A2(new_n295), .ZN(new_n417));
  OAI22_X1  g0217(.A1(new_n286), .A2(new_n202), .B1(new_n215), .B2(G68), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n292), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n415), .B1(new_n416), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n416), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n294), .A2(KEYINPUT12), .A3(new_n219), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT12), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(new_n293), .B2(G68), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n421), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n420), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n263), .A2(new_n266), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n428), .B1(new_n275), .B2(new_n220), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT13), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n231), .A2(G1698), .ZN(new_n432));
  OAI221_X1 g0232(.A(new_n432), .B1(G226), .B2(G1698), .C1(new_n251), .C2(new_n252), .ZN(new_n433));
  NAND2_X1  g0233(.A1(G33), .A2(G97), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n274), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n430), .A2(new_n431), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT73), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT13), .B1(new_n429), .B2(new_n435), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  OAI211_X1 g0240(.A(KEYINPUT73), .B(KEYINPUT13), .C1(new_n429), .C2(new_n435), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n440), .A2(G169), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT14), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(KEYINPUT75), .ZN(new_n444));
  AND2_X1   g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n444), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n440), .A2(G169), .A3(new_n441), .A4(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n437), .A2(G179), .A3(new_n439), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n427), .B1(new_n445), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n440), .A2(G200), .A3(new_n441), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT74), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT74), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n440), .A2(new_n453), .A3(G200), .A4(new_n441), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n437), .A2(G190), .A3(new_n439), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n426), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n450), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT76), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n450), .A2(new_n459), .A3(KEYINPUT76), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n414), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  OAI211_X1 g0266(.A(G244), .B(new_n247), .C1(new_n251), .C2(new_n252), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT81), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n339), .A2(KEYINPUT81), .A3(G244), .A4(new_n247), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT4), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AND2_X1   g0272(.A1(KEYINPUT4), .A2(G244), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n247), .B(new_n473), .C1(new_n251), .C2(new_n252), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT82), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n339), .A2(KEYINPUT82), .A3(new_n247), .A4(new_n473), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(G250), .B(G1698), .C1(new_n251), .C2(new_n252), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G283), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n472), .A2(new_n478), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n258), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n264), .A2(KEYINPUT83), .A3(KEYINPUT5), .ZN(new_n485));
  AOI21_X1  g0285(.A(KEYINPUT83), .B1(new_n264), .B2(KEYINPUT5), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n270), .A2(new_n272), .A3(G45), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT5), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G41), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n487), .A2(new_n488), .A3(new_n263), .A4(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n270), .A2(new_n272), .A3(new_n490), .A4(G45), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n489), .A2(G41), .ZN(new_n493));
  OAI211_X1 g0293(.A(G257), .B(new_n274), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n484), .A2(KEYINPUT85), .A3(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT85), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n481), .B1(new_n476), .B2(new_n477), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n274), .B1(new_n499), .B2(new_n472), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n498), .B1(new_n500), .B2(new_n495), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n497), .A2(new_n501), .A3(new_n375), .ZN(new_n502));
  AOI21_X1  g0302(.A(KEYINPUT7), .B1(new_n253), .B2(new_n215), .ZN(new_n503));
  INV_X1    g0303(.A(new_n334), .ZN(new_n504));
  OAI211_X1 g0304(.A(KEYINPUT80), .B(G107), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  XNOR2_X1  g0305(.A(KEYINPUT79), .B(KEYINPUT6), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n204), .A2(G107), .ZN(new_n507));
  OR2_X1    g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(G97), .A2(G107), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n506), .A2(new_n206), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(G20), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n283), .A2(G77), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n505), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n340), .A2(new_n334), .ZN(new_n514));
  AOI21_X1  g0314(.A(KEYINPUT80), .B1(new_n514), .B2(G107), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n292), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n293), .A2(G97), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n270), .A2(new_n272), .A3(G33), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n333), .A2(new_n293), .A3(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n517), .B1(new_n520), .B2(G97), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n495), .A2(KEYINPUT84), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT84), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n491), .A2(new_n494), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n526), .A2(new_n326), .A3(new_n484), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n367), .B1(new_n497), .B2(new_n501), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n523), .A2(new_n525), .B1(new_n483), .B2(new_n258), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n516), .B(new_n521), .C1(new_n530), .C2(new_n281), .ZN(new_n531));
  OAI22_X1  g0331(.A1(new_n502), .A2(new_n528), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT86), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n531), .ZN(new_n535));
  AOI21_X1  g0335(.A(KEYINPUT85), .B1(new_n484), .B2(new_n496), .ZN(new_n536));
  NOR3_X1   g0336(.A1(new_n500), .A2(new_n498), .A3(new_n495), .ZN(new_n537));
  OAI21_X1  g0337(.A(G190), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n326), .A2(new_n530), .B1(new_n516), .B2(new_n521), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n497), .A2(new_n501), .A3(new_n375), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n539), .A2(KEYINPUT86), .A3(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT87), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n339), .A2(G244), .A3(G1698), .ZN(new_n545));
  OAI211_X1 g0345(.A(G238), .B(new_n247), .C1(new_n251), .C2(new_n252), .ZN(new_n546));
  NAND2_X1  g0346(.A1(G33), .A2(G116), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n258), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n488), .A2(new_n260), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n270), .A2(new_n272), .A3(G45), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n258), .B1(new_n551), .B2(new_n222), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n544), .B1(new_n554), .B2(new_n367), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n548), .A2(new_n258), .B1(new_n550), .B2(new_n552), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n556), .A2(KEYINPUT87), .A3(G190), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n556), .A2(new_n281), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n339), .A2(new_n215), .A3(G68), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT19), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n215), .B1(new_n434), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(G87), .B2(new_n206), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n561), .B1(new_n286), .B2(new_n204), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n560), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n292), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n294), .A2(new_n392), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n566), .B(new_n567), .C1(new_n221), .C2(new_n519), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n559), .A2(new_n568), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n549), .A2(new_n326), .A3(new_n553), .ZN(new_n570));
  AOI21_X1  g0370(.A(G169), .B1(new_n549), .B2(new_n553), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n566), .B(new_n567), .C1(new_n392), .C2(new_n519), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n558), .A2(new_n569), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n534), .A2(new_n543), .A3(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(G257), .B(G1698), .C1(new_n251), .C2(new_n252), .ZN(new_n576));
  NAND2_X1  g0376(.A1(G33), .A2(G294), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT90), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n580), .B1(new_n255), .B2(G250), .ZN(new_n581));
  OAI211_X1 g0381(.A(G250), .B(new_n247), .C1(new_n251), .C2(new_n252), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n582), .A2(KEYINPUT90), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n579), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n258), .ZN(new_n585));
  OAI211_X1 g0385(.A(G264), .B(new_n274), .C1(new_n492), .C2(new_n493), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n585), .A2(new_n326), .A3(new_n491), .A4(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n255), .A2(new_n580), .A3(G250), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n582), .A2(KEYINPUT90), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n578), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n491), .B(new_n586), .C1(new_n590), .C2(new_n274), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n375), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n215), .B(G87), .C1(new_n251), .C2(new_n252), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(KEYINPUT22), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT22), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n339), .A2(new_n595), .A3(new_n215), .A4(G87), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT23), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(new_n215), .B2(G107), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n205), .A2(KEYINPUT23), .A3(G20), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n391), .A2(G116), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT24), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT24), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n597), .A2(new_n604), .A3(new_n601), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n333), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  XNOR2_X1  g0406(.A(KEYINPUT89), .B(KEYINPUT25), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n294), .A2(new_n205), .A3(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT89), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n609), .B(KEYINPUT25), .C1(new_n293), .C2(G107), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n608), .B(new_n610), .C1(new_n519), .C2(new_n205), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n587), .B(new_n592), .C1(new_n606), .C2(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n333), .A2(G116), .A3(new_n293), .A4(new_n518), .ZN(new_n613));
  INV_X1    g0413(.A(G116), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n294), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(G20), .B1(G33), .B2(G283), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n362), .A2(G97), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n616), .A2(new_n617), .B1(G20), .B2(new_n614), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n292), .A2(KEYINPUT20), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(KEYINPUT20), .B1(new_n292), .B2(new_n618), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n613), .B(new_n615), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  OAI211_X1 g0421(.A(G264), .B(G1698), .C1(new_n251), .C2(new_n252), .ZN(new_n622));
  OAI211_X1 g0422(.A(G257), .B(new_n247), .C1(new_n251), .C2(new_n252), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n248), .A2(G303), .A3(new_n249), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n258), .ZN(new_n626));
  OAI211_X1 g0426(.A(G270), .B(new_n274), .C1(new_n492), .C2(new_n493), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(new_n491), .A3(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n621), .A2(KEYINPUT21), .A3(new_n628), .A4(G169), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n626), .A2(new_n491), .A3(new_n627), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n630), .A2(G179), .A3(new_n621), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n621), .A2(G169), .A3(new_n628), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT21), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n612), .A2(new_n632), .A3(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n605), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n604), .B1(new_n597), .B2(new_n601), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n292), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n585), .A2(G190), .A3(new_n491), .A4(new_n586), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n591), .A2(G200), .ZN(new_n641));
  INV_X1    g0441(.A(new_n611), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n639), .A2(new_n640), .A3(new_n641), .A4(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT88), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n621), .B1(new_n630), .B2(G190), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n628), .A2(G200), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n621), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n626), .A2(G190), .A3(new_n491), .A4(new_n627), .ZN(new_n649));
  AND4_X1   g0449(.A1(new_n644), .A2(new_n648), .A3(new_n646), .A4(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n643), .B1(new_n647), .B2(new_n650), .ZN(new_n651));
  NOR4_X1   g0451(.A1(new_n466), .A2(new_n575), .A3(new_n636), .A4(new_n651), .ZN(G372));
  AND2_X1   g0452(.A1(new_n378), .A2(new_n384), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT92), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n408), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n399), .A2(KEYINPUT92), .A3(new_n407), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n459), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(new_n450), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n355), .A2(new_n369), .A3(KEYINPUT17), .ZN(new_n661));
  AOI21_X1  g0461(.A(KEYINPUT17), .B1(new_n355), .B2(new_n369), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n654), .B1(new_n660), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n325), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n329), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n558), .A2(new_n569), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n572), .A2(new_n573), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n668), .A2(new_n643), .A3(new_n669), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n670), .A2(new_n539), .A3(new_n542), .A4(new_n636), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n669), .ZN(new_n672));
  AND4_X1   g0472(.A1(KEYINPUT26), .A2(new_n574), .A3(new_n541), .A4(new_n540), .ZN(new_n673));
  OAI21_X1  g0473(.A(KEYINPUT91), .B1(new_n502), .B2(new_n528), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT91), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n540), .A2(new_n675), .A3(new_n541), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n674), .A2(new_n574), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT26), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n673), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n465), .B1(new_n672), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n667), .A2(new_n680), .ZN(G369));
  AND2_X1   g0481(.A1(new_n632), .A2(new_n635), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n215), .A2(G13), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n298), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT27), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n298), .A2(new_n686), .A3(new_n683), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n685), .A2(G213), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(G343), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(KEYINPUT93), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT93), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n688), .A2(new_n691), .A3(G343), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n621), .ZN(new_n694));
  OAI211_X1 g0494(.A(new_n682), .B(new_n694), .C1(new_n647), .C2(new_n650), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n682), .B2(new_n694), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n612), .A2(new_n693), .ZN(new_n699));
  INV_X1    g0499(.A(new_n693), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n606), .A2(new_n611), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n643), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n699), .B1(new_n702), .B2(new_n612), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n682), .A2(new_n693), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n699), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n704), .A2(new_n706), .ZN(G399));
  NAND3_X1  g0507(.A1(new_n209), .A2(KEYINPUT94), .A3(new_n264), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(KEYINPUT94), .B1(new_n209), .B2(new_n264), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n711), .A2(new_n269), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n714), .B1(new_n213), .B2(new_n711), .ZN(new_n715));
  XOR2_X1   g0515(.A(KEYINPUT95), .B(KEYINPUT28), .Z(new_n716));
  XNOR2_X1  g0516(.A(new_n715), .B(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(G330), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT31), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n591), .A2(new_n326), .A3(new_n554), .A4(new_n628), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(new_n530), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n586), .B1(new_n590), .B2(new_n274), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n626), .A2(G179), .A3(new_n491), .A4(new_n627), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n722), .A2(new_n723), .A3(new_n554), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n724), .B1(new_n536), .B2(new_n537), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT30), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n721), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI211_X1 g0527(.A(KEYINPUT30), .B(new_n724), .C1(new_n536), .C2(new_n537), .ZN(new_n728));
  AOI211_X1 g0528(.A(new_n719), .B(new_n700), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n725), .A2(new_n726), .ZN(new_n730));
  INV_X1    g0530(.A(new_n721), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n730), .A2(new_n728), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(KEYINPUT31), .B1(new_n732), .B2(new_n693), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n651), .A2(new_n636), .A3(new_n693), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n735), .A2(new_n534), .A3(new_n543), .A4(new_n574), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n718), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n671), .A2(new_n669), .ZN(new_n738));
  INV_X1    g0538(.A(new_n574), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n678), .B1(new_n739), .B2(new_n542), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(new_n677), .B2(new_n678), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n742), .A2(KEYINPUT29), .A3(new_n700), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n700), .B1(new_n679), .B2(new_n672), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT29), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n737), .B1(new_n743), .B2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n717), .B1(new_n748), .B2(new_n269), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT96), .ZN(G364));
  AOI21_X1  g0550(.A(new_n269), .B1(new_n683), .B2(G45), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n711), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n698), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n754), .B1(G330), .B2(new_n696), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n339), .A2(new_n209), .ZN(new_n756));
  INV_X1    g0556(.A(G355), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n756), .A2(new_n757), .B1(G116), .B2(new_n209), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n245), .A2(G45), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n253), .A2(new_n209), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n760), .B1(new_n265), .B2(new_n213), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n758), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G13), .A2(G33), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(G20), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n214), .B1(G20), .B2(new_n375), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n753), .B1(new_n762), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(G20), .A2(G179), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n770), .A2(new_n367), .A3(G200), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G322), .ZN(new_n772));
  NOR3_X1   g0572(.A1(new_n770), .A2(new_n367), .A3(new_n281), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G326), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n772), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n770), .ZN(new_n777));
  NOR2_X1   g0577(.A1(G190), .A2(G200), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n339), .B(new_n776), .C1(G311), .C2(new_n780), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n326), .A2(new_n281), .A3(G190), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G20), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G294), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n770), .A2(new_n281), .A3(G190), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  XNOR2_X1  g0586(.A(KEYINPUT33), .B(G317), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT98), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n789), .B1(new_n788), .B2(new_n787), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n215), .A2(G179), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n791), .A2(G190), .A3(G200), .ZN(new_n792));
  INV_X1    g0592(.A(G303), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n791), .A2(new_n778), .ZN(new_n794));
  INV_X1    g0594(.A(G329), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n792), .A2(new_n793), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n791), .A2(new_n367), .A3(G200), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n796), .B1(G283), .B2(new_n798), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n781), .A2(new_n784), .A3(new_n790), .A4(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n783), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n204), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(G68), .B2(new_n785), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT97), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n792), .A2(new_n221), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n774), .A2(new_n295), .B1(new_n779), .B2(new_n202), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n805), .B(new_n806), .C1(G58), .C2(new_n771), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT32), .ZN(new_n808));
  INV_X1    g0608(.A(new_n794), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n808), .B1(new_n809), .B2(G159), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n339), .B1(new_n797), .B2(new_n205), .ZN(new_n811));
  NOR3_X1   g0611(.A1(new_n794), .A2(KEYINPUT32), .A3(new_n347), .ZN(new_n812));
  NOR3_X1   g0612(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n807), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n800), .B1(new_n804), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n769), .B1(new_n815), .B2(new_n766), .ZN(new_n816));
  INV_X1    g0616(.A(new_n765), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n816), .B1(new_n696), .B2(new_n817), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n755), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(G396));
  AND2_X1   g0620(.A1(new_n399), .A2(new_n693), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n656), .A2(new_n821), .A3(new_n657), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n412), .B2(new_n821), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n744), .A2(new_n824), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n823), .B(new_n700), .C1(new_n679), .C2(new_n672), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n732), .A2(new_n693), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n719), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n732), .A2(KEYINPUT31), .A3(new_n693), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n736), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(G330), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n827), .A2(new_n832), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT101), .Z(new_n834));
  AOI21_X1  g0634(.A(new_n753), .B1(new_n827), .B2(new_n832), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n753), .ZN(new_n837));
  INV_X1    g0637(.A(new_n766), .ZN(new_n838));
  INV_X1    g0638(.A(G283), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n774), .A2(new_n793), .B1(new_n786), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(G116), .B2(new_n780), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n841), .B(KEYINPUT99), .Z(new_n842));
  AOI22_X1  g0642(.A1(new_n809), .A2(G311), .B1(G294), .B2(new_n771), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n205), .B2(new_n792), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n253), .B1(new_n797), .B2(new_n221), .ZN(new_n845));
  OR4_X1    g0645(.A1(new_n802), .A2(new_n842), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  AOI22_X1  g0646(.A1(G137), .A2(new_n773), .B1(new_n785), .B2(G150), .ZN(new_n847));
  INV_X1    g0647(.A(G143), .ZN(new_n848));
  INV_X1    g0648(.A(new_n771), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n847), .B1(new_n848), .B2(new_n849), .C1(new_n347), .C2(new_n779), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n850), .B(KEYINPUT100), .Z(new_n851));
  OR2_X1    g0651(.A1(new_n851), .A2(KEYINPUT34), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(KEYINPUT34), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n339), .B1(new_n792), .B2(new_n295), .ZN(new_n854));
  INV_X1    g0654(.A(G132), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n797), .A2(new_n219), .B1(new_n794), .B2(new_n855), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n854), .B(new_n856), .C1(G58), .C2(new_n783), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n852), .A2(new_n853), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n838), .B1(new_n846), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n766), .A2(new_n763), .ZN(new_n860));
  AOI211_X1 g0660(.A(new_n837), .B(new_n859), .C1(new_n202), .C2(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(new_n823), .B2(new_n764), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n836), .A2(new_n862), .ZN(G384));
  NAND2_X1  g0663(.A1(new_n508), .A2(new_n510), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT35), .ZN(new_n865));
  OAI211_X1 g0665(.A(G116), .B(new_n216), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(new_n865), .B2(new_n864), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(KEYINPUT36), .ZN(new_n868));
  OAI21_X1  g0668(.A(G77), .B1(new_n343), .B2(new_n219), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n869), .A2(new_n212), .B1(G50), .B2(new_n219), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n298), .A2(G13), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n868), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n688), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n654), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n408), .A2(new_n693), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n826), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n693), .A2(new_n427), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n450), .A2(new_n459), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n457), .B1(new_n452), .B2(new_n454), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n442), .A2(new_n444), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n881), .A2(new_n448), .A3(new_n447), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n427), .B(new_n693), .C1(new_n880), .C2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n877), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT38), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT37), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n382), .A2(new_n292), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n349), .B1(new_n341), .B2(G68), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n889), .A2(KEYINPUT16), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n331), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n891), .A2(new_n688), .B1(new_n355), .B2(new_n369), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n380), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n887), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n380), .B1(new_n383), .B2(new_n332), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n688), .B1(new_n383), .B2(new_n332), .ZN(new_n896));
  AND4_X1   g0696(.A1(new_n887), .A2(new_n895), .A3(new_n896), .A4(new_n370), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n891), .A2(new_n688), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n899), .B1(new_n653), .B2(new_n663), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n886), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT102), .ZN(new_n902));
  INV_X1    g0702(.A(new_n899), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n386), .A2(new_n903), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n904), .B(KEYINPUT38), .C1(new_n897), .C2(new_n894), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n901), .A2(new_n902), .A3(new_n905), .ZN(new_n906));
  OAI211_X1 g0706(.A(KEYINPUT102), .B(new_n886), .C1(new_n898), .C2(new_n900), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n874), .B1(new_n885), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT103), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n450), .A2(new_n693), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT39), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n895), .A2(new_n896), .A3(new_n370), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(KEYINPUT37), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n895), .A2(new_n896), .A3(new_n887), .A4(new_n370), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n896), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n386), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT38), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT104), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n921), .A2(new_n922), .A3(new_n905), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n913), .B1(new_n908), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n921), .A2(new_n905), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n925), .A2(new_n922), .A3(KEYINPUT39), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n912), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  OAI211_X1 g0727(.A(KEYINPUT103), .B(new_n874), .C1(new_n885), .C2(new_n908), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n911), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n743), .A2(new_n746), .A3(new_n465), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT105), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n743), .A2(new_n746), .A3(new_n465), .A4(KEYINPUT105), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n667), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n929), .B(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT40), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n831), .A2(new_n823), .A3(new_n884), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n937), .B1(new_n908), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n884), .A2(new_n823), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(new_n736), .B2(new_n734), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n937), .B1(new_n921), .B2(new_n905), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n939), .A2(new_n943), .ZN(new_n944));
  AND2_X1   g0744(.A1(new_n465), .A2(new_n831), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n718), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n944), .B2(new_n945), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n936), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n298), .B2(new_n683), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n936), .A2(new_n947), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n872), .B1(new_n949), .B2(new_n950), .ZN(G367));
  NAND2_X1  g0751(.A1(new_n693), .A2(new_n522), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n539), .A2(new_n542), .A3(new_n952), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n953), .A2(new_n612), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n693), .B1(new_n954), .B2(new_n542), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n703), .A2(new_n705), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n540), .A2(new_n541), .A3(new_n693), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n953), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n955), .B1(KEYINPUT42), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(KEYINPUT42), .B2(new_n960), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n693), .A2(new_n568), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n574), .B(new_n963), .Z(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n962), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n967), .B(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n959), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n704), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n969), .B(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n699), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n956), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT45), .ZN(new_n975));
  NOR3_X1   g0775(.A1(new_n974), .A2(new_n970), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(KEYINPUT45), .B1(new_n706), .B2(new_n959), .ZN(new_n977));
  AOI21_X1  g0777(.A(KEYINPUT44), .B1(new_n974), .B2(new_n970), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT44), .ZN(new_n979));
  NOR3_X1   g0779(.A1(new_n706), .A2(new_n959), .A3(new_n979), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n976), .A2(new_n977), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(KEYINPUT106), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n704), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n703), .A2(new_n705), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n957), .A2(new_n984), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(new_n697), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n981), .A2(KEYINPUT106), .A3(new_n698), .A4(new_n703), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n983), .A2(new_n747), .A3(new_n986), .A4(new_n987), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n988), .A2(new_n747), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n711), .B(KEYINPUT41), .Z(new_n990));
  OAI21_X1  g0790(.A(new_n751), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n972), .A2(new_n991), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n767), .B1(new_n209), .B2(new_n392), .C1(new_n237), .C2(new_n760), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n753), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT107), .Z(new_n995));
  INV_X1    g0795(.A(G137), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n774), .A2(new_n848), .B1(new_n794), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(G150), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n849), .A2(new_n998), .B1(new_n779), .B2(new_n295), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n783), .A2(G68), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n792), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n253), .B1(new_n1002), .B2(G58), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n798), .A2(G77), .B1(new_n785), .B2(G159), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n1000), .A2(new_n1001), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(KEYINPUT46), .B1(new_n1002), .B2(G116), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n339), .B(new_n1006), .C1(G294), .C2(new_n785), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n797), .A2(new_n204), .ZN(new_n1008));
  INV_X1    g0808(.A(G317), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n849), .A2(new_n793), .B1(new_n794), .B2(new_n1009), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1008), .B(new_n1010), .C1(G311), .C2(new_n773), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1002), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1007), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n780), .A2(G283), .B1(new_n783), .B2(G107), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT108), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1005), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  AND2_X1   g0817(.A1(new_n1017), .A2(KEYINPUT47), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n766), .B1(new_n1017), .B2(KEYINPUT47), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n995), .B1(new_n1018), .B2(new_n1019), .C1(new_n965), .C2(new_n817), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n992), .A2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT109), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(G387));
  INV_X1    g0823(.A(new_n711), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(new_n747), .B2(new_n986), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n747), .B2(new_n986), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n756), .A2(new_n712), .B1(G107), .B2(new_n209), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n234), .A2(new_n265), .ZN(new_n1028));
  AOI211_X1 g0828(.A(G45), .B(new_n713), .C1(G68), .C2(G77), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n285), .A2(G50), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT50), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n760), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1027), .B1(new_n1028), .B2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1008), .A2(new_n253), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n219), .B2(new_n779), .C1(new_n202), .C2(new_n792), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n774), .A2(new_n347), .B1(new_n794), .B2(new_n998), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n849), .A2(new_n295), .B1(new_n786), .B2(new_n285), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n801), .A2(new_n392), .ZN(new_n1038));
  NOR4_X1   g0838(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(G322), .A2(new_n773), .B1(new_n785), .B2(G311), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n793), .B2(new_n779), .C1(new_n1009), .C2(new_n849), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT48), .ZN(new_n1042));
  INV_X1    g0842(.A(G294), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n801), .A2(new_n839), .B1(new_n792), .B2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT110), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1042), .A2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g0846(.A(KEYINPUT111), .B(KEYINPUT49), .Z(new_n1047));
  XNOR2_X1  g0847(.A(new_n1046), .B(new_n1047), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1048), .A2(KEYINPUT112), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n253), .B1(new_n794), .B2(new_n775), .C1(new_n614), .C2(new_n797), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n1048), .B2(KEYINPUT112), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1039), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n753), .B1(new_n768), .B2(new_n1033), .C1(new_n1052), .C2(new_n838), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n703), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1053), .B1(new_n1054), .B2(new_n765), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n752), .B2(new_n986), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1026), .A2(new_n1056), .ZN(G393));
  XOR2_X1   g0857(.A(new_n981), .B(new_n704), .Z(new_n1058));
  NAND2_X1  g0858(.A1(new_n747), .A2(new_n986), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1060), .A2(new_n711), .A3(new_n988), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(KEYINPUT116), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT116), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1060), .A2(new_n988), .A3(new_n1063), .A4(new_n711), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n767), .B1(new_n204), .B2(new_n209), .C1(new_n242), .C2(new_n760), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n837), .B1(new_n1066), .B2(KEYINPUT113), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(KEYINPUT113), .B2(new_n1066), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n809), .A2(G322), .B1(G303), .B2(new_n785), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1069), .B1(new_n839), .B2(new_n792), .C1(new_n1043), .C2(new_n779), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G317), .A2(new_n773), .B1(new_n771), .B2(G311), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1071), .B(new_n1072), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n253), .B1(new_n797), .B2(new_n205), .C1(new_n801), .C2(new_n614), .ZN(new_n1074));
  NOR3_X1   g0874(.A1(new_n1070), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  OR2_X1    g0876(.A1(new_n1076), .A2(KEYINPUT115), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n801), .A2(new_n202), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n253), .B(new_n1078), .C1(G87), .C2(new_n798), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G150), .A2(new_n773), .B1(new_n771), .B2(G159), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT51), .Z(new_n1081));
  OAI22_X1  g0881(.A1(new_n786), .A2(new_n295), .B1(new_n779), .B2(new_n285), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n792), .A2(new_n219), .B1(new_n794), .B2(new_n848), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1079), .A2(new_n1081), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1076), .A2(KEYINPUT115), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1077), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1068), .B1(new_n766), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n959), .B2(new_n817), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n1058), .B2(new_n751), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1065), .A2(new_n1091), .ZN(G390));
  AND4_X1   g0892(.A1(G330), .A2(new_n831), .A3(new_n823), .A4(new_n884), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n912), .B1(new_n877), .B2(new_n884), .ZN(new_n1094));
  NOR3_X1   g0894(.A1(new_n924), .A2(new_n1094), .A3(new_n926), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n912), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n693), .B1(new_n738), .B2(new_n741), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n875), .B1(new_n1097), .B2(new_n823), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n884), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1096), .B(new_n925), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1093), .B1(new_n1095), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1093), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n898), .A2(new_n900), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n920), .B1(KEYINPUT38), .B2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1105), .A2(KEYINPUT104), .A3(new_n913), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n922), .A2(new_n1105), .B1(new_n906), .B2(new_n907), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1106), .B1(new_n1107), .B2(new_n913), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1103), .B(new_n1100), .C1(new_n1108), .C2(new_n1094), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1102), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(KEYINPUT118), .B1(new_n1110), .B2(new_n751), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT118), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1102), .A2(new_n1112), .A3(new_n752), .A4(new_n1109), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n884), .B1(new_n737), .B2(new_n823), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n877), .B1(new_n1115), .B2(new_n1093), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(KEYINPUT117), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1115), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1118), .A2(new_n1103), .A3(new_n1098), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT117), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1120), .B(new_n877), .C1(new_n1115), .C2(new_n1093), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1117), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n466), .A2(new_n832), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n666), .B(new_n1123), .C1(new_n932), .C2(new_n933), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1110), .A2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1102), .A2(new_n1122), .A3(new_n1109), .A4(new_n1124), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1126), .A2(new_n711), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n837), .B1(new_n285), .B2(new_n860), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(G107), .A2(new_n785), .B1(new_n771), .B2(G116), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1130), .B1(new_n204), .B2(new_n779), .C1(new_n839), .C2(new_n774), .ZN(new_n1131));
  NOR4_X1   g0931(.A1(new_n1131), .A2(new_n339), .A3(new_n805), .A4(new_n1078), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n797), .A2(new_n219), .B1(new_n794), .B2(new_n1043), .ZN(new_n1133));
  XOR2_X1   g0933(.A(new_n1133), .B(KEYINPUT120), .Z(new_n1134));
  NAND2_X1  g0934(.A1(new_n1002), .A2(G150), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT53), .ZN(new_n1136));
  XOR2_X1   g0936(.A(KEYINPUT54), .B(G143), .Z(new_n1137));
  AOI22_X1  g0937(.A1(new_n780), .A2(new_n1137), .B1(G137), .B2(new_n785), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(G128), .A2(new_n773), .B1(new_n771), .B2(G132), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1138), .B(new_n1139), .C1(new_n347), .C2(new_n801), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1136), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(G125), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n339), .B1(new_n794), .B2(new_n1142), .C1(new_n295), .C2(new_n797), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT119), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1132), .A2(new_n1134), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n1129), .B1(new_n838), .B2(new_n1145), .C1(new_n1108), .C2(new_n764), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1114), .A2(new_n1128), .A3(new_n1146), .ZN(G378));
  AND2_X1   g0947(.A1(new_n325), .A2(new_n329), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n873), .B1(new_n306), .B2(new_n301), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n325), .A2(new_n329), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n1149), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n1151), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1154), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n763), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n774), .A2(new_n1142), .B1(new_n779), .B2(new_n996), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(G128), .A2(new_n771), .B1(new_n785), .B2(G132), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n998), .B2(new_n801), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n1159), .B(new_n1161), .C1(new_n1002), .C2(new_n1137), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT59), .ZN(new_n1163));
  OR2_X1    g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1165));
  AOI211_X1 g0965(.A(G33), .B(G41), .C1(new_n798), .C2(G159), .ZN(new_n1166));
  INV_X1    g0966(.A(G124), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1166), .B1(new_n1167), .B2(new_n794), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT121), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1164), .A2(new_n1165), .A3(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n797), .A2(new_n343), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n774), .A2(new_n614), .B1(new_n786), .B2(new_n204), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1171), .B(new_n1172), .C1(G107), .C2(new_n771), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n253), .A2(new_n264), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n1002), .B2(G77), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(G283), .A2(new_n809), .B1(new_n780), .B2(new_n393), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1173), .A2(new_n1001), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT58), .ZN(new_n1178));
  AOI21_X1  g0978(.A(G50), .B1(new_n362), .B2(new_n264), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1177), .A2(new_n1178), .B1(new_n1174), .B2(new_n1179), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1170), .B(new_n1180), .C1(new_n1178), .C2(new_n1177), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n766), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n860), .A2(new_n295), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1158), .A2(new_n753), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n929), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n718), .B1(new_n941), .B2(new_n942), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n939), .A2(KEYINPUT122), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(KEYINPUT122), .B1(new_n939), .B2(new_n1187), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n1188), .A2(new_n1189), .A3(new_n1157), .ZN(new_n1190));
  AND4_X1   g0990(.A1(KEYINPUT122), .A2(new_n1157), .A3(new_n939), .A4(new_n1187), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1186), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1189), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n939), .A2(new_n1187), .A3(KEYINPUT122), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1157), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1188), .B1(new_n1189), .B2(new_n1157), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1196), .A2(new_n929), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1192), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1185), .B1(new_n1199), .B2(new_n752), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1127), .A2(new_n1124), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(KEYINPUT57), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n1196), .A2(new_n929), .A3(new_n1197), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n929), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1204));
  OAI21_X1  g1004(.A(KEYINPUT123), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT123), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1192), .A2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1202), .B1(new_n1205), .B2(new_n1207), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n1192), .A2(new_n1198), .B1(new_n1127), .B2(new_n1124), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n711), .B1(new_n1209), .B2(KEYINPUT57), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1200), .B1(new_n1208), .B2(new_n1210), .ZN(G375));
  NAND2_X1  g1011(.A1(new_n1099), .A2(new_n763), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n766), .A2(G68), .A3(new_n763), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n774), .A2(new_n1043), .B1(new_n794), .B2(new_n793), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n339), .B(new_n1214), .C1(G77), .C2(new_n798), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1038), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n780), .A2(G107), .B1(G116), .B2(new_n785), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n1002), .A2(G97), .B1(G283), .B2(new_n771), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n780), .A2(G150), .B1(new_n783), .B2(G50), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1220), .B(KEYINPUT124), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1171), .A2(new_n253), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1002), .A2(G159), .B1(new_n1137), .B2(new_n785), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n773), .A2(G132), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n809), .A2(G128), .B1(G137), .B2(new_n771), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .A4(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1219), .B1(new_n1221), .B2(new_n1226), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n837), .B(new_n1213), .C1(new_n1227), .C2(new_n766), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n1122), .A2(new_n752), .B1(new_n1212), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n990), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1125), .A2(new_n1230), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1229), .B1(new_n1231), .B2(new_n1232), .ZN(G381));
  INV_X1    g1033(.A(G378), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1026), .A2(new_n819), .A3(new_n1056), .ZN(new_n1235));
  NOR4_X1   g1035(.A1(G390), .A2(G381), .A3(G384), .A4(new_n1235), .ZN(new_n1236));
  AND3_X1   g1036(.A1(new_n1022), .A2(new_n1234), .A3(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT125), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1200), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT57), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1024), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1206), .B1(new_n1192), .B2(new_n1198), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1204), .A2(KEYINPUT123), .ZN(new_n1244));
  OAI211_X1 g1044(.A(KEYINPUT57), .B(new_n1201), .C1(new_n1243), .C2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1239), .B1(new_n1242), .B2(new_n1245), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n1237), .A2(new_n1238), .A3(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1238), .B1(new_n1237), .B2(new_n1246), .ZN(new_n1248));
  OR2_X1    g1048(.A1(new_n1247), .A2(new_n1248), .ZN(G407));
  OR3_X1    g1049(.A1(G375), .A2(G343), .A3(G378), .ZN(new_n1250));
  OAI211_X1 g1050(.A(G213), .B(new_n1250), .C1(new_n1247), .C2(new_n1248), .ZN(G409));
  OAI211_X1 g1051(.A(G378), .B(new_n1200), .C1(new_n1208), .C2(new_n1210), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1184), .B1(new_n1240), .B2(new_n990), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n751), .B1(new_n1205), .B2(new_n1207), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1234), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1252), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(G213), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1257), .A2(G343), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1123), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n934), .A2(new_n667), .A3(new_n1261), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1260), .A2(new_n1262), .A3(KEYINPUT60), .A4(new_n1117), .ZN(new_n1263));
  AND2_X1   g1063(.A1(new_n1263), .A2(new_n711), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT60), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1264), .B1(new_n1232), .B2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1267), .A2(G384), .A3(new_n1229), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1266), .A2(new_n1232), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1263), .A2(new_n711), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1229), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(G384), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1268), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1256), .A2(new_n1259), .A3(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(KEYINPUT62), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT61), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1258), .B1(new_n1252), .B2(new_n1255), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT62), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1279), .A2(new_n1280), .A3(new_n1275), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1258), .A2(G2897), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1268), .A2(new_n1273), .A3(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1282), .B1(new_n1268), .B2(new_n1273), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1185), .B1(new_n1209), .B2(new_n1230), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n752), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1288));
  AOI21_X1  g1088(.A(G378), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1289), .B1(new_n1246), .B2(G378), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1286), .B1(new_n1290), .B2(new_n1258), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1277), .A2(new_n1278), .A3(new_n1281), .A4(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(G393), .A2(G396), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n1235), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(G390), .A2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT109), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1294), .A2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1297), .A2(new_n1065), .A3(new_n1091), .ZN(new_n1298));
  AND3_X1   g1098(.A1(new_n1295), .A2(new_n1021), .A3(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1021), .B1(new_n1295), .B2(new_n1298), .ZN(new_n1300));
  OR2_X1    g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1292), .A2(new_n1301), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1282), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1274), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1283), .ZN(new_n1306));
  OAI211_X1 g1106(.A(new_n1303), .B(new_n1278), .C1(new_n1279), .C2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  AOI211_X1 g1108(.A(new_n1258), .B(new_n1274), .C1(new_n1252), .C2(new_n1255), .ZN(new_n1309));
  OAI21_X1  g1109(.A(KEYINPUT126), .B1(new_n1309), .B2(KEYINPUT63), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(KEYINPUT63), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT126), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT63), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1276), .A2(new_n1312), .A3(new_n1313), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1308), .A2(new_n1310), .A3(new_n1311), .A4(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1302), .A2(new_n1315), .ZN(G405));
  NOR2_X1   g1116(.A1(new_n1275), .A2(KEYINPUT127), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1301), .A2(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1303), .B1(KEYINPUT127), .B2(new_n1275), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(G375), .A2(new_n1234), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n1252), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1322), .B1(KEYINPUT127), .B2(new_n1275), .ZN(new_n1323));
  XNOR2_X1  g1123(.A(new_n1320), .B(new_n1323), .ZN(G402));
endmodule


