

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U556 ( .A1(n539), .A2(G2104), .ZN(n877) );
  INV_X1 U557 ( .A(KEYINPUT17), .ZN(n543) );
  XNOR2_X1 U558 ( .A(KEYINPUT23), .B(KEYINPUT65), .ZN(n550) );
  XNOR2_X1 U559 ( .A(n737), .B(n736), .ZN(n749) );
  NOR2_X1 U560 ( .A1(n735), .A2(n734), .ZN(n737) );
  XOR2_X1 U561 ( .A(KEYINPUT98), .B(n726), .Z(n771) );
  NOR2_X1 U562 ( .A1(G651), .A2(G543), .ZN(n656) );
  NOR2_X1 U563 ( .A1(n557), .A2(n556), .ZN(G160) );
  AND2_X1 U564 ( .A1(n779), .A2(n778), .ZN(n521) );
  NAND2_X1 U565 ( .A1(n794), .A2(n815), .ZN(n522) );
  NOR2_X1 U566 ( .A1(n704), .A2(n703), .ZN(n710) );
  INV_X1 U567 ( .A(KEYINPUT103), .ZN(n713) );
  XNOR2_X1 U568 ( .A(n714), .B(n713), .ZN(n717) );
  INV_X1 U569 ( .A(KEYINPUT104), .ZN(n736) );
  NAND2_X1 U570 ( .A1(n782), .A2(n692), .ZN(n738) );
  INV_X1 U571 ( .A(n771), .ZN(n776) );
  NOR2_X1 U572 ( .A1(G164), .A2(G1384), .ZN(n782) );
  AND2_X1 U573 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U574 ( .A(n582), .B(KEYINPUT76), .ZN(n583) );
  XNOR2_X1 U575 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U576 ( .A(n543), .B(KEYINPUT66), .ZN(n544) );
  NOR2_X1 U577 ( .A1(n522), .A2(n818), .ZN(n813) );
  NOR2_X1 U578 ( .A1(n647), .A2(n529), .ZN(n653) );
  NOR2_X2 U579 ( .A1(G2104), .A2(n539), .ZN(n873) );
  XNOR2_X1 U580 ( .A(n551), .B(n550), .ZN(n553) );
  NOR2_X1 U581 ( .A1(n549), .A2(n548), .ZN(G164) );
  INV_X1 U582 ( .A(G651), .ZN(n529) );
  NOR2_X1 U583 ( .A1(G543), .A2(n529), .ZN(n523) );
  XOR2_X2 U584 ( .A(KEYINPUT1), .B(n523), .Z(n655) );
  NAND2_X1 U585 ( .A1(G63), .A2(n655), .ZN(n526) );
  XNOR2_X1 U586 ( .A(G543), .B(KEYINPUT0), .ZN(n524) );
  XNOR2_X1 U587 ( .A(n524), .B(KEYINPUT67), .ZN(n647) );
  NOR2_X2 U588 ( .A1(G651), .A2(n647), .ZN(n659) );
  NAND2_X1 U589 ( .A1(G51), .A2(n659), .ZN(n525) );
  NAND2_X1 U590 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U591 ( .A(KEYINPUT6), .B(n527), .ZN(n534) );
  NAND2_X1 U592 ( .A1(n656), .A2(G89), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n528), .B(KEYINPUT4), .ZN(n531) );
  NAND2_X1 U594 ( .A1(G76), .A2(n653), .ZN(n530) );
  NAND2_X1 U595 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U596 ( .A(n532), .B(KEYINPUT5), .Z(n533) );
  NOR2_X1 U597 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U598 ( .A(KEYINPUT81), .B(n535), .Z(n536) );
  XOR2_X1 U599 ( .A(KEYINPUT7), .B(n536), .Z(G168) );
  XOR2_X1 U600 ( .A(G168), .B(KEYINPUT8), .Z(n537) );
  XNOR2_X1 U601 ( .A(KEYINPUT82), .B(n537), .ZN(G286) );
  INV_X1 U602 ( .A(G2105), .ZN(n539) );
  NAND2_X1 U603 ( .A1(G126), .A2(n873), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n538), .B(KEYINPUT92), .ZN(n542) );
  NAND2_X1 U605 ( .A1(G102), .A2(n877), .ZN(n540) );
  XOR2_X1 U606 ( .A(KEYINPUT93), .B(n540), .Z(n541) );
  NAND2_X1 U607 ( .A1(n542), .A2(n541), .ZN(n549) );
  NOR2_X1 U608 ( .A1(G2104), .A2(G2105), .ZN(n545) );
  XNOR2_X2 U609 ( .A(n545), .B(n544), .ZN(n621) );
  NAND2_X1 U610 ( .A1(G138), .A2(n621), .ZN(n547) );
  AND2_X1 U611 ( .A1(G2104), .A2(G2105), .ZN(n872) );
  NAND2_X1 U612 ( .A1(n872), .A2(G114), .ZN(n546) );
  NAND2_X1 U613 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U614 ( .A1(G101), .A2(n877), .ZN(n551) );
  NAND2_X1 U615 ( .A1(G113), .A2(n872), .ZN(n552) );
  NAND2_X1 U616 ( .A1(n553), .A2(n552), .ZN(n557) );
  NAND2_X1 U617 ( .A1(G137), .A2(n621), .ZN(n555) );
  NAND2_X1 U618 ( .A1(n873), .A2(G125), .ZN(n554) );
  NAND2_X1 U619 ( .A1(n555), .A2(n554), .ZN(n556) );
  AND2_X1 U620 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U621 ( .A(G132), .ZN(G219) );
  INV_X1 U622 ( .A(G82), .ZN(G220) );
  INV_X1 U623 ( .A(G120), .ZN(G236) );
  NAND2_X1 U624 ( .A1(G88), .A2(n656), .ZN(n559) );
  NAND2_X1 U625 ( .A1(G75), .A2(n653), .ZN(n558) );
  NAND2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n563) );
  NAND2_X1 U627 ( .A1(G62), .A2(n655), .ZN(n561) );
  NAND2_X1 U628 ( .A1(G50), .A2(n659), .ZN(n560) );
  NAND2_X1 U629 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U630 ( .A1(n563), .A2(n562), .ZN(G166) );
  XNOR2_X1 U631 ( .A(KEYINPUT71), .B(KEYINPUT72), .ZN(n568) );
  NAND2_X1 U632 ( .A1(G90), .A2(n656), .ZN(n565) );
  NAND2_X1 U633 ( .A1(G77), .A2(n653), .ZN(n564) );
  NAND2_X1 U634 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U635 ( .A(n566), .B(KEYINPUT9), .ZN(n567) );
  XNOR2_X1 U636 ( .A(n568), .B(n567), .ZN(n573) );
  NAND2_X1 U637 ( .A1(n655), .A2(G64), .ZN(n569) );
  XNOR2_X1 U638 ( .A(n569), .B(KEYINPUT70), .ZN(n571) );
  NAND2_X1 U639 ( .A1(G52), .A2(n659), .ZN(n570) );
  NAND2_X1 U640 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U641 ( .A1(n573), .A2(n572), .ZN(G171) );
  INV_X1 U642 ( .A(G171), .ZN(G301) );
  NAND2_X1 U643 ( .A1(G7), .A2(G661), .ZN(n574) );
  XNOR2_X1 U644 ( .A(n574), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U645 ( .A(G223), .ZN(n831) );
  NAND2_X1 U646 ( .A1(n831), .A2(G567), .ZN(n575) );
  XOR2_X1 U647 ( .A(KEYINPUT11), .B(n575), .Z(G234) );
  INV_X1 U648 ( .A(G860), .ZN(n610) );
  NAND2_X1 U649 ( .A1(n655), .A2(G56), .ZN(n576) );
  XNOR2_X1 U650 ( .A(n576), .B(KEYINPUT14), .ZN(n578) );
  NAND2_X1 U651 ( .A1(G43), .A2(n659), .ZN(n577) );
  NAND2_X1 U652 ( .A1(n578), .A2(n577), .ZN(n586) );
  NAND2_X1 U653 ( .A1(G68), .A2(n653), .ZN(n581) );
  NAND2_X1 U654 ( .A1(n656), .A2(G81), .ZN(n579) );
  XNOR2_X1 U655 ( .A(n579), .B(KEYINPUT12), .ZN(n580) );
  NAND2_X1 U656 ( .A1(n581), .A2(n580), .ZN(n584) );
  INV_X1 U657 ( .A(KEYINPUT13), .ZN(n582) );
  NOR2_X2 U658 ( .A1(n586), .A2(n585), .ZN(n960) );
  INV_X1 U659 ( .A(n960), .ZN(n614) );
  NOR2_X1 U660 ( .A1(n610), .A2(n614), .ZN(n587) );
  XNOR2_X1 U661 ( .A(n587), .B(KEYINPUT77), .ZN(G153) );
  NAND2_X1 U662 ( .A1(G868), .A2(G301), .ZN(n599) );
  NAND2_X1 U663 ( .A1(G79), .A2(n653), .ZN(n596) );
  NAND2_X1 U664 ( .A1(G54), .A2(n659), .ZN(n588) );
  XNOR2_X1 U665 ( .A(n588), .B(KEYINPUT80), .ZN(n591) );
  NAND2_X1 U666 ( .A1(G92), .A2(n656), .ZN(n589) );
  XOR2_X1 U667 ( .A(KEYINPUT79), .B(n589), .Z(n590) );
  NAND2_X1 U668 ( .A1(n591), .A2(n590), .ZN(n594) );
  NAND2_X1 U669 ( .A1(n655), .A2(G66), .ZN(n592) );
  XOR2_X1 U670 ( .A(KEYINPUT78), .B(n592), .Z(n593) );
  NOR2_X1 U671 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U672 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X2 U673 ( .A(n597), .B(KEYINPUT15), .ZN(n898) );
  INV_X1 U674 ( .A(n898), .ZN(n951) );
  INV_X1 U675 ( .A(G868), .ZN(n673) );
  NAND2_X1 U676 ( .A1(n951), .A2(n673), .ZN(n598) );
  NAND2_X1 U677 ( .A1(n599), .A2(n598), .ZN(G284) );
  NAND2_X1 U678 ( .A1(G65), .A2(n655), .ZN(n600) );
  XOR2_X1 U679 ( .A(KEYINPUT74), .B(n600), .Z(n605) );
  NAND2_X1 U680 ( .A1(G91), .A2(n656), .ZN(n602) );
  NAND2_X1 U681 ( .A1(G78), .A2(n653), .ZN(n601) );
  NAND2_X1 U682 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U683 ( .A(KEYINPUT73), .B(n603), .Z(n604) );
  NOR2_X1 U684 ( .A1(n605), .A2(n604), .ZN(n607) );
  NAND2_X1 U685 ( .A1(n659), .A2(G53), .ZN(n606) );
  NAND2_X1 U686 ( .A1(n607), .A2(n606), .ZN(G299) );
  NAND2_X1 U687 ( .A1(G868), .A2(G286), .ZN(n609) );
  NAND2_X1 U688 ( .A1(G299), .A2(n673), .ZN(n608) );
  NAND2_X1 U689 ( .A1(n609), .A2(n608), .ZN(G297) );
  NAND2_X1 U690 ( .A1(n610), .A2(G559), .ZN(n611) );
  NAND2_X1 U691 ( .A1(n611), .A2(n898), .ZN(n612) );
  XNOR2_X1 U692 ( .A(n612), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U693 ( .A1(n898), .A2(G868), .ZN(n613) );
  NOR2_X1 U694 ( .A1(G559), .A2(n613), .ZN(n616) );
  NOR2_X1 U695 ( .A1(G868), .A2(n614), .ZN(n615) );
  NOR2_X1 U696 ( .A1(n616), .A2(n615), .ZN(G282) );
  NAND2_X1 U697 ( .A1(G111), .A2(n872), .ZN(n626) );
  NAND2_X1 U698 ( .A1(G123), .A2(n873), .ZN(n617) );
  XNOR2_X1 U699 ( .A(n617), .B(KEYINPUT18), .ZN(n620) );
  NAND2_X1 U700 ( .A1(G99), .A2(n877), .ZN(n618) );
  XNOR2_X1 U701 ( .A(n618), .B(KEYINPUT84), .ZN(n619) );
  NAND2_X1 U702 ( .A1(n620), .A2(n619), .ZN(n624) );
  NAND2_X1 U703 ( .A1(G135), .A2(n621), .ZN(n622) );
  XNOR2_X1 U704 ( .A(KEYINPUT83), .B(n622), .ZN(n623) );
  NOR2_X1 U705 ( .A1(n624), .A2(n623), .ZN(n625) );
  NAND2_X1 U706 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U707 ( .A(n627), .B(KEYINPUT85), .ZN(n999) );
  XOR2_X1 U708 ( .A(G2096), .B(n999), .Z(n628) );
  NOR2_X1 U709 ( .A1(G2100), .A2(n628), .ZN(n629) );
  XOR2_X1 U710 ( .A(KEYINPUT86), .B(n629), .Z(G156) );
  NAND2_X1 U711 ( .A1(G67), .A2(n655), .ZN(n631) );
  NAND2_X1 U712 ( .A1(G55), .A2(n659), .ZN(n630) );
  NAND2_X1 U713 ( .A1(n631), .A2(n630), .ZN(n635) );
  NAND2_X1 U714 ( .A1(G93), .A2(n656), .ZN(n633) );
  NAND2_X1 U715 ( .A1(G80), .A2(n653), .ZN(n632) );
  NAND2_X1 U716 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U717 ( .A1(n635), .A2(n634), .ZN(n674) );
  NAND2_X1 U718 ( .A1(n898), .A2(G559), .ZN(n671) );
  XOR2_X1 U719 ( .A(n960), .B(n671), .Z(n636) );
  NOR2_X1 U720 ( .A1(G860), .A2(n636), .ZN(n637) );
  XNOR2_X1 U721 ( .A(n674), .B(n637), .ZN(G145) );
  NAND2_X1 U722 ( .A1(n655), .A2(G61), .ZN(n638) );
  XOR2_X1 U723 ( .A(KEYINPUT87), .B(n638), .Z(n640) );
  NAND2_X1 U724 ( .A1(n656), .A2(G86), .ZN(n639) );
  NAND2_X1 U725 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U726 ( .A(KEYINPUT88), .B(n641), .ZN(n644) );
  NAND2_X1 U727 ( .A1(G73), .A2(n653), .ZN(n642) );
  XOR2_X1 U728 ( .A(KEYINPUT2), .B(n642), .Z(n643) );
  NOR2_X1 U729 ( .A1(n644), .A2(n643), .ZN(n646) );
  NAND2_X1 U730 ( .A1(n659), .A2(G48), .ZN(n645) );
  NAND2_X1 U731 ( .A1(n646), .A2(n645), .ZN(G305) );
  NAND2_X1 U732 ( .A1(G49), .A2(n659), .ZN(n649) );
  NAND2_X1 U733 ( .A1(G87), .A2(n647), .ZN(n648) );
  NAND2_X1 U734 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U735 ( .A1(n655), .A2(n650), .ZN(n652) );
  NAND2_X1 U736 ( .A1(G651), .A2(G74), .ZN(n651) );
  NAND2_X1 U737 ( .A1(n652), .A2(n651), .ZN(G288) );
  NAND2_X1 U738 ( .A1(G72), .A2(n653), .ZN(n654) );
  XNOR2_X1 U739 ( .A(n654), .B(KEYINPUT68), .ZN(n664) );
  NAND2_X1 U740 ( .A1(G60), .A2(n655), .ZN(n658) );
  NAND2_X1 U741 ( .A1(G85), .A2(n656), .ZN(n657) );
  NAND2_X1 U742 ( .A1(n658), .A2(n657), .ZN(n662) );
  NAND2_X1 U743 ( .A1(G47), .A2(n659), .ZN(n660) );
  XNOR2_X1 U744 ( .A(KEYINPUT69), .B(n660), .ZN(n661) );
  NOR2_X1 U745 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U746 ( .A1(n664), .A2(n663), .ZN(G290) );
  INV_X1 U747 ( .A(G299), .ZN(n943) );
  XNOR2_X1 U748 ( .A(KEYINPUT19), .B(G288), .ZN(n665) );
  XNOR2_X1 U749 ( .A(n665), .B(G290), .ZN(n666) );
  XOR2_X1 U750 ( .A(n674), .B(n666), .Z(n668) );
  XNOR2_X1 U751 ( .A(n960), .B(G166), .ZN(n667) );
  XNOR2_X1 U752 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U753 ( .A(n943), .B(n669), .ZN(n670) );
  XNOR2_X1 U754 ( .A(G305), .B(n670), .ZN(n897) );
  XOR2_X1 U755 ( .A(n897), .B(n671), .Z(n672) );
  NOR2_X1 U756 ( .A1(n673), .A2(n672), .ZN(n676) );
  NOR2_X1 U757 ( .A1(G868), .A2(n674), .ZN(n675) );
  NOR2_X1 U758 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U759 ( .A(KEYINPUT89), .B(n677), .ZN(G295) );
  NAND2_X1 U760 ( .A1(G2078), .A2(G2084), .ZN(n678) );
  XOR2_X1 U761 ( .A(KEYINPUT20), .B(n678), .Z(n679) );
  NAND2_X1 U762 ( .A1(G2090), .A2(n679), .ZN(n680) );
  XNOR2_X1 U763 ( .A(KEYINPUT21), .B(n680), .ZN(n681) );
  NAND2_X1 U764 ( .A1(n681), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U765 ( .A(KEYINPUT75), .B(G57), .ZN(G237) );
  XNOR2_X1 U766 ( .A(KEYINPUT90), .B(G44), .ZN(n682) );
  XNOR2_X1 U767 ( .A(n682), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U768 ( .A1(G237), .A2(G236), .ZN(n683) );
  NAND2_X1 U769 ( .A1(G69), .A2(n683), .ZN(n684) );
  XNOR2_X1 U770 ( .A(KEYINPUT91), .B(n684), .ZN(n685) );
  NAND2_X1 U771 ( .A1(n685), .A2(G108), .ZN(n836) );
  NAND2_X1 U772 ( .A1(n836), .A2(G567), .ZN(n690) );
  NOR2_X1 U773 ( .A1(G220), .A2(G219), .ZN(n686) );
  XOR2_X1 U774 ( .A(KEYINPUT22), .B(n686), .Z(n687) );
  NOR2_X1 U775 ( .A1(G218), .A2(n687), .ZN(n688) );
  NAND2_X1 U776 ( .A1(G96), .A2(n688), .ZN(n837) );
  NAND2_X1 U777 ( .A1(n837), .A2(G2106), .ZN(n689) );
  NAND2_X1 U778 ( .A1(n690), .A2(n689), .ZN(n838) );
  NAND2_X1 U779 ( .A1(G483), .A2(G661), .ZN(n691) );
  NOR2_X1 U780 ( .A1(n838), .A2(n691), .ZN(n835) );
  NAND2_X1 U781 ( .A1(n835), .A2(G36), .ZN(G176) );
  INV_X1 U782 ( .A(G166), .ZN(G303) );
  INV_X1 U783 ( .A(KEYINPUT100), .ZN(n697) );
  NAND2_X1 U784 ( .A1(G160), .A2(G40), .ZN(n781) );
  INV_X1 U785 ( .A(n781), .ZN(n692) );
  NAND2_X1 U786 ( .A1(G1956), .A2(n738), .ZN(n695) );
  AND2_X1 U787 ( .A1(n692), .A2(n782), .ZN(n699) );
  NAND2_X1 U788 ( .A1(n699), .A2(G2072), .ZN(n693) );
  XOR2_X1 U789 ( .A(KEYINPUT27), .B(n693), .Z(n694) );
  NAND2_X1 U790 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U791 ( .A(n697), .B(n696), .ZN(n715) );
  NOR2_X1 U792 ( .A1(n943), .A2(n715), .ZN(n698) );
  XOR2_X1 U793 ( .A(n698), .B(KEYINPUT28), .Z(n719) );
  NAND2_X1 U794 ( .A1(n699), .A2(G1996), .ZN(n700) );
  XNOR2_X1 U795 ( .A(n700), .B(KEYINPUT26), .ZN(n701) );
  NAND2_X1 U796 ( .A1(n701), .A2(n960), .ZN(n704) );
  NAND2_X1 U797 ( .A1(G1341), .A2(n738), .ZN(n702) );
  XNOR2_X1 U798 ( .A(n702), .B(KEYINPUT101), .ZN(n703) );
  NAND2_X1 U799 ( .A1(n710), .A2(n898), .ZN(n708) );
  NOR2_X1 U800 ( .A1(n699), .A2(G1348), .ZN(n706) );
  NOR2_X1 U801 ( .A1(G2067), .A2(n738), .ZN(n705) );
  NOR2_X1 U802 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U803 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U804 ( .A(n709), .B(KEYINPUT102), .ZN(n712) );
  OR2_X1 U805 ( .A1(n710), .A2(n898), .ZN(n711) );
  NAND2_X1 U806 ( .A1(n712), .A2(n711), .ZN(n714) );
  NAND2_X1 U807 ( .A1(n943), .A2(n715), .ZN(n716) );
  NAND2_X1 U808 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U809 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U810 ( .A(n720), .B(KEYINPUT29), .ZN(n725) );
  NOR2_X1 U811 ( .A1(n699), .A2(G1961), .ZN(n721) );
  XOR2_X1 U812 ( .A(KEYINPUT99), .B(n721), .Z(n723) );
  XOR2_X1 U813 ( .A(G2078), .B(KEYINPUT25), .Z(n929) );
  NOR2_X1 U814 ( .A1(n929), .A2(n738), .ZN(n722) );
  NOR2_X1 U815 ( .A1(n723), .A2(n722), .ZN(n730) );
  NOR2_X1 U816 ( .A1(G301), .A2(n730), .ZN(n724) );
  NOR2_X1 U817 ( .A1(n725), .A2(n724), .ZN(n735) );
  NAND2_X1 U818 ( .A1(n738), .A2(G8), .ZN(n726) );
  NOR2_X1 U819 ( .A1(n776), .A2(G1966), .ZN(n751) );
  NOR2_X1 U820 ( .A1(G2084), .A2(n738), .ZN(n748) );
  NOR2_X1 U821 ( .A1(n751), .A2(n748), .ZN(n727) );
  NAND2_X1 U822 ( .A1(G8), .A2(n727), .ZN(n728) );
  XNOR2_X1 U823 ( .A(KEYINPUT30), .B(n728), .ZN(n729) );
  NOR2_X1 U824 ( .A1(G168), .A2(n729), .ZN(n732) );
  AND2_X1 U825 ( .A1(G301), .A2(n730), .ZN(n731) );
  NOR2_X1 U826 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U827 ( .A(n733), .B(KEYINPUT31), .ZN(n734) );
  NAND2_X1 U828 ( .A1(n749), .A2(G286), .ZN(n744) );
  NOR2_X1 U829 ( .A1(n776), .A2(G1971), .ZN(n740) );
  NOR2_X1 U830 ( .A1(G2090), .A2(n738), .ZN(n739) );
  NOR2_X1 U831 ( .A1(n740), .A2(n739), .ZN(n741) );
  XOR2_X1 U832 ( .A(KEYINPUT105), .B(n741), .Z(n742) );
  NAND2_X1 U833 ( .A1(n742), .A2(G303), .ZN(n743) );
  NAND2_X1 U834 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U835 ( .A(n745), .B(KEYINPUT106), .ZN(n746) );
  NAND2_X1 U836 ( .A1(n746), .A2(G8), .ZN(n747) );
  XNOR2_X1 U837 ( .A(n747), .B(KEYINPUT32), .ZN(n755) );
  NAND2_X1 U838 ( .A1(G8), .A2(n748), .ZN(n753) );
  INV_X1 U839 ( .A(n749), .ZN(n750) );
  NOR2_X1 U840 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U841 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U842 ( .A1(n755), .A2(n754), .ZN(n775) );
  NOR2_X1 U843 ( .A1(G1971), .A2(G303), .ZN(n756) );
  XNOR2_X1 U844 ( .A(KEYINPUT107), .B(n756), .ZN(n757) );
  NOR2_X1 U845 ( .A1(G1976), .A2(G288), .ZN(n944) );
  NAND2_X1 U846 ( .A1(n944), .A2(n771), .ZN(n763) );
  AND2_X1 U847 ( .A1(n757), .A2(n763), .ZN(n758) );
  NAND2_X1 U848 ( .A1(n775), .A2(n758), .ZN(n760) );
  NAND2_X1 U849 ( .A1(G1976), .A2(G288), .ZN(n945) );
  AND2_X1 U850 ( .A1(n945), .A2(n771), .ZN(n759) );
  NAND2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U852 ( .A(n761), .B(KEYINPUT64), .ZN(n762) );
  INV_X1 U853 ( .A(KEYINPUT33), .ZN(n764) );
  NAND2_X1 U854 ( .A1(n762), .A2(n764), .ZN(n769) );
  NOR2_X1 U855 ( .A1(n764), .A2(n763), .ZN(n765) );
  XOR2_X1 U856 ( .A(n765), .B(KEYINPUT108), .Z(n767) );
  XNOR2_X1 U857 ( .A(G1981), .B(G305), .ZN(n941) );
  INV_X1 U858 ( .A(n941), .ZN(n766) );
  NAND2_X1 U859 ( .A1(n769), .A2(n768), .ZN(n780) );
  NOR2_X1 U860 ( .A1(G1981), .A2(G305), .ZN(n770) );
  XNOR2_X1 U861 ( .A(KEYINPUT24), .B(n770), .ZN(n772) );
  NAND2_X1 U862 ( .A1(n772), .A2(n771), .ZN(n779) );
  NOR2_X1 U863 ( .A1(G2090), .A2(G303), .ZN(n773) );
  NAND2_X1 U864 ( .A1(G8), .A2(n773), .ZN(n774) );
  NAND2_X1 U865 ( .A1(n775), .A2(n774), .ZN(n777) );
  NAND2_X1 U866 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U867 ( .A1(n780), .A2(n521), .ZN(n814) );
  XNOR2_X1 U868 ( .A(G1986), .B(G290), .ZN(n958) );
  NOR2_X1 U869 ( .A1(n782), .A2(n781), .ZN(n823) );
  NAND2_X1 U870 ( .A1(n958), .A2(n823), .ZN(n794) );
  XOR2_X1 U871 ( .A(KEYINPUT37), .B(G2067), .Z(n822) );
  NAND2_X1 U872 ( .A1(G140), .A2(n621), .ZN(n783) );
  XNOR2_X1 U873 ( .A(n783), .B(KEYINPUT94), .ZN(n785) );
  NAND2_X1 U874 ( .A1(G104), .A2(n877), .ZN(n784) );
  NAND2_X1 U875 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U876 ( .A(KEYINPUT34), .B(n786), .ZN(n792) );
  NAND2_X1 U877 ( .A1(G116), .A2(n872), .ZN(n788) );
  NAND2_X1 U878 ( .A1(G128), .A2(n873), .ZN(n787) );
  NAND2_X1 U879 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U880 ( .A(KEYINPUT95), .B(n789), .ZN(n790) );
  XNOR2_X1 U881 ( .A(KEYINPUT35), .B(n790), .ZN(n791) );
  NOR2_X1 U882 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U883 ( .A(KEYINPUT36), .B(n793), .Z(n893) );
  AND2_X1 U884 ( .A1(n822), .A2(n893), .ZN(n1008) );
  NAND2_X1 U885 ( .A1(n1008), .A2(n823), .ZN(n815) );
  NAND2_X1 U886 ( .A1(G95), .A2(n877), .ZN(n796) );
  NAND2_X1 U887 ( .A1(G107), .A2(n872), .ZN(n795) );
  NAND2_X1 U888 ( .A1(n796), .A2(n795), .ZN(n800) );
  NAND2_X1 U889 ( .A1(n873), .A2(G119), .ZN(n798) );
  NAND2_X1 U890 ( .A1(G131), .A2(n621), .ZN(n797) );
  NAND2_X1 U891 ( .A1(n798), .A2(n797), .ZN(n799) );
  OR2_X1 U892 ( .A1(n800), .A2(n799), .ZN(n886) );
  NAND2_X1 U893 ( .A1(G1991), .A2(n886), .ZN(n801) );
  XOR2_X1 U894 ( .A(KEYINPUT96), .B(n801), .Z(n811) );
  NAND2_X1 U895 ( .A1(G105), .A2(n877), .ZN(n802) );
  XNOR2_X1 U896 ( .A(n802), .B(KEYINPUT38), .ZN(n809) );
  NAND2_X1 U897 ( .A1(G117), .A2(n872), .ZN(n804) );
  NAND2_X1 U898 ( .A1(G129), .A2(n873), .ZN(n803) );
  NAND2_X1 U899 ( .A1(n804), .A2(n803), .ZN(n807) );
  NAND2_X1 U900 ( .A1(G141), .A2(n621), .ZN(n805) );
  XNOR2_X1 U901 ( .A(KEYINPUT97), .B(n805), .ZN(n806) );
  NOR2_X1 U902 ( .A1(n807), .A2(n806), .ZN(n808) );
  NAND2_X1 U903 ( .A1(n809), .A2(n808), .ZN(n885) );
  AND2_X1 U904 ( .A1(G1996), .A2(n885), .ZN(n810) );
  NOR2_X1 U905 ( .A1(n811), .A2(n810), .ZN(n1001) );
  INV_X1 U906 ( .A(n823), .ZN(n812) );
  NOR2_X1 U907 ( .A1(n1001), .A2(n812), .ZN(n818) );
  NAND2_X1 U908 ( .A1(n814), .A2(n813), .ZN(n829) );
  INV_X1 U909 ( .A(n815), .ZN(n827) );
  NOR2_X1 U910 ( .A1(G1996), .A2(n885), .ZN(n1005) );
  NOR2_X1 U911 ( .A1(G1986), .A2(G290), .ZN(n816) );
  NOR2_X1 U912 ( .A1(G1991), .A2(n886), .ZN(n1003) );
  NOR2_X1 U913 ( .A1(n816), .A2(n1003), .ZN(n817) );
  NOR2_X1 U914 ( .A1(n818), .A2(n817), .ZN(n819) );
  NOR2_X1 U915 ( .A1(n1005), .A2(n819), .ZN(n820) );
  XNOR2_X1 U916 ( .A(KEYINPUT39), .B(n820), .ZN(n821) );
  NAND2_X1 U917 ( .A1(n821), .A2(n823), .ZN(n825) );
  NOR2_X1 U918 ( .A1(n822), .A2(n893), .ZN(n1012) );
  NAND2_X1 U919 ( .A1(n1012), .A2(n823), .ZN(n824) );
  AND2_X1 U920 ( .A1(n825), .A2(n824), .ZN(n826) );
  OR2_X1 U921 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U922 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U923 ( .A(n830), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n831), .ZN(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n832) );
  NAND2_X1 U926 ( .A1(G661), .A2(n832), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n833) );
  XOR2_X1 U928 ( .A(KEYINPUT111), .B(n833), .Z(n834) );
  NAND2_X1 U929 ( .A1(n835), .A2(n834), .ZN(G188) );
  INV_X1 U931 ( .A(G108), .ZN(G238) );
  INV_X1 U932 ( .A(G96), .ZN(G221) );
  NOR2_X1 U933 ( .A1(n837), .A2(n836), .ZN(G325) );
  INV_X1 U934 ( .A(G325), .ZN(G261) );
  INV_X1 U935 ( .A(n838), .ZN(G319) );
  XOR2_X1 U936 ( .A(G2100), .B(G2096), .Z(n840) );
  XNOR2_X1 U937 ( .A(KEYINPUT42), .B(G2678), .ZN(n839) );
  XNOR2_X1 U938 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U939 ( .A(KEYINPUT43), .B(G2090), .Z(n842) );
  XNOR2_X1 U940 ( .A(G2067), .B(G2072), .ZN(n841) );
  XNOR2_X1 U941 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U942 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U943 ( .A(G2078), .B(G2084), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n846), .B(n845), .ZN(G227) );
  XOR2_X1 U945 ( .A(G1986), .B(G1976), .Z(n848) );
  XNOR2_X1 U946 ( .A(G1961), .B(G1971), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U948 ( .A(n849), .B(G2474), .Z(n851) );
  XNOR2_X1 U949 ( .A(G1996), .B(G1991), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U951 ( .A(KEYINPUT41), .B(G1956), .Z(n853) );
  XNOR2_X1 U952 ( .A(G1981), .B(G1966), .ZN(n852) );
  XNOR2_X1 U953 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(G229) );
  NAND2_X1 U955 ( .A1(G124), .A2(n873), .ZN(n856) );
  XNOR2_X1 U956 ( .A(n856), .B(KEYINPUT44), .ZN(n858) );
  NAND2_X1 U957 ( .A1(n872), .A2(G112), .ZN(n857) );
  NAND2_X1 U958 ( .A1(n858), .A2(n857), .ZN(n862) );
  NAND2_X1 U959 ( .A1(n877), .A2(G100), .ZN(n860) );
  NAND2_X1 U960 ( .A1(G136), .A2(n621), .ZN(n859) );
  NAND2_X1 U961 ( .A1(n860), .A2(n859), .ZN(n861) );
  NOR2_X1 U962 ( .A1(n862), .A2(n861), .ZN(G162) );
  NAND2_X1 U963 ( .A1(n877), .A2(G103), .ZN(n864) );
  NAND2_X1 U964 ( .A1(G139), .A2(n621), .ZN(n863) );
  NAND2_X1 U965 ( .A1(n864), .A2(n863), .ZN(n869) );
  NAND2_X1 U966 ( .A1(G115), .A2(n872), .ZN(n866) );
  NAND2_X1 U967 ( .A1(G127), .A2(n873), .ZN(n865) );
  NAND2_X1 U968 ( .A1(n866), .A2(n865), .ZN(n867) );
  XOR2_X1 U969 ( .A(KEYINPUT47), .B(n867), .Z(n868) );
  NOR2_X1 U970 ( .A1(n869), .A2(n868), .ZN(n1015) );
  XOR2_X1 U971 ( .A(G162), .B(n1015), .Z(n871) );
  XNOR2_X1 U972 ( .A(G160), .B(G164), .ZN(n870) );
  XNOR2_X1 U973 ( .A(n871), .B(n870), .ZN(n884) );
  NAND2_X1 U974 ( .A1(G118), .A2(n872), .ZN(n875) );
  NAND2_X1 U975 ( .A1(G130), .A2(n873), .ZN(n874) );
  NAND2_X1 U976 ( .A1(n875), .A2(n874), .ZN(n882) );
  NAND2_X1 U977 ( .A1(G142), .A2(n621), .ZN(n876) );
  XNOR2_X1 U978 ( .A(n876), .B(KEYINPUT112), .ZN(n879) );
  NAND2_X1 U979 ( .A1(G106), .A2(n877), .ZN(n878) );
  NAND2_X1 U980 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U981 ( .A(n880), .B(KEYINPUT45), .Z(n881) );
  NOR2_X1 U982 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U983 ( .A(n884), .B(n883), .Z(n889) );
  XNOR2_X1 U984 ( .A(n999), .B(n885), .ZN(n887) );
  XNOR2_X1 U985 ( .A(n887), .B(n886), .ZN(n888) );
  XOR2_X1 U986 ( .A(n889), .B(n888), .Z(n895) );
  XOR2_X1 U987 ( .A(KEYINPUT48), .B(KEYINPUT114), .Z(n891) );
  XNOR2_X1 U988 ( .A(KEYINPUT46), .B(KEYINPUT113), .ZN(n890) );
  XNOR2_X1 U989 ( .A(n891), .B(n890), .ZN(n892) );
  XNOR2_X1 U990 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U991 ( .A(n895), .B(n894), .ZN(n896) );
  NOR2_X1 U992 ( .A1(G37), .A2(n896), .ZN(G395) );
  XNOR2_X1 U993 ( .A(n897), .B(KEYINPUT115), .ZN(n900) );
  XNOR2_X1 U994 ( .A(G171), .B(n898), .ZN(n899) );
  XNOR2_X1 U995 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U996 ( .A(n901), .B(G286), .ZN(n902) );
  NOR2_X1 U997 ( .A1(G37), .A2(n902), .ZN(G397) );
  XNOR2_X1 U998 ( .A(G2451), .B(G2446), .ZN(n912) );
  XOR2_X1 U999 ( .A(G2430), .B(KEYINPUT110), .Z(n904) );
  XNOR2_X1 U1000 ( .A(G2454), .B(G2435), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n908) );
  XOR2_X1 U1002 ( .A(G2438), .B(KEYINPUT109), .Z(n906) );
  XNOR2_X1 U1003 ( .A(G1341), .B(G1348), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1005 ( .A(n908), .B(n907), .Z(n910) );
  XNOR2_X1 U1006 ( .A(G2443), .B(G2427), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(n910), .B(n909), .ZN(n911) );
  XNOR2_X1 U1008 ( .A(n912), .B(n911), .ZN(n913) );
  NAND2_X1 U1009 ( .A1(n913), .A2(G14), .ZN(n919) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n919), .ZN(n916) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n914) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n914), .ZN(n915) );
  NOR2_X1 U1013 ( .A1(n916), .A2(n915), .ZN(n918) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1015 ( .A1(n918), .A2(n917), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(G69), .ZN(G235) );
  INV_X1 U1018 ( .A(n919), .ZN(G401) );
  XNOR2_X1 U1019 ( .A(KEYINPUT121), .B(G2067), .ZN(n920) );
  XNOR2_X1 U1020 ( .A(n920), .B(G26), .ZN(n928) );
  XNOR2_X1 U1021 ( .A(G1996), .B(G32), .ZN(n922) );
  XNOR2_X1 U1022 ( .A(G1991), .B(G25), .ZN(n921) );
  NOR2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1024 ( .A1(G28), .A2(n923), .ZN(n926) );
  XNOR2_X1 U1025 ( .A(KEYINPUT122), .B(G2072), .ZN(n924) );
  XNOR2_X1 U1026 ( .A(G33), .B(n924), .ZN(n925) );
  NOR2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n931) );
  XNOR2_X1 U1029 ( .A(G27), .B(n929), .ZN(n930) );
  NOR2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1031 ( .A(KEYINPUT53), .B(n932), .Z(n935) );
  XOR2_X1 U1032 ( .A(G34), .B(KEYINPUT54), .Z(n933) );
  XNOR2_X1 U1033 ( .A(G2084), .B(n933), .ZN(n934) );
  NAND2_X1 U1034 ( .A1(n935), .A2(n934), .ZN(n937) );
  XNOR2_X1 U1035 ( .A(G35), .B(G2090), .ZN(n936) );
  NOR2_X1 U1036 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1037 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n1023) );
  XNOR2_X1 U1038 ( .A(n938), .B(n1023), .ZN(n939) );
  NOR2_X1 U1039 ( .A1(G29), .A2(n939), .ZN(n994) );
  XNOR2_X1 U1040 ( .A(G16), .B(KEYINPUT56), .ZN(n966) );
  XOR2_X1 U1041 ( .A(G168), .B(G1966), .Z(n940) );
  NOR2_X1 U1042 ( .A1(n941), .A2(n940), .ZN(n942) );
  XOR2_X1 U1043 ( .A(KEYINPUT57), .B(n942), .Z(n964) );
  XNOR2_X1 U1044 ( .A(n943), .B(G1956), .ZN(n956) );
  XNOR2_X1 U1045 ( .A(G166), .B(G1971), .ZN(n950) );
  INV_X1 U1046 ( .A(n944), .ZN(n946) );
  NAND2_X1 U1047 ( .A1(n946), .A2(n945), .ZN(n948) );
  XNOR2_X1 U1048 ( .A(G1961), .B(G301), .ZN(n947) );
  NOR2_X1 U1049 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1050 ( .A1(n950), .A2(n949), .ZN(n954) );
  XOR2_X1 U1051 ( .A(G1348), .B(n951), .Z(n952) );
  XNOR2_X1 U1052 ( .A(KEYINPUT123), .B(n952), .ZN(n953) );
  NOR2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1054 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1056 ( .A(KEYINPUT124), .B(n959), .Z(n962) );
  XOR2_X1 U1057 ( .A(n960), .B(G1341), .Z(n961) );
  NOR2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n992) );
  INV_X1 U1061 ( .A(G16), .ZN(n990) );
  XOR2_X1 U1062 ( .A(G1961), .B(G5), .Z(n974) );
  XNOR2_X1 U1063 ( .A(G1971), .B(G22), .ZN(n968) );
  XNOR2_X1 U1064 ( .A(G23), .B(G1976), .ZN(n967) );
  NOR2_X1 U1065 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1066 ( .A(KEYINPUT126), .B(n969), .Z(n971) );
  XNOR2_X1 U1067 ( .A(G1986), .B(G24), .ZN(n970) );
  NOR2_X1 U1068 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1069 ( .A(KEYINPUT58), .B(n972), .ZN(n973) );
  NAND2_X1 U1070 ( .A1(n974), .A2(n973), .ZN(n987) );
  XOR2_X1 U1071 ( .A(G1966), .B(G21), .Z(n985) );
  XNOR2_X1 U1072 ( .A(G1348), .B(KEYINPUT59), .ZN(n975) );
  XNOR2_X1 U1073 ( .A(n975), .B(G4), .ZN(n979) );
  XNOR2_X1 U1074 ( .A(G1956), .B(G20), .ZN(n977) );
  XNOR2_X1 U1075 ( .A(G19), .B(G1341), .ZN(n976) );
  NOR2_X1 U1076 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1077 ( .A1(n979), .A2(n978), .ZN(n982) );
  XOR2_X1 U1078 ( .A(KEYINPUT125), .B(G1981), .Z(n980) );
  XNOR2_X1 U1079 ( .A(G6), .B(n980), .ZN(n981) );
  NOR2_X1 U1080 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1081 ( .A(n983), .B(KEYINPUT60), .ZN(n984) );
  NAND2_X1 U1082 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1083 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1084 ( .A(KEYINPUT61), .B(n988), .ZN(n989) );
  NAND2_X1 U1085 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1086 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1088 ( .A1(G11), .A2(n995), .ZN(n996) );
  XNOR2_X1 U1089 ( .A(n996), .B(KEYINPUT127), .ZN(n1027) );
  XOR2_X1 U1090 ( .A(G160), .B(G2084), .Z(n997) );
  XNOR2_X1 U1091 ( .A(KEYINPUT116), .B(n997), .ZN(n998) );
  NOR2_X1 U1092 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1093 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NOR2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1010) );
  XOR2_X1 U1095 ( .A(G2090), .B(G162), .Z(n1004) );
  NOR2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1097 ( .A(n1006), .B(KEYINPUT51), .ZN(n1007) );
  NOR2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1101 ( .A(KEYINPUT117), .B(n1013), .Z(n1020) );
  XOR2_X1 U1102 ( .A(G164), .B(G2078), .Z(n1014) );
  XNOR2_X1 U1103 ( .A(KEYINPUT118), .B(n1014), .ZN(n1017) );
  XOR2_X1 U1104 ( .A(G2072), .B(n1015), .Z(n1016) );
  NOR2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1106 ( .A(KEYINPUT50), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1108 ( .A(n1021), .B(KEYINPUT119), .ZN(n1022) );
  XNOR2_X1 U1109 ( .A(n1022), .B(KEYINPUT52), .ZN(n1024) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1111 ( .A1(G29), .A2(n1025), .ZN(n1026) );
  NAND2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XOR2_X1 U1113 ( .A(KEYINPUT62), .B(n1028), .Z(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

