

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587;

  XNOR2_X1 U327 ( .A(n452), .B(n451), .ZN(n527) );
  NOR2_X1 U328 ( .A1(n453), .A2(n527), .ZN(n563) );
  XOR2_X1 U329 ( .A(n554), .B(KEYINPUT82), .Z(n537) );
  XNOR2_X1 U330 ( .A(KEYINPUT48), .B(KEYINPUT116), .ZN(n378) );
  XNOR2_X1 U331 ( .A(n379), .B(n378), .ZN(n526) );
  XNOR2_X1 U332 ( .A(n413), .B(KEYINPUT64), .ZN(n570) );
  INV_X1 U333 ( .A(G190GAT), .ZN(n454) );
  XOR2_X1 U334 ( .A(KEYINPUT95), .B(n466), .Z(n541) );
  XNOR2_X1 U335 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U336 ( .A(n457), .B(n456), .ZN(G1351GAT) );
  XOR2_X1 U337 ( .A(KEYINPUT65), .B(KEYINPUT11), .Z(n296) );
  XNOR2_X1 U338 ( .A(KEYINPUT67), .B(KEYINPUT78), .ZN(n295) );
  XNOR2_X1 U339 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U340 ( .A(KEYINPUT80), .B(KEYINPUT9), .Z(n298) );
  XNOR2_X1 U341 ( .A(KEYINPUT81), .B(KEYINPUT10), .ZN(n297) );
  XNOR2_X1 U342 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U343 ( .A(n300), .B(n299), .Z(n305) );
  XNOR2_X1 U344 ( .A(G50GAT), .B(KEYINPUT77), .ZN(n301) );
  XNOR2_X1 U345 ( .A(n301), .B(G162GAT), .ZN(n414) );
  XOR2_X1 U346 ( .A(G92GAT), .B(G218GAT), .Z(n303) );
  XNOR2_X1 U347 ( .A(G36GAT), .B(G190GAT), .ZN(n302) );
  XNOR2_X1 U348 ( .A(n303), .B(n302), .ZN(n387) );
  XNOR2_X1 U349 ( .A(n414), .B(n387), .ZN(n304) );
  XNOR2_X1 U350 ( .A(n305), .B(n304), .ZN(n310) );
  XNOR2_X1 U351 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n306) );
  XNOR2_X1 U352 ( .A(n306), .B(KEYINPUT7), .ZN(n344) );
  XOR2_X1 U353 ( .A(KEYINPUT79), .B(n344), .Z(n308) );
  NAND2_X1 U354 ( .A1(G232GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U355 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U356 ( .A(n310), .B(n309), .Z(n314) );
  XNOR2_X1 U357 ( .A(G29GAT), .B(G134GAT), .ZN(n311) );
  XNOR2_X1 U358 ( .A(n311), .B(G85GAT), .ZN(n409) );
  XNOR2_X1 U359 ( .A(G99GAT), .B(G106GAT), .ZN(n312) );
  XNOR2_X1 U360 ( .A(n312), .B(KEYINPUT75), .ZN(n323) );
  XNOR2_X1 U361 ( .A(n409), .B(n323), .ZN(n313) );
  XNOR2_X1 U362 ( .A(n314), .B(n313), .ZN(n554) );
  XOR2_X1 U363 ( .A(KEYINPUT33), .B(G92GAT), .Z(n316) );
  XNOR2_X1 U364 ( .A(G78GAT), .B(G85GAT), .ZN(n315) );
  XNOR2_X1 U365 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U366 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n318) );
  XNOR2_X1 U367 ( .A(KEYINPUT74), .B(KEYINPUT76), .ZN(n317) );
  XNOR2_X1 U368 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U369 ( .A(n320), .B(n319), .ZN(n330) );
  XOR2_X1 U370 ( .A(G176GAT), .B(G204GAT), .Z(n383) );
  XOR2_X1 U371 ( .A(G71GAT), .B(KEYINPUT13), .Z(n367) );
  INV_X1 U372 ( .A(n367), .ZN(n321) );
  XNOR2_X1 U373 ( .A(n383), .B(n321), .ZN(n328) );
  XNOR2_X1 U374 ( .A(G120GAT), .B(G148GAT), .ZN(n322) );
  XNOR2_X1 U375 ( .A(n322), .B(G57GAT), .ZN(n397) );
  XOR2_X1 U376 ( .A(n323), .B(G64GAT), .Z(n325) );
  NAND2_X1 U377 ( .A1(G230GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U378 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U379 ( .A(n397), .B(n326), .ZN(n327) );
  XNOR2_X1 U380 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U381 ( .A(n330), .B(n329), .ZN(n575) );
  XNOR2_X1 U382 ( .A(KEYINPUT41), .B(n575), .ZN(n562) );
  XOR2_X1 U383 ( .A(G197GAT), .B(G113GAT), .Z(n332) );
  XNOR2_X1 U384 ( .A(G169GAT), .B(G50GAT), .ZN(n331) );
  XNOR2_X1 U385 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U386 ( .A(KEYINPUT72), .B(KEYINPUT73), .Z(n334) );
  XNOR2_X1 U387 ( .A(G22GAT), .B(G141GAT), .ZN(n333) );
  XNOR2_X1 U388 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U389 ( .A(n336), .B(n335), .Z(n341) );
  XOR2_X1 U390 ( .A(KEYINPUT30), .B(G8GAT), .Z(n338) );
  NAND2_X1 U391 ( .A1(G229GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U392 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U393 ( .A(KEYINPUT29), .B(n339), .ZN(n340) );
  XNOR2_X1 U394 ( .A(n341), .B(n340), .ZN(n350) );
  XOR2_X1 U395 ( .A(KEYINPUT68), .B(G1GAT), .Z(n343) );
  XNOR2_X1 U396 ( .A(KEYINPUT69), .B(KEYINPUT71), .ZN(n342) );
  XNOR2_X1 U397 ( .A(n343), .B(n342), .ZN(n348) );
  XOR2_X1 U398 ( .A(G15GAT), .B(KEYINPUT70), .Z(n366) );
  XOR2_X1 U399 ( .A(n366), .B(G36GAT), .Z(n346) );
  XNOR2_X1 U400 ( .A(n344), .B(G29GAT), .ZN(n345) );
  XNOR2_X1 U401 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U402 ( .A(n348), .B(n347), .Z(n349) );
  XOR2_X1 U403 ( .A(n350), .B(n349), .Z(n544) );
  INV_X1 U404 ( .A(n544), .ZN(n571) );
  NAND2_X1 U405 ( .A1(n562), .A2(n571), .ZN(n352) );
  XNOR2_X1 U406 ( .A(KEYINPUT46), .B(KEYINPUT114), .ZN(n351) );
  XNOR2_X1 U407 ( .A(n352), .B(n351), .ZN(n369) );
  XOR2_X1 U408 ( .A(KEYINPUT12), .B(KEYINPUT83), .Z(n354) );
  NAND2_X1 U409 ( .A1(G231GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U410 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U411 ( .A(n355), .B(KEYINPUT15), .Z(n360) );
  XNOR2_X1 U412 ( .A(G22GAT), .B(G155GAT), .ZN(n356) );
  XNOR2_X1 U413 ( .A(n356), .B(G78GAT), .ZN(n428) );
  XOR2_X1 U414 ( .A(G64GAT), .B(G211GAT), .Z(n358) );
  XNOR2_X1 U415 ( .A(G8GAT), .B(G183GAT), .ZN(n357) );
  XNOR2_X1 U416 ( .A(n358), .B(n357), .ZN(n380) );
  XNOR2_X1 U417 ( .A(n428), .B(n380), .ZN(n359) );
  XNOR2_X1 U418 ( .A(n360), .B(n359), .ZN(n362) );
  INV_X1 U419 ( .A(KEYINPUT14), .ZN(n361) );
  XNOR2_X1 U420 ( .A(n362), .B(n361), .ZN(n364) );
  XOR2_X1 U421 ( .A(G1GAT), .B(G127GAT), .Z(n402) );
  XNOR2_X1 U422 ( .A(G57GAT), .B(n402), .ZN(n363) );
  XNOR2_X1 U423 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U424 ( .A(n366), .B(n365), .ZN(n368) );
  XNOR2_X1 U425 ( .A(n368), .B(n367), .ZN(n550) );
  XOR2_X1 U426 ( .A(KEYINPUT113), .B(n550), .Z(n567) );
  NAND2_X1 U427 ( .A1(n369), .A2(n567), .ZN(n370) );
  NOR2_X1 U428 ( .A1(n554), .A2(n370), .ZN(n372) );
  XNOR2_X1 U429 ( .A(KEYINPUT47), .B(KEYINPUT115), .ZN(n371) );
  XNOR2_X1 U430 ( .A(n372), .B(n371), .ZN(n377) );
  XNOR2_X1 U431 ( .A(KEYINPUT36), .B(n537), .ZN(n585) );
  NOR2_X1 U432 ( .A1(n550), .A2(n585), .ZN(n373) );
  XNOR2_X1 U433 ( .A(n373), .B(KEYINPUT45), .ZN(n374) );
  NAND2_X1 U434 ( .A1(n374), .A2(n575), .ZN(n375) );
  NOR2_X1 U435 ( .A1(n571), .A2(n375), .ZN(n376) );
  NOR2_X1 U436 ( .A1(n377), .A2(n376), .ZN(n379) );
  XOR2_X1 U437 ( .A(G197GAT), .B(KEYINPUT21), .Z(n420) );
  XOR2_X1 U438 ( .A(n380), .B(n420), .Z(n382) );
  NAND2_X1 U439 ( .A1(G226GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U440 ( .A(n382), .B(n381), .ZN(n384) );
  XOR2_X1 U441 ( .A(n384), .B(n383), .Z(n389) );
  XOR2_X1 U442 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n386) );
  XNOR2_X1 U443 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n385) );
  XNOR2_X1 U444 ( .A(n386), .B(n385), .ZN(n437) );
  XNOR2_X1 U445 ( .A(n437), .B(n387), .ZN(n388) );
  XNOR2_X1 U446 ( .A(n389), .B(n388), .ZN(n517) );
  XNOR2_X1 U447 ( .A(n517), .B(KEYINPUT120), .ZN(n390) );
  NOR2_X1 U448 ( .A1(n526), .A2(n390), .ZN(n391) );
  XNOR2_X1 U449 ( .A(n391), .B(KEYINPUT54), .ZN(n412) );
  XOR2_X1 U450 ( .A(KEYINPUT1), .B(KEYINPUT5), .Z(n393) );
  NAND2_X1 U451 ( .A1(G225GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U452 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U453 ( .A(n394), .B(KEYINPUT4), .Z(n399) );
  XOR2_X1 U454 ( .A(KEYINPUT89), .B(KEYINPUT3), .Z(n396) );
  XNOR2_X1 U455 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n395) );
  XNOR2_X1 U456 ( .A(n396), .B(n395), .ZN(n427) );
  XNOR2_X1 U457 ( .A(n427), .B(n397), .ZN(n398) );
  XNOR2_X1 U458 ( .A(n399), .B(n398), .ZN(n407) );
  XOR2_X1 U459 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n401) );
  XNOR2_X1 U460 ( .A(KEYINPUT6), .B(KEYINPUT94), .ZN(n400) );
  XNOR2_X1 U461 ( .A(n401), .B(n400), .ZN(n403) );
  XOR2_X1 U462 ( .A(n403), .B(n402), .Z(n405) );
  XNOR2_X1 U463 ( .A(G155GAT), .B(G162GAT), .ZN(n404) );
  XNOR2_X1 U464 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U465 ( .A(n407), .B(n406), .Z(n411) );
  XNOR2_X1 U466 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n408) );
  XNOR2_X1 U467 ( .A(n408), .B(KEYINPUT84), .ZN(n436) );
  XNOR2_X1 U468 ( .A(n436), .B(n409), .ZN(n410) );
  XNOR2_X1 U469 ( .A(n411), .B(n410), .ZN(n466) );
  NAND2_X1 U470 ( .A1(n412), .A2(n541), .ZN(n413) );
  XOR2_X1 U471 ( .A(n414), .B(KEYINPUT91), .Z(n416) );
  NAND2_X1 U472 ( .A1(G228GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U473 ( .A(n416), .B(n415), .ZN(n432) );
  XOR2_X1 U474 ( .A(KEYINPUT24), .B(G211GAT), .Z(n418) );
  XNOR2_X1 U475 ( .A(KEYINPUT23), .B(KEYINPUT90), .ZN(n417) );
  XNOR2_X1 U476 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U477 ( .A(n419), .B(G106GAT), .Z(n422) );
  XNOR2_X1 U478 ( .A(n420), .B(G218GAT), .ZN(n421) );
  XNOR2_X1 U479 ( .A(n422), .B(n421), .ZN(n426) );
  XOR2_X1 U480 ( .A(G204GAT), .B(G148GAT), .Z(n424) );
  XNOR2_X1 U481 ( .A(KEYINPUT22), .B(KEYINPUT88), .ZN(n423) );
  XNOR2_X1 U482 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U483 ( .A(n426), .B(n425), .Z(n430) );
  XNOR2_X1 U484 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U485 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U486 ( .A(n432), .B(n431), .ZN(n469) );
  NOR2_X1 U487 ( .A1(n570), .A2(n469), .ZN(n433) );
  XNOR2_X1 U488 ( .A(n433), .B(KEYINPUT55), .ZN(n453) );
  XOR2_X1 U489 ( .A(G176GAT), .B(KEYINPUT85), .Z(n435) );
  XNOR2_X1 U490 ( .A(KEYINPUT86), .B(KEYINPUT87), .ZN(n434) );
  XNOR2_X1 U491 ( .A(n435), .B(n434), .ZN(n452) );
  XNOR2_X1 U492 ( .A(n437), .B(n436), .ZN(n450) );
  XOR2_X1 U493 ( .A(G190GAT), .B(G134GAT), .Z(n439) );
  XNOR2_X1 U494 ( .A(G43GAT), .B(G99GAT), .ZN(n438) );
  XNOR2_X1 U495 ( .A(n439), .B(n438), .ZN(n443) );
  XOR2_X1 U496 ( .A(KEYINPUT20), .B(G71GAT), .Z(n441) );
  XNOR2_X1 U497 ( .A(G15GAT), .B(G183GAT), .ZN(n440) );
  XNOR2_X1 U498 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U499 ( .A(n443), .B(n442), .Z(n448) );
  XOR2_X1 U500 ( .A(G127GAT), .B(G120GAT), .Z(n445) );
  NAND2_X1 U501 ( .A1(G227GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U502 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U503 ( .A(KEYINPUT66), .B(n446), .ZN(n447) );
  XNOR2_X1 U504 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U505 ( .A(n450), .B(n449), .ZN(n451) );
  INV_X1 U506 ( .A(n563), .ZN(n566) );
  NOR2_X1 U507 ( .A1(n537), .A2(n566), .ZN(n457) );
  XNOR2_X1 U508 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n455) );
  NAND2_X1 U509 ( .A1(n575), .A2(n571), .ZN(n491) );
  XOR2_X1 U510 ( .A(KEYINPUT26), .B(KEYINPUT97), .Z(n459) );
  NAND2_X1 U511 ( .A1(n469), .A2(n527), .ZN(n458) );
  XNOR2_X1 U512 ( .A(n459), .B(n458), .ZN(n569) );
  XOR2_X1 U513 ( .A(n517), .B(KEYINPUT27), .Z(n470) );
  INV_X1 U514 ( .A(n470), .ZN(n460) );
  NOR2_X1 U515 ( .A1(n569), .A2(n460), .ZN(n543) );
  NOR2_X1 U516 ( .A1(n517), .A2(n527), .ZN(n461) );
  XNOR2_X1 U517 ( .A(n461), .B(KEYINPUT98), .ZN(n462) );
  NOR2_X1 U518 ( .A1(n469), .A2(n462), .ZN(n463) );
  XOR2_X1 U519 ( .A(KEYINPUT25), .B(n463), .Z(n464) );
  NOR2_X1 U520 ( .A1(n543), .A2(n464), .ZN(n465) );
  XNOR2_X1 U521 ( .A(KEYINPUT99), .B(n465), .ZN(n467) );
  NAND2_X1 U522 ( .A1(n467), .A2(n466), .ZN(n468) );
  XNOR2_X1 U523 ( .A(n468), .B(KEYINPUT100), .ZN(n474) );
  XOR2_X1 U524 ( .A(KEYINPUT28), .B(n469), .Z(n522) );
  NAND2_X1 U525 ( .A1(n470), .A2(n522), .ZN(n471) );
  NOR2_X1 U526 ( .A1(n541), .A2(n471), .ZN(n529) );
  XNOR2_X1 U527 ( .A(KEYINPUT96), .B(n529), .ZN(n472) );
  NAND2_X1 U528 ( .A1(n472), .A2(n527), .ZN(n473) );
  NAND2_X1 U529 ( .A1(n474), .A2(n473), .ZN(n488) );
  INV_X1 U530 ( .A(n550), .ZN(n580) );
  NAND2_X1 U531 ( .A1(n537), .A2(n580), .ZN(n475) );
  XOR2_X1 U532 ( .A(KEYINPUT16), .B(n475), .Z(n476) );
  NAND2_X1 U533 ( .A1(n488), .A2(n476), .ZN(n477) );
  XOR2_X1 U534 ( .A(KEYINPUT101), .B(n477), .Z(n503) );
  OR2_X1 U535 ( .A1(n491), .A2(n503), .ZN(n486) );
  NOR2_X1 U536 ( .A1(n541), .A2(n486), .ZN(n479) );
  XNOR2_X1 U537 ( .A(KEYINPUT102), .B(KEYINPUT34), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n479), .B(n478), .ZN(n480) );
  XOR2_X1 U539 ( .A(G1GAT), .B(n480), .Z(G1324GAT) );
  NOR2_X1 U540 ( .A1(n517), .A2(n486), .ZN(n482) );
  XNOR2_X1 U541 ( .A(G8GAT), .B(KEYINPUT103), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n482), .B(n481), .ZN(G1325GAT) );
  NOR2_X1 U543 ( .A1(n527), .A2(n486), .ZN(n484) );
  XNOR2_X1 U544 ( .A(KEYINPUT35), .B(KEYINPUT104), .ZN(n483) );
  XNOR2_X1 U545 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U546 ( .A(G15GAT), .B(n485), .ZN(G1326GAT) );
  NOR2_X1 U547 ( .A1(n522), .A2(n486), .ZN(n487) );
  XOR2_X1 U548 ( .A(G22GAT), .B(n487), .Z(G1327GAT) );
  XNOR2_X1 U549 ( .A(KEYINPUT105), .B(KEYINPUT39), .ZN(n494) );
  NAND2_X1 U550 ( .A1(n550), .A2(n488), .ZN(n489) );
  NOR2_X1 U551 ( .A1(n585), .A2(n489), .ZN(n490) );
  XNOR2_X1 U552 ( .A(KEYINPUT37), .B(n490), .ZN(n515) );
  NOR2_X1 U553 ( .A1(n515), .A2(n491), .ZN(n492) );
  XOR2_X1 U554 ( .A(KEYINPUT38), .B(n492), .Z(n500) );
  NOR2_X1 U555 ( .A1(n541), .A2(n500), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U557 ( .A(G29GAT), .B(n495), .Z(G1328GAT) );
  NOR2_X1 U558 ( .A1(n517), .A2(n500), .ZN(n496) );
  XOR2_X1 U559 ( .A(KEYINPUT106), .B(n496), .Z(n497) );
  XNOR2_X1 U560 ( .A(G36GAT), .B(n497), .ZN(G1329GAT) );
  NOR2_X1 U561 ( .A1(n500), .A2(n527), .ZN(n498) );
  XOR2_X1 U562 ( .A(KEYINPUT40), .B(n498), .Z(n499) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(n499), .ZN(G1330GAT) );
  NOR2_X1 U564 ( .A1(n500), .A2(n522), .ZN(n501) );
  XOR2_X1 U565 ( .A(G50GAT), .B(n501), .Z(G1331GAT) );
  NAND2_X1 U566 ( .A1(n562), .A2(n544), .ZN(n502) );
  XOR2_X1 U567 ( .A(KEYINPUT107), .B(n502), .Z(n514) );
  OR2_X1 U568 ( .A1(n503), .A2(n514), .ZN(n510) );
  NOR2_X1 U569 ( .A1(n541), .A2(n510), .ZN(n505) );
  XNOR2_X1 U570 ( .A(KEYINPUT108), .B(KEYINPUT42), .ZN(n504) );
  XNOR2_X1 U571 ( .A(n505), .B(n504), .ZN(n506) );
  XOR2_X1 U572 ( .A(G57GAT), .B(n506), .Z(G1332GAT) );
  NOR2_X1 U573 ( .A1(n517), .A2(n510), .ZN(n507) );
  XOR2_X1 U574 ( .A(G64GAT), .B(n507), .Z(G1333GAT) );
  NOR2_X1 U575 ( .A1(n527), .A2(n510), .ZN(n509) );
  XNOR2_X1 U576 ( .A(G71GAT), .B(KEYINPUT109), .ZN(n508) );
  XNOR2_X1 U577 ( .A(n509), .B(n508), .ZN(G1334GAT) );
  NOR2_X1 U578 ( .A1(n522), .A2(n510), .ZN(n512) );
  XNOR2_X1 U579 ( .A(KEYINPUT110), .B(KEYINPUT43), .ZN(n511) );
  XNOR2_X1 U580 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U581 ( .A(G78GAT), .B(n513), .ZN(G1335GAT) );
  OR2_X1 U582 ( .A1(n515), .A2(n514), .ZN(n521) );
  NOR2_X1 U583 ( .A1(n541), .A2(n521), .ZN(n516) );
  XOR2_X1 U584 ( .A(G85GAT), .B(n516), .Z(G1336GAT) );
  NOR2_X1 U585 ( .A1(n517), .A2(n521), .ZN(n518) );
  XOR2_X1 U586 ( .A(G92GAT), .B(n518), .Z(G1337GAT) );
  NOR2_X1 U587 ( .A1(n527), .A2(n521), .ZN(n520) );
  XNOR2_X1 U588 ( .A(G99GAT), .B(KEYINPUT111), .ZN(n519) );
  XNOR2_X1 U589 ( .A(n520), .B(n519), .ZN(G1338GAT) );
  NOR2_X1 U590 ( .A1(n522), .A2(n521), .ZN(n524) );
  XNOR2_X1 U591 ( .A(KEYINPUT112), .B(KEYINPUT44), .ZN(n523) );
  XNOR2_X1 U592 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U593 ( .A(G106GAT), .B(n525), .Z(G1339GAT) );
  NOR2_X1 U594 ( .A1(n526), .A2(n527), .ZN(n528) );
  NAND2_X1 U595 ( .A1(n529), .A2(n528), .ZN(n536) );
  NOR2_X1 U596 ( .A1(n544), .A2(n536), .ZN(n530) );
  XOR2_X1 U597 ( .A(G113GAT), .B(n530), .Z(G1340GAT) );
  INV_X1 U598 ( .A(n562), .ZN(n546) );
  NOR2_X1 U599 ( .A1(n546), .A2(n536), .ZN(n532) );
  XNOR2_X1 U600 ( .A(KEYINPUT49), .B(KEYINPUT117), .ZN(n531) );
  XNOR2_X1 U601 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U602 ( .A(G120GAT), .B(n533), .Z(G1341GAT) );
  NOR2_X1 U603 ( .A1(n567), .A2(n536), .ZN(n534) );
  XOR2_X1 U604 ( .A(KEYINPUT50), .B(n534), .Z(n535) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  NOR2_X1 U606 ( .A1(n537), .A2(n536), .ZN(n539) );
  XNOR2_X1 U607 ( .A(KEYINPUT51), .B(KEYINPUT118), .ZN(n538) );
  XNOR2_X1 U608 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U609 ( .A(G134GAT), .B(n540), .ZN(G1343GAT) );
  NOR2_X1 U610 ( .A1(n541), .A2(n526), .ZN(n542) );
  NAND2_X1 U611 ( .A1(n543), .A2(n542), .ZN(n553) );
  NOR2_X1 U612 ( .A1(n544), .A2(n553), .ZN(n545) );
  XOR2_X1 U613 ( .A(G141GAT), .B(n545), .Z(G1344GAT) );
  NOR2_X1 U614 ( .A1(n546), .A2(n553), .ZN(n548) );
  XNOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n547) );
  XNOR2_X1 U616 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(n549), .ZN(G1345GAT) );
  NOR2_X1 U618 ( .A1(n550), .A2(n553), .ZN(n552) );
  XNOR2_X1 U619 ( .A(G155GAT), .B(KEYINPUT119), .ZN(n551) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(G1346GAT) );
  INV_X1 U621 ( .A(n553), .ZN(n555) );
  NAND2_X1 U622 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U624 ( .A(G169GAT), .B(KEYINPUT121), .Z(n558) );
  NAND2_X1 U625 ( .A1(n563), .A2(n571), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n558), .B(n557), .ZN(G1348GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n560) );
  XNOR2_X1 U628 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n559) );
  XNOR2_X1 U629 ( .A(n560), .B(n559), .ZN(n561) );
  XOR2_X1 U630 ( .A(KEYINPUT56), .B(n561), .Z(n565) );
  NAND2_X1 U631 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(G1349GAT) );
  NOR2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U634 ( .A(G183GAT), .B(n568), .Z(G1350GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n573) );
  NOR2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n579) );
  NAND2_X1 U637 ( .A1(n579), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(n574), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n577) );
  INV_X1 U641 ( .A(n579), .ZN(n584) );
  OR2_X1 U642 ( .A1(n584), .A2(n575), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n578) );
  XOR2_X1 U644 ( .A(G204GAT), .B(n578), .Z(G1353GAT) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n583) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(n587) );
  NOR2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U651 ( .A(n587), .B(n586), .Z(G1355GAT) );
endmodule

