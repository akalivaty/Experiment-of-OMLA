//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 0 1 1 1 0 1 0 0 0 0 0 1 0 0 0 1 1 0 1 1 1 0 1 0 1 0 0 1 1 0 0 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(new_n206), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n222));
  INV_X1    g0022(.A(G77), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  INV_X1    g0024(.A(G107), .ZN(new_n225));
  INV_X1    g0025(.A(G264), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n208), .B1(new_n221), .B2(new_n227), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n211), .B1(new_n214), .B2(new_n215), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G87), .B(G97), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT64), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  NOR3_X1   g0046(.A1(new_n206), .A2(KEYINPUT23), .A3(G107), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT83), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT67), .B(G107), .ZN(new_n249));
  OAI21_X1  g0049(.A(KEYINPUT23), .B1(new_n249), .B2(new_n206), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT22), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT3), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n206), .A2(G87), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n251), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AND3_X1   g0058(.A1(new_n248), .A2(new_n250), .A3(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(KEYINPUT72), .B1(new_n252), .B2(KEYINPUT3), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT72), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(new_n254), .A3(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT71), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n264), .B1(new_n254), .B2(G33), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n252), .A2(KEYINPUT71), .A3(KEYINPUT3), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n251), .A2(new_n219), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n263), .A2(new_n265), .A3(new_n266), .A4(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G116), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n206), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n259), .A2(new_n271), .A3(KEYINPUT24), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT24), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n248), .A2(new_n250), .A3(new_n258), .ZN(new_n274));
  AOI21_X1  g0074(.A(G20), .B1(new_n268), .B2(new_n269), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n212), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n272), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n280));
  OAI21_X1  g0080(.A(KEYINPUT25), .B1(new_n280), .B2(G107), .ZN(new_n281));
  OR3_X1    g0081(.A1(new_n280), .A2(KEYINPUT25), .A3(G107), .ZN(new_n282));
  INV_X1    g0082(.A(new_n278), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n283), .B(new_n280), .C1(G1), .C2(new_n252), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n281), .B(new_n282), .C1(new_n284), .C2(new_n225), .ZN(new_n285));
  XNOR2_X1  g0085(.A(new_n285), .B(KEYINPUT84), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n279), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(KEYINPUT85), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT85), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n279), .A2(new_n289), .A3(new_n286), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n265), .A2(new_n266), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G250), .A2(G1698), .ZN(new_n292));
  INV_X1    g0092(.A(G257), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n292), .B1(new_n293), .B2(G1698), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n291), .A2(new_n263), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(G33), .A2(G294), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT86), .ZN(new_n300));
  INV_X1    g0100(.A(G274), .ZN(new_n301));
  INV_X1    g0101(.A(new_n212), .ZN(new_n302));
  NAND2_X1  g0102(.A1(G33), .A2(G41), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G45), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n305), .A2(G1), .ZN(new_n306));
  XNOR2_X1  g0106(.A(KEYINPUT5), .B(G41), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n304), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  AND2_X1   g0108(.A1(KEYINPUT5), .A2(G41), .ZN(new_n309));
  NOR2_X1   g0109(.A1(KEYINPUT5), .A2(G41), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n306), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n303), .A2(G1), .A3(G13), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n311), .A2(G264), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n308), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n299), .A2(new_n300), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n312), .B1(new_n295), .B2(new_n296), .ZN(new_n317));
  OAI21_X1  g0117(.A(KEYINPUT86), .B1(new_n317), .B2(new_n314), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n316), .A2(G169), .A3(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n317), .A2(new_n314), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G179), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n319), .A2(KEYINPUT87), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(KEYINPUT87), .B1(new_n319), .B2(new_n321), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n288), .B(new_n290), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT88), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n319), .A2(new_n321), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT87), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n319), .A2(KEYINPUT87), .A3(new_n321), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AND3_X1   g0131(.A1(new_n279), .A2(new_n289), .A3(new_n286), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n289), .B1(new_n279), .B2(new_n286), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n331), .A2(new_n334), .A3(KEYINPUT88), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n316), .A2(new_n318), .ZN(new_n336));
  OAI22_X1  g0136(.A1(new_n336), .A2(G190), .B1(G200), .B2(new_n320), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n337), .A2(new_n286), .A3(new_n279), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n326), .A2(new_n335), .A3(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(G257), .A2(G1698), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n340), .B1(new_n226), .B2(G1698), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n263), .A2(new_n341), .A3(new_n265), .A4(new_n266), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n256), .A2(G303), .ZN(new_n343));
  AND3_X1   g0143(.A1(new_n342), .A2(KEYINPUT81), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(KEYINPUT81), .B1(new_n342), .B2(new_n343), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n298), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n311), .A2(G270), .A3(new_n312), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n308), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n280), .A2(G116), .ZN(new_n349));
  INV_X1    g0149(.A(new_n280), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n252), .A2(G1), .ZN(new_n351));
  NOR3_X1   g0151(.A1(new_n350), .A2(new_n278), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n349), .B1(new_n352), .B2(G116), .ZN(new_n353));
  AOI21_X1  g0153(.A(G20), .B1(new_n252), .B2(G97), .ZN(new_n354));
  NAND2_X1  g0154(.A1(G33), .A2(G283), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT77), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(KEYINPUT77), .B1(G33), .B2(G283), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n354), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G116), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n277), .A2(new_n212), .B1(G20), .B2(new_n360), .ZN(new_n361));
  AND3_X1   g0161(.A1(new_n359), .A2(KEYINPUT20), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(KEYINPUT20), .B1(new_n359), .B2(new_n361), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n353), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n346), .A2(G179), .A3(new_n348), .A4(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(G169), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n366), .B1(new_n348), .B2(new_n346), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n365), .B1(new_n367), .B2(KEYINPUT21), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n346), .A2(new_n348), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n369), .A2(KEYINPUT21), .A3(G169), .A4(new_n364), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT82), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT82), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n367), .A2(new_n372), .A3(KEYINPUT21), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n368), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n364), .B1(new_n369), .B2(G200), .ZN(new_n375));
  INV_X1    g0175(.A(G190), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n375), .B1(new_n376), .B2(new_n369), .ZN(new_n377));
  AND2_X1   g0177(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n280), .A2(G97), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n379), .B1(new_n352), .B2(G97), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT6), .ZN(new_n381));
  INV_X1    g0181(.A(G97), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n382), .A2(new_n225), .ZN(new_n383));
  NOR2_X1   g0183(.A1(G97), .A2(G107), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n381), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n225), .A2(KEYINPUT6), .A3(G97), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(G20), .A2(G33), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n387), .A2(G20), .B1(G77), .B2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT7), .B1(new_n256), .B2(new_n206), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT7), .ZN(new_n391));
  AOI211_X1 g0191(.A(new_n391), .B(G20), .C1(new_n253), .C2(new_n255), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n249), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  AND2_X1   g0193(.A1(new_n389), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n380), .B1(new_n394), .B2(new_n283), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n311), .A2(new_n312), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n308), .B1(new_n396), .B2(new_n293), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  XNOR2_X1  g0198(.A(new_n355), .B(new_n356), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT4), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n400), .A2(new_n224), .ZN(new_n401));
  INV_X1    g0201(.A(G1698), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n401), .A2(new_n402), .A3(new_n253), .A4(new_n255), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n253), .A2(new_n255), .A3(G250), .A4(G1698), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n399), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n291), .A2(G244), .A3(new_n402), .A4(new_n263), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n405), .B1(new_n406), .B2(new_n400), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n398), .B1(new_n407), .B2(new_n312), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n395), .B1(G190), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT78), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  OAI211_X1 g0212(.A(KEYINPUT78), .B(new_n398), .C1(new_n407), .C2(new_n312), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(G200), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n304), .A2(new_n306), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n306), .A2(new_n220), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n312), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT79), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n263), .A2(new_n265), .A3(new_n266), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n218), .A2(G1698), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n421), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n291), .A2(G244), .A3(G1698), .A4(new_n263), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n291), .A2(KEYINPUT79), .A3(new_n263), .A4(new_n423), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n425), .A2(new_n269), .A3(new_n426), .A4(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n420), .B1(new_n428), .B2(new_n298), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(G190), .ZN(new_n430));
  XOR2_X1   g0230(.A(KEYINPUT15), .B(G87), .Z(new_n431));
  NOR2_X1   g0231(.A1(new_n431), .A2(new_n280), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n284), .A2(new_n219), .ZN(new_n433));
  NAND2_X1  g0233(.A1(G33), .A2(G97), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT19), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n206), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT80), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI211_X1 g0238(.A(KEYINPUT80), .B(new_n206), .C1(new_n434), .C2(new_n435), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n219), .A2(new_n382), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n438), .B(new_n439), .C1(new_n440), .C2(new_n249), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n252), .A2(G20), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n435), .B1(new_n443), .B2(new_n382), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n206), .A2(G68), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n441), .B(new_n444), .C1(new_n422), .C2(new_n445), .ZN(new_n446));
  AOI211_X1 g0246(.A(new_n432), .B(new_n433), .C1(new_n446), .C2(new_n278), .ZN(new_n447));
  INV_X1    g0247(.A(G200), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n430), .B(new_n447), .C1(new_n448), .C2(new_n429), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n428), .A2(new_n298), .ZN(new_n450));
  INV_X1    g0250(.A(G179), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n450), .A2(new_n451), .A3(new_n419), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n432), .B1(new_n446), .B2(new_n278), .ZN(new_n453));
  INV_X1    g0253(.A(new_n431), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n453), .B1(new_n454), .B2(new_n284), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n452), .B(new_n455), .C1(G169), .C2(new_n429), .ZN(new_n456));
  INV_X1    g0256(.A(G169), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n408), .A2(new_n457), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n451), .B(new_n398), .C1(new_n407), .C2(new_n312), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n395), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  AND4_X1   g0260(.A1(new_n415), .A2(new_n449), .A3(new_n456), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n378), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n256), .ZN(new_n463));
  NOR2_X1   g0263(.A1(G222), .A2(G1698), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n402), .A2(G223), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n312), .B1(new_n256), .B2(new_n223), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n298), .A2(new_n469), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n466), .A2(new_n467), .B1(G226), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n469), .A2(new_n312), .A3(G274), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT65), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n304), .A2(KEYINPUT65), .A3(new_n469), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n471), .A2(G190), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n448), .B1(new_n471), .B2(new_n476), .ZN(new_n478));
  NOR3_X1   g0278(.A1(new_n477), .A2(new_n478), .A3(KEYINPUT10), .ZN(new_n479));
  XNOR2_X1  g0279(.A(KEYINPUT8), .B(G58), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(KEYINPUT66), .ZN(new_n481));
  INV_X1    g0281(.A(G58), .ZN(new_n482));
  NOR3_X1   g0282(.A1(new_n482), .A2(KEYINPUT66), .A3(KEYINPUT8), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n481), .A2(new_n484), .A3(new_n442), .ZN(new_n485));
  INV_X1    g0285(.A(G150), .ZN(new_n486));
  INV_X1    g0286(.A(new_n388), .ZN(new_n487));
  OAI22_X1  g0287(.A1(new_n486), .A2(new_n487), .B1(new_n201), .B2(new_n206), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n283), .B1(new_n485), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n350), .A2(new_n278), .ZN(new_n491));
  INV_X1    g0291(.A(G50), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n492), .B1(new_n205), .B2(G20), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n491), .A2(new_n493), .B1(new_n492), .B2(new_n350), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(KEYINPUT9), .B1(new_n490), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT68), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT9), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n483), .B1(new_n480), .B2(KEYINPUT66), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n488), .B1(new_n499), .B2(new_n442), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n498), .B(new_n494), .C1(new_n500), .C2(new_n283), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n496), .A2(new_n497), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n497), .B1(new_n496), .B2(new_n501), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n479), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT69), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT69), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n479), .B(new_n506), .C1(new_n502), .C2(new_n503), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  OR2_X1    g0308(.A1(new_n477), .A2(new_n478), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n496), .A2(new_n501), .ZN(new_n510));
  OAI21_X1  g0310(.A(KEYINPUT10), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n490), .A2(new_n495), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n471), .A2(new_n476), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n513), .B1(new_n457), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n471), .A2(new_n451), .A3(new_n476), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n512), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n350), .A2(new_n217), .ZN(new_n520));
  XNOR2_X1  g0320(.A(new_n520), .B(KEYINPUT12), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n205), .A2(G20), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n491), .A2(G68), .A3(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n443), .A2(new_n223), .ZN(new_n524));
  OAI22_X1  g0324(.A1(new_n487), .A2(new_n492), .B1(new_n206), .B2(G68), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n278), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT11), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n521), .B(new_n523), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  AND2_X1   g0328(.A1(new_n526), .A2(new_n527), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  NOR4_X1   g0331(.A1(new_n298), .A2(new_n468), .A3(new_n473), .A4(new_n301), .ZN(new_n532));
  AOI21_X1  g0332(.A(KEYINPUT65), .B1(new_n304), .B2(new_n469), .ZN(new_n533));
  OAI21_X1  g0333(.A(KEYINPUT70), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OR2_X1    g0334(.A1(G226), .A2(G1698), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(G232), .B2(new_n402), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n434), .B1(new_n536), .B2(new_n256), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n537), .A2(new_n298), .B1(new_n470), .B2(G238), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT70), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n474), .A2(new_n539), .A3(new_n475), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n534), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT13), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT13), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n534), .A2(new_n538), .A3(new_n540), .A4(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT14), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n546), .A3(G169), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n542), .A2(G179), .A3(new_n544), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n546), .B1(new_n545), .B2(G169), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n531), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n545), .A2(G200), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n542), .A2(G190), .A3(new_n544), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n552), .A2(new_n530), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n463), .A2(G232), .A3(new_n402), .ZN(new_n556));
  INV_X1    g0356(.A(new_n249), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n556), .B1(new_n463), .B2(new_n557), .ZN(new_n558));
  NOR3_X1   g0358(.A1(new_n256), .A2(new_n218), .A3(new_n402), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n298), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n474), .A2(new_n475), .B1(G244), .B2(new_n470), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(G200), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n491), .A2(G77), .A3(new_n522), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(G77), .B2(new_n280), .ZN(new_n565));
  NAND2_X1  g0365(.A1(G20), .A2(G77), .ZN(new_n566));
  OAI221_X1 g0366(.A(new_n566), .B1(new_n480), .B2(new_n487), .C1(new_n454), .C2(new_n443), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n565), .B1(new_n278), .B2(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n563), .B(new_n568), .C1(new_n376), .C2(new_n562), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n568), .B1(new_n562), .B2(new_n457), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n560), .A2(new_n451), .A3(new_n561), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n551), .A2(new_n555), .A3(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n519), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT76), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n499), .A2(new_n522), .ZN(new_n577));
  AOI211_X1 g0377(.A(new_n350), .B(new_n278), .C1(new_n577), .C2(KEYINPUT74), .ZN(new_n578));
  OR2_X1    g0378(.A1(new_n577), .A2(KEYINPUT74), .ZN(new_n579));
  INV_X1    g0379(.A(new_n499), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n578), .A2(new_n579), .B1(new_n350), .B2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  AND2_X1   g0382(.A1(new_n260), .A2(new_n262), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n265), .A2(new_n266), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n391), .B(new_n206), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(G68), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n391), .B1(new_n422), .B2(new_n206), .ZN(new_n587));
  OAI21_X1  g0387(.A(KEYINPUT73), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n583), .A2(new_n584), .ZN(new_n589));
  OAI21_X1  g0389(.A(KEYINPUT7), .B1(new_n589), .B2(G20), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT73), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n590), .A2(new_n591), .A3(G68), .A4(new_n585), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n482), .A2(new_n217), .ZN(new_n594));
  NOR2_X1   g0394(.A1(G58), .A2(G68), .ZN(new_n595));
  OR2_X1    g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n596), .A2(G20), .B1(G159), .B2(new_n388), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(KEYINPUT16), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n283), .B1(new_n593), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(G68), .B1(new_n390), .B2(new_n392), .ZN(new_n601));
  AOI21_X1  g0401(.A(KEYINPUT16), .B1(new_n601), .B2(new_n597), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n582), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT75), .ZN(new_n605));
  NAND2_X1  g0405(.A1(G226), .A2(G1698), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n605), .B1(new_n422), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n606), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n291), .A2(KEYINPUT75), .A3(new_n263), .A4(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n402), .A2(G223), .ZN(new_n611));
  OAI22_X1  g0411(.A1(new_n422), .A2(new_n611), .B1(new_n252), .B2(new_n219), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n312), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n474), .A2(new_n475), .B1(G232), .B2(new_n470), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(G169), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n612), .B1(new_n607), .B2(new_n609), .ZN(new_n618));
  OAI211_X1 g0418(.A(G179), .B(new_n615), .C1(new_n618), .C2(new_n312), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(KEYINPUT18), .B1(new_n604), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(G20), .B1(new_n291), .B2(new_n263), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n217), .B1(new_n623), .B2(new_n391), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n591), .B1(new_n624), .B2(new_n590), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n586), .A2(KEYINPUT73), .A3(new_n587), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n599), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n627), .A2(new_n278), .A3(new_n603), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n448), .B1(new_n614), .B2(new_n616), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n376), .B(new_n615), .C1(new_n618), .C2(new_n312), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n628), .A2(new_n631), .A3(new_n581), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT17), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n604), .A2(KEYINPUT17), .A3(new_n631), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT18), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n598), .B1(new_n588), .B2(new_n592), .ZN(new_n637));
  NOR3_X1   g0437(.A1(new_n637), .A2(new_n283), .A3(new_n602), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n636), .B(new_n620), .C1(new_n638), .C2(new_n582), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n622), .A2(new_n634), .A3(new_n635), .A4(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n575), .A2(new_n576), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n550), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n643), .A2(new_n548), .A3(new_n547), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n554), .B1(new_n644), .B2(new_n531), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n645), .A2(new_n512), .A3(new_n518), .A4(new_n573), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT76), .B1(new_n646), .B2(new_n640), .ZN(new_n647));
  AOI211_X1 g0447(.A(new_n339), .B(new_n462), .C1(new_n642), .C2(new_n647), .ZN(G372));
  NAND2_X1  g0448(.A1(new_n642), .A2(new_n647), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n447), .B1(new_n429), .B2(new_n448), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT89), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n447), .B(KEYINPUT89), .C1(new_n429), .C2(new_n448), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(new_n430), .A3(new_n653), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n395), .A2(new_n458), .A3(new_n459), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(new_n655), .A3(new_n456), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT26), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(KEYINPUT90), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT90), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n656), .A2(new_n660), .A3(new_n657), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n449), .A2(new_n456), .A3(KEYINPUT26), .A4(new_n655), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n659), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n456), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n655), .B1(new_n414), .B2(new_n410), .ZN(new_n665));
  AND4_X1   g0465(.A1(new_n338), .A2(new_n665), .A3(new_n654), .A4(new_n456), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n327), .A2(new_n287), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n374), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n664), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n663), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n649), .A2(new_n670), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n622), .A2(new_n639), .ZN(new_n672));
  AOI21_X1  g0472(.A(KEYINPUT17), .B1(new_n604), .B2(new_n631), .ZN(new_n673));
  AND4_X1   g0473(.A1(KEYINPUT17), .A2(new_n628), .A3(new_n581), .A4(new_n631), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n572), .ZN(new_n677));
  AOI22_X1  g0477(.A1(new_n555), .A2(new_n677), .B1(new_n644), .B2(new_n531), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n672), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n517), .B1(new_n679), .B2(new_n512), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n671), .A2(new_n680), .ZN(G369));
  NAND3_X1  g0481(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G213), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(G343), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n364), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  AND3_X1   g0489(.A1(new_n374), .A2(new_n377), .A3(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n374), .A2(new_n689), .ZN(new_n691));
  OAI21_X1  g0491(.A(G330), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  OR2_X1    g0492(.A1(new_n692), .A2(KEYINPUT91), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(KEYINPUT91), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n331), .A2(new_n334), .A3(new_n687), .ZN(new_n696));
  INV_X1    g0496(.A(new_n687), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n332), .A2(new_n333), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n696), .B1(new_n339), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n371), .A2(new_n373), .ZN(new_n701));
  INV_X1    g0501(.A(new_n368), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n687), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n326), .A2(new_n703), .A3(new_n338), .A4(new_n335), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n327), .A2(new_n287), .A3(new_n697), .ZN(new_n705));
  AOI21_X1  g0505(.A(KEYINPUT92), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n704), .A2(KEYINPUT92), .A3(new_n705), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n700), .B1(new_n706), .B2(new_n708), .ZN(G399));
  INV_X1    g0509(.A(new_n209), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(G41), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n249), .A2(G116), .A3(new_n440), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(G1), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n215), .B2(new_n712), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT28), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT30), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n406), .A2(new_n400), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n298), .B1(new_n718), .B2(new_n405), .ZN(new_n719));
  INV_X1    g0519(.A(new_n313), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n308), .A2(new_n347), .A3(G179), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n317), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n719), .A2(new_n722), .A3(new_n346), .A4(new_n398), .ZN(new_n723));
  INV_X1    g0523(.A(new_n429), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n717), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n722), .A2(new_n346), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n726), .A2(KEYINPUT30), .A3(new_n409), .A4(new_n429), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n320), .A2(G179), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n724), .A2(new_n369), .A3(new_n408), .A4(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n725), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n730), .A2(KEYINPUT31), .A3(new_n687), .ZN(new_n731));
  AOI21_X1  g0531(.A(KEYINPUT31), .B1(new_n730), .B2(new_n687), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n461), .A2(new_n374), .A3(new_n377), .A4(new_n697), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n733), .B1(new_n734), .B2(new_n339), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n735), .A2(G330), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT94), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n326), .A2(new_n335), .A3(new_n374), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(new_n666), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n456), .A2(KEYINPUT93), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n724), .A2(new_n457), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT93), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n741), .A2(new_n742), .A3(new_n452), .A4(new_n455), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n449), .A2(new_n456), .A3(new_n657), .A4(new_n655), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n746), .B1(KEYINPUT26), .B2(new_n656), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n739), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n737), .B1(new_n748), .B2(new_n697), .ZN(new_n749));
  AOI211_X1 g0549(.A(KEYINPUT94), .B(new_n687), .C1(new_n739), .C2(new_n747), .ZN(new_n750));
  OAI21_X1  g0550(.A(KEYINPUT29), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n670), .A2(new_n697), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT29), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n736), .B1(new_n751), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n716), .B1(new_n755), .B2(G1), .ZN(G364));
  INV_X1    g0556(.A(G13), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n205), .B1(new_n758), .B2(G45), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n711), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n209), .A2(new_n463), .ZN(new_n762));
  INV_X1    g0562(.A(G355), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n762), .A2(new_n763), .B1(G116), .B2(new_n209), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n422), .A2(new_n209), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT95), .Z(new_n766));
  NOR2_X1   g0566(.A1(new_n215), .A2(G45), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n767), .B1(new_n245), .B2(G45), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n764), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G13), .A2(G33), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  XOR2_X1   g0572(.A(new_n772), .B(KEYINPUT96), .Z(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n212), .B1(G20), .B2(new_n457), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n761), .B1(new_n769), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n206), .A2(new_n451), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n376), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n206), .A2(G179), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n783), .A2(new_n376), .A3(G200), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n782), .A2(new_n492), .B1(new_n784), .B2(new_n225), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n376), .A2(G179), .A3(G200), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n206), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n783), .A2(G190), .A3(G200), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n787), .A2(new_n382), .B1(new_n788), .B2(new_n219), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G190), .A2(G200), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n779), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n779), .A2(G190), .A3(new_n448), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n463), .B1(new_n792), .B2(new_n223), .C1(new_n482), .C2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(KEYINPUT32), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n783), .A2(new_n791), .ZN(new_n796));
  INV_X1    g0596(.A(G159), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n796), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n799), .A2(KEYINPUT32), .A3(G159), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n794), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n780), .A2(G190), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n802), .A2(KEYINPUT97), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n802), .A2(KEYINPUT97), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n790), .B(new_n801), .C1(new_n217), .C2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n788), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n781), .A2(G326), .B1(new_n807), .B2(G303), .ZN(new_n808));
  INV_X1    g0608(.A(G283), .ZN(new_n809));
  INV_X1    g0609(.A(G294), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n808), .B1(new_n809), .B2(new_n784), .C1(new_n810), .C2(new_n787), .ZN(new_n811));
  INV_X1    g0611(.A(new_n792), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G311), .A2(new_n812), .B1(new_n799), .B2(G329), .ZN(new_n813));
  INV_X1    g0613(.A(G322), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n813), .B(new_n256), .C1(new_n814), .C2(new_n793), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n805), .ZN(new_n817));
  XNOR2_X1  g0617(.A(KEYINPUT99), .B(KEYINPUT33), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(G317), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  AOI22_X1  g0620(.A1(KEYINPUT98), .A2(new_n806), .B1(new_n816), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(KEYINPUT98), .B2(new_n806), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n778), .B1(new_n822), .B2(new_n775), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n690), .A2(new_n691), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n823), .B1(new_n824), .B2(new_n773), .ZN(new_n825));
  INV_X1    g0625(.A(new_n761), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n824), .B2(G330), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n825), .B1(new_n695), .B2(new_n827), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT100), .Z(G396));
  NOR2_X1   g0629(.A1(new_n784), .A2(new_n219), .ZN(new_n830));
  INV_X1    g0630(.A(G303), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n782), .A2(new_n831), .B1(new_n788), .B2(new_n225), .ZN(new_n832));
  INV_X1    g0632(.A(new_n787), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n830), .B(new_n832), .C1(G97), .C2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(G311), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n792), .A2(new_n360), .B1(new_n796), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n793), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n463), .B(new_n836), .C1(G294), .C2(new_n837), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n834), .B(new_n838), .C1(new_n809), .C2(new_n805), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT102), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n837), .A2(G143), .B1(new_n812), .B2(G159), .ZN(new_n841));
  INV_X1    g0641(.A(G137), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n841), .B1(new_n842), .B2(new_n782), .C1(new_n805), .C2(new_n486), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT34), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n843), .A2(new_n844), .ZN(new_n846));
  INV_X1    g0646(.A(G132), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n589), .B1(new_n847), .B2(new_n796), .ZN(new_n848));
  INV_X1    g0648(.A(new_n784), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n807), .A2(G50), .B1(new_n849), .B2(G68), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n482), .B2(new_n787), .ZN(new_n851));
  NOR4_X1   g0651(.A1(new_n845), .A2(new_n846), .A3(new_n848), .A4(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n775), .B1(new_n840), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n775), .A2(new_n770), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n854), .B(KEYINPUT101), .Z(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n826), .B1(new_n856), .B2(new_n223), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n569), .B1(new_n568), .B2(new_n697), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n572), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n677), .A2(new_n697), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n853), .B(new_n857), .C1(new_n862), .C2(new_n771), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n687), .B(new_n861), .C1(new_n663), .C2(new_n669), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n864), .A2(KEYINPUT103), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n752), .A2(new_n861), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n865), .B(new_n866), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n867), .A2(new_n736), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n826), .B1(new_n867), .B2(new_n736), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n863), .B1(new_n868), .B2(new_n869), .ZN(G384));
  OAI21_X1  g0670(.A(new_n597), .B1(new_n625), .B2(new_n626), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT16), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n582), .B1(new_n873), .B2(new_n600), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n632), .B1(new_n874), .B2(new_n685), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n874), .A2(new_n621), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT37), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n620), .B1(new_n638), .B2(new_n582), .ZN(new_n878));
  INV_X1    g0678(.A(new_n685), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n638), .B2(new_n582), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT37), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n878), .A2(new_n880), .A3(new_n881), .A4(new_n632), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n877), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n627), .A2(new_n278), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT16), .B1(new_n593), .B2(new_n597), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n581), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n879), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n640), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n883), .A2(KEYINPUT38), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n878), .A2(new_n880), .A3(new_n632), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT37), .ZN(new_n892));
  INV_X1    g0692(.A(new_n880), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n882), .A2(new_n892), .B1(new_n640), .B2(new_n893), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n890), .B(KEYINPUT105), .C1(KEYINPUT38), .C2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT39), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT105), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n883), .A2(new_n889), .A3(new_n897), .A4(KEYINPUT38), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n895), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n644), .A2(new_n531), .A3(new_n697), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT38), .ZN(new_n902));
  AND4_X1   g0702(.A1(new_n881), .A2(new_n878), .A3(new_n880), .A4(new_n632), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n887), .B(new_n632), .C1(new_n621), .C2(new_n874), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n903), .B1(KEYINPUT37), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n887), .B1(new_n672), .B2(new_n675), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n902), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n907), .A2(KEYINPUT39), .A3(new_n890), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n899), .A2(new_n901), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n907), .A2(new_n890), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n551), .B(new_n555), .C1(new_n530), .C2(new_n697), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n531), .B(new_n687), .C1(new_n644), .C2(new_n554), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n860), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n910), .B(new_n913), .C1(new_n864), .C2(new_n914), .ZN(new_n915));
  OR2_X1    g0715(.A1(new_n672), .A2(new_n879), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n909), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n751), .A2(new_n754), .A3(new_n649), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n680), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n917), .B(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT40), .ZN(new_n921));
  INV_X1    g0721(.A(new_n890), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT38), .B1(new_n883), .B2(new_n889), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n861), .B1(new_n911), .B2(new_n912), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n735), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n921), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n735), .A2(KEYINPUT40), .A3(new_n925), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n895), .A2(new_n898), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n649), .A2(new_n735), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n930), .A2(new_n931), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n932), .A2(G330), .A3(new_n933), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n920), .A2(new_n934), .B1(new_n205), .B2(new_n758), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT106), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n935), .A2(new_n936), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n920), .A2(new_n934), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AOI211_X1 g0740(.A(new_n360), .B(new_n214), .C1(new_n387), .C2(KEYINPUT35), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(KEYINPUT35), .B2(new_n387), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT36), .ZN(new_n943));
  NOR3_X1   g0743(.A1(new_n594), .A2(new_n215), .A3(new_n223), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n944), .A2(KEYINPUT104), .B1(new_n492), .B2(G68), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(KEYINPUT104), .B2(new_n944), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n946), .A2(G1), .A3(new_n757), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n940), .A2(new_n943), .A3(new_n947), .ZN(G367));
  OR2_X1    g0748(.A1(new_n447), .A2(new_n697), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n654), .A2(new_n456), .A3(new_n949), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n456), .A2(new_n949), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n774), .ZN(new_n954));
  INV_X1    g0754(.A(new_n766), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n955), .A2(new_n237), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n776), .B1(new_n209), .B2(new_n454), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n761), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n589), .B1(G311), .B2(new_n781), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n833), .A2(new_n249), .B1(new_n849), .B2(G97), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n959), .B(new_n960), .C1(new_n805), .C2(new_n810), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n837), .A2(G303), .B1(new_n799), .B2(G317), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n807), .A2(KEYINPUT46), .A3(G116), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT46), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n788), .B2(new_n360), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n812), .A2(G283), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n962), .A2(new_n963), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n805), .A2(new_n797), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n833), .A2(G68), .B1(new_n849), .B2(G77), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n781), .A2(G143), .B1(new_n807), .B2(G58), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n256), .B1(new_n837), .B2(G150), .ZN(new_n971));
  AOI22_X1  g0771(.A1(G50), .A2(new_n812), .B1(new_n799), .B2(G137), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n969), .A2(new_n970), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n961), .A2(new_n967), .B1(new_n968), .B2(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT47), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n958), .B1(new_n975), .B2(new_n775), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n954), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT109), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n711), .B(KEYINPUT41), .Z(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n704), .A2(new_n705), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT92), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n395), .A2(new_n687), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n665), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n655), .A2(new_n687), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n983), .A2(new_n707), .A3(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT108), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT44), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n990), .A2(new_n991), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n983), .A2(new_n707), .A3(new_n988), .A4(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n992), .A2(new_n993), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n987), .B1(new_n708), .B2(new_n706), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT45), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI211_X1 g0799(.A(KEYINPUT45), .B(new_n987), .C1(new_n708), .C2(new_n706), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n996), .A2(new_n1001), .A3(new_n700), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n700), .B1(new_n996), .B2(new_n1001), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n699), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n703), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n704), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n695), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1007), .A2(new_n693), .A3(new_n694), .A4(new_n704), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n755), .A2(new_n1011), .ZN(new_n1012));
  NOR3_X1   g0812(.A1(new_n1003), .A2(new_n1004), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n755), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n980), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n759), .ZN(new_n1016));
  OAI21_X1  g0816(.A(KEYINPUT42), .B1(new_n704), .B2(new_n988), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n326), .A2(new_n335), .B1(new_n414), .B2(new_n410), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n697), .B1(new_n1018), .B2(new_n655), .ZN(new_n1019));
  AND2_X1   g0819(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(KEYINPUT107), .ZN(new_n1021));
  OR3_X1    g0821(.A1(new_n704), .A2(new_n988), .A3(KEYINPUT42), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT43), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1020), .A2(KEYINPUT107), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1024), .A2(new_n1025), .A3(new_n953), .A4(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n700), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n987), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n953), .A2(new_n1025), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n952), .A2(KEYINPUT43), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1032), .B(new_n1033), .C1(new_n1023), .C2(new_n1026), .ZN(new_n1034));
  AND3_X1   g0834(.A1(new_n1028), .A2(new_n1031), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1031), .B1(new_n1028), .B2(new_n1034), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n978), .B1(new_n1016), .B2(new_n1037), .ZN(new_n1038));
  AND2_X1   g0838(.A1(new_n755), .A2(new_n1011), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n996), .A2(new_n1001), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n1029), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1039), .A2(new_n1041), .A3(new_n1002), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n979), .B1(new_n1042), .B2(new_n755), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n978), .B(new_n1037), .C1(new_n1043), .C2(new_n760), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n977), .B1(new_n1038), .B2(new_n1045), .ZN(G387));
  OAI21_X1  g0846(.A(new_n766), .B1(new_n234), .B2(new_n305), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n713), .B2(new_n762), .ZN(new_n1048));
  OR3_X1    g0848(.A1(new_n480), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1049));
  AOI21_X1  g0849(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1050));
  OAI21_X1  g0850(.A(KEYINPUT50), .B1(new_n480), .B2(G50), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1049), .A2(new_n713), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n1048), .A2(new_n1052), .B1(new_n225), .B2(new_n710), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n761), .B1(new_n1053), .B2(new_n777), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n817), .A2(new_n499), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n782), .A2(new_n797), .B1(new_n454), .B2(new_n787), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n788), .A2(new_n223), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n793), .A2(new_n492), .B1(new_n796), .B2(new_n486), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(G68), .B2(new_n812), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n422), .B1(G97), .B2(new_n849), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1055), .A2(new_n1058), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n589), .B1(G326), .B2(new_n799), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n837), .A2(G317), .B1(new_n812), .B2(G303), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1064), .B1(new_n814), .B2(new_n782), .C1(new_n805), .C2(new_n835), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT48), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n833), .A2(G283), .B1(new_n807), .B2(G294), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT49), .Z(new_n1071));
  INV_X1    g0871(.A(KEYINPUT110), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1063), .B1(new_n360), .B2(new_n784), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1062), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1054), .B1(new_n1075), .B2(new_n775), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT111), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1005), .A2(new_n774), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1077), .A2(new_n1078), .B1(new_n760), .B2(new_n1011), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1012), .A2(new_n711), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n755), .A2(new_n1011), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1079), .B1(new_n1080), .B2(new_n1081), .ZN(G393));
  NAND3_X1  g0882(.A1(new_n1041), .A2(new_n760), .A3(new_n1002), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n775), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G317), .A2(new_n781), .B1(new_n837), .B2(G311), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT52), .Z(new_n1086));
  OAI22_X1  g0886(.A1(new_n788), .A2(new_n809), .B1(new_n796), .B2(new_n814), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT112), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n817), .A2(G303), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n256), .B1(new_n792), .B2(new_n810), .C1(new_n225), .C2(new_n784), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(G116), .B2(new_n833), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1086), .A2(new_n1088), .A3(new_n1089), .A4(new_n1091), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n782), .A2(new_n486), .B1(new_n797), .B2(new_n793), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT51), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n817), .A2(G50), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n792), .A2(new_n480), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n1096), .B(new_n422), .C1(G143), .C2(new_n799), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n788), .A2(new_n217), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n830), .B(new_n1098), .C1(G77), .C2(new_n833), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1094), .A2(new_n1095), .A3(new_n1097), .A4(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1084), .B1(new_n1092), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n766), .A2(new_n242), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n777), .B1(G97), .B2(new_n710), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n826), .B(new_n1101), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n987), .B2(new_n773), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1083), .A2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1013), .A2(new_n712), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1012), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1106), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(G390));
  NAND2_X1  g0910(.A1(new_n899), .A2(new_n908), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n770), .ZN(new_n1112));
  INV_X1    g0912(.A(G128), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n782), .A2(new_n1113), .B1(new_n847), .B2(new_n793), .ZN(new_n1114));
  OR2_X1    g0914(.A1(new_n1114), .A2(KEYINPUT116), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(KEYINPUT116), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1115), .B(new_n1116), .C1(new_n805), .C2(new_n842), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n788), .A2(new_n486), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1118), .B(KEYINPUT53), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(KEYINPUT54), .B(G143), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n812), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n256), .B1(new_n799), .B2(G125), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n833), .A2(G159), .B1(new_n849), .B2(G50), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1119), .A2(new_n1122), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1117), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1127), .A2(KEYINPUT117), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n817), .A2(new_n249), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n792), .A2(new_n382), .B1(new_n796), .B2(new_n810), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n463), .B(new_n1130), .C1(G116), .C2(new_n837), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n807), .A2(G87), .B1(new_n849), .B2(G68), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(G77), .A2(new_n833), .B1(new_n781), .B2(G283), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1129), .A2(new_n1131), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT117), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1134), .B1(new_n1126), .B2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n775), .B1(new_n1128), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n826), .B1(new_n856), .B2(new_n580), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1112), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n735), .A2(G330), .A3(new_n862), .A4(new_n913), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n895), .A2(new_n900), .A3(new_n898), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n859), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n749), .A2(new_n750), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1143), .B1(new_n1144), .B2(new_n860), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1142), .B1(new_n1145), .B2(new_n913), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n913), .B1(new_n864), .B2(new_n914), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n1147), .A2(new_n900), .B1(new_n908), .B2(new_n899), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1141), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n687), .B1(new_n739), .B2(new_n747), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1150), .B(new_n737), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n859), .B(new_n913), .C1(new_n1151), .C2(new_n914), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1142), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n687), .B1(new_n663), .B2(new_n669), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n914), .B1(new_n1155), .B2(new_n862), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n913), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n900), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n1111), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1154), .A2(new_n1159), .A3(new_n1140), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1149), .A2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1139), .B1(new_n1161), .B2(new_n759), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n649), .A2(new_n736), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(KEYINPUT113), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT113), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n649), .A2(new_n736), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n1167), .A2(new_n918), .A3(new_n680), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n860), .B1(new_n752), .B2(new_n1143), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n735), .A2(G330), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1157), .B1(new_n1170), .B2(new_n861), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(new_n1140), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1173), .B(KEYINPUT114), .C1(new_n1145), .C2(new_n1172), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n859), .B1(new_n1151), .B2(new_n914), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT114), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1175), .A2(new_n1176), .A3(new_n1140), .A4(new_n1171), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1168), .A2(new_n1174), .A3(new_n1177), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n1146), .A2(new_n1148), .A3(new_n1141), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1140), .B1(new_n1154), .B2(new_n1159), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1178), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT115), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1161), .A2(KEYINPUT115), .A3(new_n1178), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1174), .A2(new_n1177), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1186), .A2(new_n1149), .A3(new_n1160), .A4(new_n1168), .ZN(new_n1187));
  AND2_X1   g0987(.A1(new_n1187), .A2(new_n711), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1162), .B1(new_n1185), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(G378));
  OAI21_X1  g0990(.A(new_n1168), .B1(new_n1161), .B2(new_n1178), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n926), .B1(new_n907), .B2(new_n890), .ZN(new_n1192));
  OAI21_X1  g0992(.A(G330), .B1(new_n1192), .B2(KEYINPUT40), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n895), .A2(new_n898), .A3(new_n928), .ZN(new_n1194));
  OAI21_X1  g0994(.A(KEYINPUT120), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT120), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n927), .A2(new_n1196), .A3(G330), .A4(new_n929), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n513), .A2(new_n685), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1198), .B(KEYINPUT55), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n519), .B(new_n1199), .ZN(new_n1200));
  XOR2_X1   g1000(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1201));
  XNOR2_X1  g1001(.A(new_n1200), .B(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1195), .A2(new_n1197), .A3(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1205), .A2(new_n1196), .A3(new_n1202), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1204), .A2(KEYINPUT121), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n917), .A2(KEYINPUT122), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT122), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n909), .A2(new_n915), .A3(new_n1209), .A4(new_n916), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1208), .A2(new_n1210), .ZN(new_n1211));
  AND2_X1   g1011(.A1(new_n1207), .A2(new_n1211), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1207), .A2(new_n1211), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1191), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT57), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n917), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1204), .A2(new_n1217), .A3(new_n1206), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1217), .B1(new_n1204), .B2(new_n1206), .ZN(new_n1220));
  NOR3_X1   g1020(.A1(new_n1219), .A2(new_n1220), .A3(new_n1215), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n712), .B1(new_n1221), .B2(new_n1191), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1216), .A2(new_n1222), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1204), .A2(KEYINPUT121), .A3(new_n1206), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n1208), .A2(new_n1210), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1207), .A2(new_n1211), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n759), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT123), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n761), .B1(new_n855), .B2(G50), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n589), .A2(G41), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n492), .B1(G33), .B2(G41), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n782), .A2(new_n360), .B1(new_n784), .B2(new_n482), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n1057), .B(new_n1234), .C1(G68), .C2(new_n833), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n817), .A2(G97), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n793), .A2(new_n225), .B1(new_n796), .B2(new_n809), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n431), .B2(new_n812), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1235), .A2(new_n1236), .A3(new_n1231), .A4(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT58), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1233), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n793), .A2(new_n1113), .B1(new_n792), .B2(new_n842), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(G150), .B2(new_n833), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n781), .A2(G125), .B1(new_n807), .B2(new_n1121), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1243), .B(new_n1244), .C1(new_n805), .C2(new_n847), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1245), .A2(KEYINPUT59), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(KEYINPUT59), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n849), .A2(G159), .ZN(new_n1248));
  AOI211_X1 g1048(.A(G33), .B(G41), .C1(new_n799), .C2(G124), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1247), .A2(new_n1248), .A3(new_n1249), .ZN(new_n1250));
  OAI221_X1 g1050(.A(new_n1241), .B1(new_n1240), .B2(new_n1239), .C1(new_n1246), .C2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1230), .B1(new_n1251), .B2(new_n775), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n1203), .B2(new_n771), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(new_n1253), .B(KEYINPUT119), .ZN(new_n1254));
  NOR3_X1   g1054(.A1(new_n1228), .A2(new_n1229), .A3(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n760), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1254), .ZN(new_n1257));
  AOI21_X1  g1057(.A(KEYINPUT123), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1223), .B1(new_n1255), .B2(new_n1258), .ZN(G375));
  INV_X1    g1059(.A(KEYINPUT126), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1174), .A2(new_n1177), .A3(new_n760), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n826), .B1(new_n856), .B2(new_n217), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n817), .A2(G116), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n793), .A2(new_n809), .B1(new_n796), .B2(new_n831), .ZN(new_n1264));
  AOI211_X1 g1064(.A(new_n463), .B(new_n1264), .C1(new_n249), .C2(new_n812), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n833), .A2(new_n431), .B1(new_n849), .B2(G77), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n781), .A2(G294), .B1(new_n807), .B2(G97), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1263), .A2(new_n1265), .A3(new_n1266), .A4(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT124), .ZN(new_n1269));
  OAI22_X1  g1069(.A1(new_n788), .A2(new_n797), .B1(new_n796), .B2(new_n1113), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n817), .A2(new_n1121), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1271), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n781), .A2(G132), .B1(new_n849), .B2(G58), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n837), .A2(G137), .B1(new_n812), .B2(G150), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n833), .A2(G50), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1273), .A2(new_n1274), .A3(new_n589), .A4(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1268), .B1(new_n1272), .B2(new_n1276), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1277), .A2(KEYINPUT125), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(KEYINPUT125), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n775), .ZN(new_n1280));
  OAI221_X1 g1080(.A(new_n1262), .B1(new_n1278), .B2(new_n1280), .C1(new_n913), .C2(new_n771), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1260), .B1(new_n1261), .B2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1261), .A2(new_n1260), .A3(new_n1281), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1168), .B1(new_n1174), .B2(new_n1177), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1178), .A2(new_n980), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1285), .B1(new_n1286), .B2(new_n1287), .ZN(G381));
  OAI21_X1  g1088(.A(new_n1229), .B1(new_n1228), .B2(new_n1254), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1256), .A2(KEYINPUT123), .A3(new_n1257), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1291), .A2(new_n1189), .A3(new_n1223), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1037), .B1(new_n1043), .B2(new_n760), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(KEYINPUT109), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1044), .ZN(new_n1296));
  OR2_X1    g1096(.A1(G393), .A2(G396), .ZN(new_n1297));
  NOR4_X1   g1097(.A1(G381), .A2(G390), .A3(new_n1297), .A4(G384), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1293), .A2(new_n1296), .A3(new_n977), .A4(new_n1298), .ZN(G407));
  OAI211_X1 g1099(.A(G407), .B(G213), .C1(G343), .C2(new_n1292), .ZN(G409));
  AND2_X1   g1100(.A1(new_n686), .A2(G213), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n917), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1303), .A2(new_n760), .A3(new_n1218), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1257), .ZN(new_n1305));
  AOI22_X1  g1105(.A1(new_n1226), .A2(new_n1227), .B1(new_n1187), .B2(new_n1168), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1305), .B1(new_n1306), .B2(new_n980), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1301), .B1(new_n1307), .B2(new_n1189), .ZN(new_n1308));
  AOI22_X1  g1108(.A1(new_n1289), .A2(new_n1290), .B1(new_n1216), .B2(new_n1222), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1308), .B1(new_n1309), .B2(new_n1189), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1286), .B1(KEYINPUT60), .B2(new_n1178), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1174), .A2(new_n1177), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1168), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1312), .A2(new_n1313), .A3(KEYINPUT60), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n711), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1284), .ZN(new_n1316));
  OAI22_X1  g1116(.A1(new_n1311), .A2(new_n1315), .B1(new_n1316), .B2(new_n1282), .ZN(new_n1317));
  INV_X1    g1117(.A(G384), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1285), .B(G384), .C1(new_n1311), .C2(new_n1315), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1301), .A2(G2897), .ZN(new_n1321));
  AND3_X1   g1121(.A1(new_n1319), .A2(new_n1320), .A3(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1321), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(KEYINPUT61), .B1(new_n1310), .B2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(G375), .A2(G378), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT62), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1328), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1326), .A2(new_n1327), .A3(new_n1308), .A4(new_n1329), .ZN(new_n1330));
  OAI211_X1 g1130(.A(new_n1308), .B(new_n1329), .C1(new_n1309), .C2(new_n1189), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(KEYINPUT62), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1325), .A2(new_n1330), .A3(new_n1332), .ZN(new_n1333));
  XOR2_X1   g1133(.A(G393), .B(G396), .Z(new_n1334));
  INV_X1    g1134(.A(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(G390), .B1(new_n1296), .B2(new_n977), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n977), .ZN(new_n1337));
  AOI211_X1 g1137(.A(new_n1337), .B(new_n1109), .C1(new_n1295), .C2(new_n1044), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1335), .B1(new_n1336), .B2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(G387), .A2(new_n1109), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1296), .A2(new_n977), .A3(G390), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1340), .A2(new_n1334), .A3(new_n1341), .ZN(new_n1342));
  AND2_X1   g1142(.A1(new_n1339), .A2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1333), .A2(new_n1344), .ZN(new_n1345));
  NAND4_X1  g1145(.A1(new_n1326), .A2(KEYINPUT63), .A3(new_n1308), .A4(new_n1329), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT63), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1331), .A2(new_n1347), .ZN(new_n1348));
  NAND4_X1  g1148(.A1(new_n1343), .A2(new_n1325), .A3(new_n1346), .A4(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1345), .A2(new_n1349), .ZN(G405));
  NOR2_X1   g1150(.A1(new_n1309), .A2(new_n1189), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1329), .B1(new_n1293), .B2(new_n1351), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1326), .A2(new_n1292), .A3(new_n1328), .ZN(new_n1353));
  AND3_X1   g1153(.A1(new_n1343), .A2(new_n1352), .A3(new_n1353), .ZN(new_n1354));
  AOI21_X1  g1154(.A(new_n1343), .B1(new_n1352), .B2(new_n1353), .ZN(new_n1355));
  NOR2_X1   g1155(.A1(new_n1354), .A2(new_n1355), .ZN(G402));
endmodule


