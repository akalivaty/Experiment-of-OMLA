//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1 1 0 1 1 0 0 1 0 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 1 1 1 1 0 0 0 1 0 0 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n883, new_n884,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952;
  INV_X1    g000(.A(KEYINPUT29), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT26), .B(G101), .Z(new_n188));
  INV_X1    g002(.A(G237), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G210), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n188), .B(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G116), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT68), .B1(new_n195), .B2(G119), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT68), .ZN(new_n197));
  INV_X1    g011(.A(G119), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(G116), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n195), .A2(G119), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n196), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT2), .B(G113), .ZN(new_n202));
  XNOR2_X1  g016(.A(new_n201), .B(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  OR2_X1    g018(.A1(KEYINPUT0), .A2(G128), .ZN(new_n205));
  NAND2_X1  g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(G143), .B(G146), .ZN(new_n208));
  MUX2_X1   g022(.A(new_n207), .B(new_n206), .S(new_n208), .Z(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  AND2_X1   g024(.A1(KEYINPUT66), .A2(G137), .ZN(new_n211));
  NOR2_X1   g025(.A1(KEYINPUT66), .A2(G137), .ZN(new_n212));
  OAI211_X1 g026(.A(KEYINPUT11), .B(G134), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT67), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT66), .B(G137), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n216), .A2(KEYINPUT67), .A3(KEYINPUT11), .A4(G134), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n219));
  INV_X1    g033(.A(G134), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n220), .A2(G137), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n219), .B1(new_n221), .B2(KEYINPUT11), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT11), .ZN(new_n223));
  OAI211_X1 g037(.A(KEYINPUT65), .B(new_n223), .C1(new_n220), .C2(G137), .ZN(new_n224));
  AOI22_X1  g038(.A1(new_n222), .A2(new_n224), .B1(new_n220), .B2(G137), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n218), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G131), .ZN(new_n227));
  INV_X1    g041(.A(G131), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n218), .A2(new_n228), .A3(new_n225), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n210), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G128), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n231), .A2(KEYINPUT1), .ZN(new_n232));
  INV_X1    g046(.A(G146), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G143), .ZN(new_n234));
  INV_X1    g048(.A(G143), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G146), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n232), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n231), .A2(new_n233), .A3(G143), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n235), .B(G146), .C1(new_n231), .C2(KEYINPUT1), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n237), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n216), .A2(G134), .ZN(new_n241));
  OAI21_X1  g055(.A(G131), .B1(new_n241), .B2(new_n221), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n229), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT64), .B1(new_n230), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT30), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n218), .A2(new_n228), .A3(new_n225), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n228), .B1(new_n218), .B2(new_n225), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n209), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(new_n243), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(KEYINPUT64), .A3(KEYINPUT30), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n204), .B1(new_n247), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n250), .A2(new_n204), .A3(new_n243), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n187), .B(new_n194), .C1(new_n253), .C2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n204), .B1(new_n250), .B2(new_n243), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT28), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n194), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT28), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n254), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n258), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n187), .A2(KEYINPUT70), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n263), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n258), .A2(new_n259), .A3(new_n265), .A4(new_n261), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n256), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(G472), .B1(new_n267), .B2(G902), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT30), .B1(new_n251), .B2(KEYINPUT64), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT64), .ZN(new_n270));
  AOI211_X1 g084(.A(new_n270), .B(new_n246), .C1(new_n250), .C2(new_n243), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n203), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n272), .A2(new_n254), .A3(new_n259), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT31), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n251), .A2(new_n203), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n260), .B1(new_n275), .B2(new_n254), .ZN(new_n276));
  INV_X1    g090(.A(new_n261), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n194), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n273), .A2(new_n274), .A3(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G472), .ZN(new_n280));
  INV_X1    g094(.A(G902), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n272), .A2(KEYINPUT31), .A3(new_n254), .A4(new_n259), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n279), .A2(new_n280), .A3(new_n281), .A4(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT32), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n282), .A2(new_n281), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n286), .A2(KEYINPUT32), .A3(new_n280), .A4(new_n279), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n268), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n231), .A2(G119), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(KEYINPUT72), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT23), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n198), .A2(G128), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT23), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n289), .A2(KEYINPUT72), .A3(new_n293), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n291), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G110), .ZN(new_n296));
  OR2_X1    g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n292), .A2(KEYINPUT71), .ZN(new_n298));
  MUX2_X1   g112(.A(KEYINPUT71), .B(new_n298), .S(new_n289), .Z(new_n299));
  XNOR2_X1  g113(.A(KEYINPUT24), .B(G110), .ZN(new_n300));
  OR2_X1    g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G125), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G140), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT73), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT73), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n305), .A2(new_n302), .A3(G140), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  OR2_X1    g121(.A1(new_n302), .A2(G140), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n307), .A2(KEYINPUT16), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT74), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n302), .A2(G140), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT16), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n309), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n311), .B1(new_n304), .B2(new_n306), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(KEYINPUT74), .A3(KEYINPUT16), .ZN(new_n317));
  AND3_X1   g131(.A1(new_n315), .A2(G146), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(G146), .B1(new_n315), .B2(new_n317), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n297), .B(new_n301), .C1(new_n318), .C2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT75), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n315), .A2(new_n317), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n233), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n315), .A2(G146), .A3(new_n317), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n325), .A2(new_n326), .A3(new_n297), .A4(new_n301), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n321), .A2(new_n327), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n308), .A2(new_n233), .A3(new_n303), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n295), .A2(new_n296), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n299), .A2(new_n300), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n324), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT22), .B(G137), .ZN(new_n335));
  AND3_X1   g149(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n336));
  XOR2_X1   g150(.A(new_n335), .B(new_n336), .Z(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n328), .A2(new_n333), .A3(new_n337), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(new_n281), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT25), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n337), .B1(new_n328), .B2(new_n333), .ZN(new_n344));
  INV_X1    g158(.A(new_n333), .ZN(new_n345));
  AOI211_X1 g159(.A(new_n345), .B(new_n338), .C1(new_n321), .C2(new_n327), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(KEYINPUT25), .A3(new_n281), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G217), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n350), .B1(G234), .B2(new_n281), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n351), .A2(G902), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n349), .A2(new_n351), .B1(new_n347), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n288), .A2(new_n353), .ZN(new_n354));
  OR2_X1    g168(.A1(new_n354), .A2(KEYINPUT76), .ZN(new_n355));
  INV_X1    g169(.A(G221), .ZN(new_n356));
  XOR2_X1   g170(.A(KEYINPUT9), .B(G234), .Z(new_n357));
  XNOR2_X1  g171(.A(new_n357), .B(KEYINPUT77), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n356), .B1(new_n358), .B2(new_n281), .ZN(new_n359));
  INV_X1    g173(.A(G104), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT3), .B1(new_n360), .B2(G107), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT3), .ZN(new_n362));
  INV_X1    g176(.A(G107), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(new_n363), .A3(G104), .ZN(new_n364));
  INV_X1    g178(.A(G101), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n360), .A2(G107), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n361), .A2(new_n364), .A3(new_n365), .A4(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n360), .A2(G107), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n363), .A2(G104), .ZN(new_n369));
  OAI21_X1  g183(.A(G101), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n240), .A2(new_n367), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n372));
  OR2_X1    g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n361), .A2(new_n364), .A3(new_n366), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G101), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n375), .A2(KEYINPUT78), .A3(KEYINPUT4), .A4(new_n367), .ZN(new_n376));
  NAND2_X1  g190(.A1(KEYINPUT78), .A2(KEYINPUT4), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n374), .A2(G101), .A3(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(new_n209), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n371), .A2(new_n372), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n373), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n248), .A2(new_n249), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n373), .A2(new_n379), .A3(new_n380), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n227), .A2(new_n229), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(G110), .B(G140), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n190), .A2(G227), .ZN(new_n388));
  XOR2_X1   g202(.A(new_n387), .B(new_n388), .Z(new_n389));
  NAND3_X1  g203(.A1(new_n383), .A2(new_n386), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n367), .A2(new_n370), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n391), .A2(new_n238), .A3(new_n237), .A4(new_n239), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n371), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n393), .B1(new_n248), .B2(new_n249), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT12), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n393), .B(KEYINPUT12), .C1(new_n248), .C2(new_n249), .ZN(new_n397));
  AOI22_X1  g211(.A1(new_n396), .A2(new_n397), .B1(new_n381), .B2(new_n382), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n390), .B(G469), .C1(new_n398), .C2(new_n389), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(KEYINPUT12), .B1(new_n385), .B2(new_n393), .ZN(new_n401));
  INV_X1    g215(.A(new_n397), .ZN(new_n402));
  OAI21_X1  g216(.A(KEYINPUT79), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n389), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n404), .B1(new_n381), .B2(new_n382), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT79), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n396), .A2(new_n406), .A3(new_n397), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n403), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n383), .A2(new_n386), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(new_n404), .ZN(new_n410));
  AOI21_X1  g224(.A(G902), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G469), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n400), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n412), .A2(new_n281), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n359), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  XOR2_X1   g231(.A(G110), .B(G122), .Z(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n203), .A2(new_n376), .A3(new_n378), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT5), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(new_n198), .A3(G116), .ZN(new_n422));
  OAI211_X1 g236(.A(G113), .B(new_n422), .C1(new_n201), .C2(new_n421), .ZN(new_n423));
  OR2_X1    g237(.A1(new_n201), .A2(new_n202), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n423), .A2(new_n424), .A3(new_n367), .A4(new_n370), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n419), .B1(new_n420), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n420), .A2(new_n425), .A3(new_n419), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(KEYINPUT6), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n240), .A2(new_n302), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n430), .B1(new_n210), .B2(new_n302), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n190), .A2(G224), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n431), .B(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT6), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n426), .A2(KEYINPUT80), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(KEYINPUT80), .B1(new_n426), .B2(new_n434), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n429), .B(new_n433), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT81), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n432), .A2(KEYINPUT7), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n431), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n438), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n423), .A2(new_n424), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n391), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n425), .ZN(new_n445));
  XOR2_X1   g259(.A(new_n418), .B(KEYINPUT8), .Z(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n431), .A2(new_n438), .A3(new_n439), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n442), .A2(new_n447), .A3(new_n428), .A4(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n437), .A2(new_n281), .A3(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(G210), .B1(G237), .B2(G902), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n437), .A2(new_n281), .A3(new_n451), .A4(new_n449), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(G214), .B1(G237), .B2(G902), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n417), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(G116), .B(G122), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n459), .B(new_n363), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(KEYINPUT85), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT88), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n231), .A2(G143), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT87), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n464), .B1(new_n235), .B2(G128), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n231), .A2(KEYINPUT87), .A3(G143), .ZN(new_n466));
  AOI211_X1 g280(.A(new_n462), .B(new_n463), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n466), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n235), .A2(G128), .ZN(new_n469));
  AOI21_X1  g283(.A(KEYINPUT88), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n220), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  XOR2_X1   g285(.A(KEYINPUT86), .B(KEYINPUT13), .Z(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n469), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n468), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n472), .A2(new_n469), .ZN(new_n475));
  OAI21_X1  g289(.A(G134), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n461), .A2(new_n471), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n231), .A2(KEYINPUT87), .A3(G143), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT87), .B1(new_n231), .B2(G143), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n469), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n462), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n468), .A2(KEYINPUT88), .A3(new_n469), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(G134), .A3(new_n483), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n471), .A2(new_n484), .A3(KEYINPUT89), .ZN(new_n485));
  AOI21_X1  g299(.A(KEYINPUT89), .B1(new_n471), .B2(new_n484), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n459), .A2(new_n363), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n195), .A2(KEYINPUT14), .A3(G122), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT14), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n489), .B1(new_n459), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n488), .B1(G107), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(KEYINPUT90), .B1(new_n487), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT89), .ZN(new_n494));
  NOR3_X1   g308(.A1(new_n467), .A2(new_n470), .A3(new_n220), .ZN(new_n495));
  AOI21_X1  g309(.A(G134), .B1(new_n482), .B2(new_n483), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n471), .A2(new_n484), .A3(KEYINPUT89), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n497), .A2(KEYINPUT90), .A3(new_n492), .A4(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n478), .B1(new_n493), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n358), .A2(G217), .A3(new_n190), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n502), .B(KEYINPUT91), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n497), .A2(new_n492), .A3(new_n498), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT90), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n499), .ZN(new_n508));
  INV_X1    g322(.A(new_n503), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(new_n509), .A3(new_n478), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n504), .A2(new_n281), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT92), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n509), .B1(new_n508), .B2(new_n478), .ZN(new_n514));
  AOI211_X1 g328(.A(new_n503), .B(new_n477), .C1(new_n507), .C2(new_n499), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(KEYINPUT92), .A3(new_n281), .ZN(new_n517));
  INV_X1    g331(.A(G478), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n518), .A2(KEYINPUT15), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n513), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  OR2_X1    g334(.A1(new_n511), .A2(new_n519), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT19), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n308), .A2(new_n523), .A3(new_n303), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT82), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT82), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n308), .A2(new_n526), .A3(new_n523), .A4(new_n303), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n525), .B(new_n527), .C1(new_n316), .C2(new_n523), .ZN(new_n528));
  OR2_X1    g342(.A1(new_n528), .A2(G146), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n324), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT83), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n189), .A2(new_n190), .A3(G214), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n533), .B(G143), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n534), .B(G131), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n529), .A2(new_n324), .A3(KEYINPUT83), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n532), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  XNOR2_X1  g352(.A(G113), .B(G122), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(new_n360), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(KEYINPUT18), .A2(G131), .ZN(new_n542));
  XOR2_X1   g356(.A(new_n534), .B(new_n542), .Z(new_n543));
  NOR2_X1   g357(.A1(new_n316), .A2(new_n233), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n543), .B1(new_n329), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n538), .A2(new_n541), .A3(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(G475), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT17), .ZN(new_n548));
  OR3_X1    g362(.A1(new_n534), .A2(new_n548), .A3(new_n228), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n549), .B1(new_n536), .B2(KEYINPUT17), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n545), .B1(new_n550), .B2(new_n325), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n540), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n546), .A2(new_n547), .A3(new_n281), .A4(new_n552), .ZN(new_n553));
  OR2_X1    g367(.A1(new_n553), .A2(KEYINPUT20), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(KEYINPUT20), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OR2_X1    g370(.A1(new_n540), .A2(KEYINPUT84), .ZN(new_n557));
  AOI21_X1  g371(.A(G902), .B1(new_n551), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n558), .B1(new_n557), .B2(new_n551), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(G475), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(G952), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n562), .A2(KEYINPUT93), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n562), .A2(KEYINPUT93), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n190), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n565), .B1(G234), .B2(G237), .ZN(new_n566));
  XOR2_X1   g380(.A(KEYINPUT21), .B(G898), .Z(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  AOI211_X1 g382(.A(new_n281), .B(new_n190), .C1(G234), .C2(G237), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n566), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NOR3_X1   g384(.A1(new_n522), .A2(new_n561), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n354), .A2(KEYINPUT76), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n355), .A2(new_n458), .A3(new_n571), .A4(new_n572), .ZN(new_n573));
  XOR2_X1   g387(.A(KEYINPUT94), .B(G101), .Z(new_n574));
  XNOR2_X1  g388(.A(new_n573), .B(new_n574), .ZN(G3));
  AND3_X1   g389(.A1(new_n273), .A2(new_n274), .A3(new_n278), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n282), .A2(new_n281), .ZN(new_n577));
  NAND2_X1  g391(.A1(KEYINPUT95), .A2(G472), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NOR3_X1   g393(.A1(new_n576), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n578), .B1(new_n286), .B2(new_n279), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT96), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n582), .A2(new_n583), .A3(new_n353), .A4(new_n416), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n579), .B1(new_n576), .B2(new_n577), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n286), .A2(new_n279), .A3(new_n578), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(new_n416), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(KEYINPUT25), .B1(new_n347), .B2(new_n281), .ZN(new_n588));
  NOR4_X1   g402(.A1(new_n344), .A2(new_n346), .A3(new_n342), .A4(G902), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n351), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n347), .A2(new_n352), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(KEYINPUT96), .B1(new_n587), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n584), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(KEYINPUT97), .ZN(new_n595));
  AOI21_X1  g409(.A(KEYINPUT92), .B1(new_n516), .B2(new_n281), .ZN(new_n596));
  NOR4_X1   g410(.A1(new_n514), .A2(new_n515), .A3(new_n512), .A4(G902), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n518), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT98), .ZN(new_n599));
  NAND2_X1  g413(.A1(G478), .A2(G902), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n504), .A2(KEYINPUT33), .A3(new_n510), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT33), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n602), .B1(new_n514), .B2(new_n515), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n601), .A2(new_n603), .A3(G478), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n598), .A2(new_n599), .A3(new_n600), .A4(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(G478), .B1(new_n513), .B2(new_n517), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n604), .A2(new_n600), .ZN(new_n607));
  OAI21_X1  g421(.A(KEYINPUT98), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  AOI22_X1  g423(.A1(new_n554), .A2(new_n555), .B1(G475), .B2(new_n559), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n457), .A2(new_n570), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n595), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT34), .B(G104), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G6));
  NAND3_X1  g430(.A1(new_n612), .A2(new_n522), .A3(new_n610), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n595), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(KEYINPUT99), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT35), .B(G107), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G9));
  NOR2_X1   g435(.A1(new_n338), .A2(KEYINPUT36), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n334), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n352), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n590), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n571), .A2(new_n458), .A3(new_n582), .A4(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT37), .B(G110), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT100), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n626), .B(new_n628), .ZN(G12));
  NAND2_X1  g443(.A1(new_n288), .A2(new_n625), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n630), .A2(new_n457), .A3(new_n417), .ZN(new_n631));
  INV_X1    g445(.A(new_n522), .ZN(new_n632));
  INV_X1    g446(.A(new_n566), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT101), .B(G900), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n569), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n632), .A2(new_n561), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n631), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G128), .ZN(G30));
  XNOR2_X1  g454(.A(KEYINPUT104), .B(KEYINPUT39), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n636), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n416), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT105), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT40), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n632), .A2(new_n610), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT103), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n455), .B(new_n648), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n285), .A2(new_n287), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n253), .A2(new_n255), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n651), .A2(new_n194), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n275), .A2(new_n254), .A3(new_n194), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n281), .ZN(new_n654));
  OAI21_X1  g468(.A(G472), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  AOI211_X1 g469(.A(new_n625), .B(new_n649), .C1(new_n650), .C2(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n645), .A2(new_n456), .A3(new_n646), .A4(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G143), .ZN(G45));
  NAND4_X1  g472(.A1(new_n605), .A2(new_n608), .A3(new_n561), .A4(new_n636), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n631), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G146), .ZN(G48));
  NOR4_X1   g476(.A1(new_n609), .A2(new_n457), .A3(new_n610), .A4(new_n570), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n411), .B(G469), .ZN(new_n664));
  INV_X1    g478(.A(new_n359), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n288), .A2(new_n353), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT41), .B(G113), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G15));
  INV_X1    g484(.A(new_n617), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n667), .A2(KEYINPUT106), .A3(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT106), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n288), .A2(new_n353), .A3(new_n666), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n673), .B1(new_n674), .B2(new_n617), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G116), .ZN(G18));
  INV_X1    g491(.A(new_n630), .ZN(new_n678));
  INV_X1    g492(.A(new_n666), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n679), .A2(new_n457), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n678), .A2(new_n571), .A3(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT107), .B(G119), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G21));
  NAND2_X1  g497(.A1(new_n283), .A2(KEYINPUT108), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n286), .A2(new_n685), .A3(new_n280), .A4(new_n279), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g501(.A(G472), .B1(new_n576), .B2(new_n577), .ZN(new_n688));
  AND3_X1   g502(.A1(new_n687), .A2(new_n353), .A3(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n689), .A2(new_n612), .A3(new_n646), .A4(new_n666), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G122), .ZN(G24));
  NAND4_X1  g505(.A1(new_n625), .A2(new_n688), .A3(new_n684), .A4(new_n686), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(KEYINPUT109), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT109), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n687), .A2(new_n694), .A3(new_n625), .A4(new_n688), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT110), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n659), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n659), .A2(new_n697), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n696), .B(new_n680), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G125), .ZN(G27));
  NAND2_X1  g515(.A1(new_n660), .A2(KEYINPUT110), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n659), .A2(new_n697), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n456), .ZN(new_n705));
  OAI21_X1  g519(.A(KEYINPUT111), .B1(new_n455), .B2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT111), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n453), .A2(new_n707), .A3(new_n456), .A4(new_n454), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n416), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n354), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n704), .A2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT42), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n704), .A2(KEYINPUT42), .A3(new_n712), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G131), .ZN(G33));
  NAND2_X1  g532(.A1(new_n712), .A2(new_n638), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G134), .ZN(G36));
  NAND3_X1  g534(.A1(new_n605), .A2(new_n608), .A3(new_n610), .ZN(new_n721));
  NAND2_X1  g535(.A1(KEYINPUT112), .A2(KEYINPUT43), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g537(.A(KEYINPUT112), .B(KEYINPUT43), .Z(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n605), .A2(new_n608), .A3(new_n610), .A4(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n582), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n727), .A2(KEYINPUT44), .A3(new_n728), .A4(new_n625), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT113), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n582), .B1(new_n723), .B2(new_n726), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT113), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n731), .A2(new_n732), .A3(KEYINPUT44), .A4(new_n625), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT114), .B1(new_n734), .B2(new_n710), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT114), .ZN(new_n736));
  AOI211_X1 g550(.A(new_n736), .B(new_n709), .C1(new_n730), .C2(new_n733), .ZN(new_n737));
  AOI21_X1  g551(.A(KEYINPUT44), .B1(new_n731), .B2(new_n625), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n735), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n390), .B1(new_n398), .B2(new_n389), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n741), .A2(KEYINPUT45), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(KEYINPUT45), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(G469), .A3(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n744), .A2(KEYINPUT46), .A3(new_n415), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n411), .A2(new_n412), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(KEYINPUT46), .B1(new_n744), .B2(new_n415), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n665), .B(new_n642), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n739), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G137), .ZN(G39));
  OAI21_X1  g566(.A(new_n665), .B1(new_n747), .B2(new_n748), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT47), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT47), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n755), .B(new_n665), .C1(new_n747), .C2(new_n748), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n288), .A2(new_n709), .A3(new_n353), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n754), .A2(new_n660), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G140), .ZN(G42));
  NOR3_X1   g573(.A1(new_n592), .A2(new_n705), .A3(new_n359), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(KEYINPUT115), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n650), .A2(new_n655), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n721), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n664), .B(KEYINPUT49), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n763), .A2(new_n649), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  AOI22_X1  g580(.A1(new_n702), .A2(new_n703), .B1(new_n695), .B2(new_n693), .ZN(new_n767));
  NOR4_X1   g581(.A1(new_n630), .A2(new_n561), .A3(new_n522), .A4(new_n637), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n416), .B(new_n710), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n584), .A2(new_n593), .A3(new_n671), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n626), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT116), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n770), .A2(new_n626), .A3(KEYINPUT116), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n773), .A2(new_n573), .A3(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n354), .ZN(new_n776));
  AOI22_X1  g590(.A1(new_n776), .A2(new_n666), .B1(new_n584), .B2(new_n593), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n681), .B1(new_n777), .B2(new_n613), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n672), .A2(new_n675), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n769), .A2(new_n775), .A3(new_n780), .A4(new_n690), .ZN(new_n781));
  INV_X1    g595(.A(new_n716), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT42), .B1(new_n704), .B2(new_n712), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n719), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n631), .B1(new_n660), .B2(new_n638), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n700), .A2(new_n786), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n632), .A2(new_n457), .A3(new_n610), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n625), .A2(new_n637), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n788), .A2(new_n762), .A3(new_n416), .A4(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n787), .A2(KEYINPUT117), .A3(KEYINPUT52), .A4(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n700), .A2(new_n786), .A3(new_n790), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n700), .A2(KEYINPUT52), .A3(new_n786), .A4(new_n790), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n791), .A2(new_n794), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n785), .A2(KEYINPUT53), .A3(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n800));
  INV_X1    g614(.A(new_n719), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n801), .B1(new_n715), .B2(new_n716), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n773), .A2(new_n573), .A3(new_n690), .A4(new_n774), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n676), .B(new_n681), .C1(new_n613), .C2(new_n777), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n802), .A2(new_n805), .A3(new_n769), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n794), .A2(new_n795), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n800), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n799), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n785), .A2(new_n798), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n800), .ZN(new_n813));
  AND4_X1   g627(.A1(new_n690), .A2(new_n769), .A3(new_n775), .A4(new_n780), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n814), .A2(new_n807), .A3(KEYINPUT53), .A4(new_n802), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT118), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n785), .A2(new_n817), .A3(KEYINPUT53), .A4(new_n807), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n813), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n811), .B1(new_n819), .B2(KEYINPUT54), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n666), .A2(new_n706), .A3(new_n708), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT119), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n710), .A2(KEYINPUT119), .A3(new_n666), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(new_n566), .A3(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(new_n776), .A3(new_n727), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT48), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n727), .A2(new_n566), .A3(new_n689), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n754), .A2(new_n756), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n664), .A2(new_n359), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n709), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n826), .A2(new_n727), .A3(new_n696), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n650), .A2(new_n353), .A3(new_n655), .ZN(new_n836));
  OAI21_X1  g650(.A(KEYINPUT120), .B1(new_n825), .B2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n836), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n633), .B1(new_n821), .B2(new_n822), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT120), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n838), .A2(new_n839), .A3(new_n840), .A4(new_n824), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n837), .A2(new_n610), .A3(new_n609), .A4(new_n841), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n842), .A2(KEYINPUT121), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(KEYINPUT121), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n835), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n829), .A2(new_n666), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n846), .A2(KEYINPUT50), .A3(new_n705), .A4(new_n649), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT50), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n829), .A2(new_n649), .A3(new_n666), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n848), .B1(new_n849), .B2(new_n456), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n845), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT51), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n565), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n837), .A2(new_n611), .A3(new_n841), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n845), .A2(new_n851), .A3(KEYINPUT51), .ZN(new_n856));
  AND4_X1   g670(.A1(new_n828), .A2(new_n854), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n829), .A2(new_n680), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n820), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(G952), .A2(G953), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n766), .B1(new_n859), .B2(new_n860), .ZN(G75));
  AOI21_X1  g675(.A(new_n281), .B1(new_n799), .B2(new_n809), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(G210), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT56), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n429), .B1(new_n435), .B2(new_n436), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(new_n433), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(KEYINPUT55), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n868), .B1(KEYINPUT122), .B2(new_n864), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n863), .A2(new_n864), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n869), .B1(new_n863), .B2(new_n864), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n190), .A2(G952), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(G51));
  NAND2_X1  g687(.A1(new_n415), .A2(KEYINPUT57), .ZN(new_n874));
  OR2_X1    g688(.A1(new_n415), .A2(KEYINPUT57), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n810), .B1(new_n799), .B2(new_n809), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n874), .B(new_n875), .C1(new_n811), .C2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n408), .A2(new_n410), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n744), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n862), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n872), .B1(new_n879), .B2(new_n881), .ZN(G54));
  AND3_X1   g696(.A1(new_n862), .A2(KEYINPUT58), .A3(G475), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n546), .A2(new_n552), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n883), .A2(new_n884), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n885), .A2(new_n886), .A3(new_n872), .ZN(G60));
  AND2_X1   g701(.A1(new_n601), .A2(new_n603), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n600), .B(KEYINPUT59), .Z(new_n889));
  OAI21_X1  g703(.A(new_n888), .B1(new_n820), .B2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT123), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n888), .A2(new_n889), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n799), .A2(new_n809), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(KEYINPUT54), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n799), .A2(new_n809), .A3(new_n810), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n893), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n891), .B1(new_n897), .B2(new_n872), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n892), .B1(new_n811), .B2(new_n876), .ZN(new_n899));
  INV_X1    g713(.A(new_n872), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n899), .A2(KEYINPUT123), .A3(new_n900), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n890), .A2(new_n898), .A3(new_n901), .ZN(G63));
  NAND2_X1  g716(.A1(G217), .A2(G902), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT60), .Z(new_n904));
  NAND3_X1  g718(.A1(new_n894), .A2(new_n623), .A3(new_n904), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n905), .A2(new_n900), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n894), .A2(new_n904), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n907), .B1(new_n346), .B2(new_n344), .ZN(new_n908));
  XNOR2_X1  g722(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n906), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n909), .B1(new_n906), .B2(new_n908), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n910), .A2(new_n911), .ZN(G66));
  INV_X1    g726(.A(G224), .ZN(new_n913));
  OAI21_X1  g727(.A(G953), .B1(new_n568), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n914), .B1(new_n805), .B2(G953), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n915), .B(KEYINPUT125), .Z(new_n916));
  OAI21_X1  g730(.A(new_n865), .B1(G898), .B2(new_n190), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n916), .B(new_n917), .ZN(G69));
  AND2_X1   g732(.A1(new_n776), .A2(new_n788), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n750), .B1(new_n739), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n247), .A2(new_n252), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(new_n528), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n802), .A2(new_n758), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n920), .A2(new_n787), .A3(new_n923), .A4(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n787), .A2(new_n657), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT62), .Z(new_n927));
  NOR2_X1   g741(.A1(new_n632), .A2(new_n561), .ZN(new_n928));
  OR2_X1    g742(.A1(new_n611), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n709), .A2(new_n643), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n929), .A2(new_n572), .A3(new_n355), .A4(new_n930), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n931), .A2(new_n758), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n751), .A2(new_n927), .A3(new_n932), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n925), .B(new_n190), .C1(new_n933), .C2(new_n923), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n190), .B1(new_n923), .B2(G227), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n935), .B(G900), .C1(G227), .C2(new_n923), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n934), .A2(new_n936), .ZN(G72));
  NAND4_X1  g751(.A1(new_n751), .A2(new_n805), .A3(new_n927), .A4(new_n932), .ZN(new_n938));
  NAND2_X1  g752(.A1(G472), .A2(G902), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT63), .Z(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT126), .Z(new_n941));
  NAND2_X1  g755(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n652), .ZN(new_n943));
  INV_X1    g757(.A(new_n652), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n651), .A2(new_n194), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n819), .A2(new_n944), .A3(new_n940), .A4(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n943), .A2(new_n900), .A3(new_n946), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n920), .A2(new_n787), .A3(new_n805), .A4(new_n924), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n948), .A2(KEYINPUT127), .A3(new_n941), .ZN(new_n949));
  AOI21_X1  g763(.A(KEYINPUT127), .B1(new_n948), .B2(new_n941), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n945), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n947), .B1(new_n951), .B2(new_n952), .ZN(G57));
endmodule


