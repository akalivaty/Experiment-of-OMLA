

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765;

  XNOR2_X1 U376 ( .A(n623), .B(n622), .ZN(n624) );
  NOR2_X1 U377 ( .A1(n553), .A2(n556), .ZN(n534) );
  NOR2_X1 U378 ( .A1(n696), .A2(n704), .ZN(n521) );
  XNOR2_X1 U379 ( .A(n355), .B(n452), .ZN(n623) );
  XNOR2_X1 U380 ( .A(G143), .B(G113), .ZN(n497) );
  NOR2_X2 U381 ( .A1(n584), .A2(KEYINPUT44), .ZN(n582) );
  XNOR2_X1 U382 ( .A(n354), .B(n549), .ZN(n405) );
  NAND2_X1 U383 ( .A1(n765), .A2(n764), .ZN(n354) );
  NOR2_X2 U384 ( .A1(n669), .A2(n552), .ZN(n543) );
  XNOR2_X1 U385 ( .A(n460), .B(n463), .ZN(n355) );
  XNOR2_X2 U386 ( .A(n752), .B(KEYINPUT77), .ZN(n609) );
  XNOR2_X2 U387 ( .A(n444), .B(KEYINPUT3), .ZN(n402) );
  XNOR2_X2 U388 ( .A(n471), .B(n470), .ZN(n740) );
  XNOR2_X2 U389 ( .A(n402), .B(n401), .ZN(n471) );
  XNOR2_X2 U390 ( .A(n356), .B(n376), .ZN(n598) );
  NAND2_X2 U391 ( .A1(n566), .A2(n418), .ZN(n356) );
  XNOR2_X2 U392 ( .A(n503), .B(n502), .ZN(n632) );
  XNOR2_X2 U393 ( .A(n476), .B(n395), .ZN(n492) );
  AND2_X1 U394 ( .A1(n573), .A2(n687), .ZN(n691) );
  AND2_X2 U395 ( .A1(n412), .A2(n407), .ZN(n400) );
  INV_X2 U396 ( .A(n654), .ZN(n357) );
  INV_X1 U397 ( .A(G146), .ZN(n449) );
  INV_X4 U398 ( .A(G953), .ZN(n753) );
  XNOR2_X1 U399 ( .A(n415), .B(KEYINPUT39), .ZN(n552) );
  AND2_X1 U400 ( .A1(n367), .A2(n539), .ZN(n415) );
  XNOR2_X1 U401 ( .A(n463), .B(n462), .ZN(n478) );
  XNOR2_X1 U402 ( .A(n749), .B(n449), .ZN(n460) );
  XNOR2_X1 U403 ( .A(n496), .B(G134), .ZN(n749) );
  XNOR2_X1 U404 ( .A(n748), .B(n450), .ZN(n463) );
  XNOR2_X1 U405 ( .A(n505), .B(n380), .ZN(n748) );
  INV_X2 U406 ( .A(G125), .ZN(n396) );
  INV_X1 U407 ( .A(n600), .ZN(n358) );
  XNOR2_X1 U408 ( .A(n468), .B(n467), .ZN(n538) );
  BUF_X1 U409 ( .A(n740), .Z(n359) );
  INV_X1 U410 ( .A(n596), .ZN(n360) );
  XNOR2_X2 U411 ( .A(n392), .B(n364), .ZN(n566) );
  XNOR2_X1 U412 ( .A(n382), .B(KEYINPUT80), .ZN(n381) );
  OR2_X2 U413 ( .A1(n761), .A2(n361), .ZN(n382) );
  NAND2_X1 U414 ( .A1(n411), .A2(n410), .ZN(n409) );
  INV_X1 U415 ( .A(n613), .ZN(n411) );
  INV_X1 U416 ( .A(KEYINPUT67), .ZN(n410) );
  INV_X1 U417 ( .A(KEYINPUT46), .ZN(n549) );
  INV_X1 U418 ( .A(KEYINPUT66), .ZN(n397) );
  NOR2_X1 U419 ( .A1(n705), .A2(n600), .ZN(n539) );
  NOR2_X1 U420 ( .A1(n362), .A2(n541), .ZN(n367) );
  INV_X1 U421 ( .A(KEYINPUT22), .ZN(n390) );
  XNOR2_X1 U422 ( .A(n521), .B(n387), .ZN(n541) );
  INV_X1 U423 ( .A(KEYINPUT30), .ZN(n387) );
  NOR2_X1 U424 ( .A1(n531), .A2(n696), .ZN(n456) );
  BUF_X1 U425 ( .A(n658), .Z(n661) );
  NOR2_X1 U426 ( .A1(n753), .A2(G952), .ZN(n666) );
  XNOR2_X1 U427 ( .A(KEYINPUT5), .B(KEYINPUT96), .ZN(n445) );
  XNOR2_X1 U428 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n380) );
  NOR2_X1 U429 ( .A1(G953), .A2(G237), .ZN(n491) );
  INV_X1 U430 ( .A(KEYINPUT10), .ZN(n395) );
  XNOR2_X1 U431 ( .A(G119), .B(G116), .ZN(n401) );
  NAND2_X1 U432 ( .A1(n365), .A2(n408), .ZN(n407) );
  NAND2_X1 U433 ( .A1(n409), .A2(n618), .ZN(n408) );
  NAND2_X1 U434 ( .A1(n406), .A2(n366), .ZN(n399) );
  INV_X1 U435 ( .A(KEYINPUT0), .ZN(n376) );
  XNOR2_X1 U436 ( .A(G110), .B(G107), .ZN(n461) );
  XNOR2_X1 U437 ( .A(G128), .B(G110), .ZN(n423) );
  XNOR2_X1 U438 ( .A(G134), .B(G116), .ZN(n508) );
  INV_X4 U439 ( .A(KEYINPUT71), .ZN(n369) );
  XNOR2_X1 U440 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n473) );
  NAND2_X1 U441 ( .A1(n725), .A2(KEYINPUT2), .ZN(n727) );
  INV_X1 U442 ( .A(KEYINPUT100), .ZN(n517) );
  NAND2_X1 U443 ( .A1(n394), .A2(n589), .ZN(n393) );
  XNOR2_X1 U444 ( .A(n593), .B(KEYINPUT103), .ZN(n394) );
  BUF_X1 U445 ( .A(n696), .Z(n370) );
  INV_X1 U446 ( .A(n692), .ZN(n388) );
  XNOR2_X1 U447 ( .A(n464), .B(n478), .ZN(n663) );
  XNOR2_X1 U448 ( .A(n460), .B(n459), .ZN(n464) );
  AND2_X1 U449 ( .A1(n524), .A2(n384), .ZN(n526) );
  NOR2_X1 U450 ( .A1(n541), .A2(n385), .ZN(n384) );
  NOR2_X1 U451 ( .A1(n546), .A2(n560), .ZN(n682) );
  XNOR2_X1 U452 ( .A(n655), .B(n372), .ZN(n657) );
  XNOR2_X1 U453 ( .A(n374), .B(n373), .ZN(n660) );
  INV_X1 U454 ( .A(n659), .ZN(n373) );
  INV_X1 U455 ( .A(n540), .ZN(n386) );
  XOR2_X1 U456 ( .A(n528), .B(KEYINPUT82), .Z(n361) );
  NAND2_X1 U457 ( .A1(n691), .A2(n386), .ZN(n362) );
  AND2_X1 U458 ( .A1(n692), .A2(n575), .ZN(n363) );
  XOR2_X1 U459 ( .A(n488), .B(KEYINPUT19), .Z(n364) );
  OR2_X1 U460 ( .A1(n618), .A2(KEYINPUT67), .ZN(n365) );
  AND2_X1 U461 ( .A1(n618), .A2(n410), .ZN(n366) );
  XNOR2_X1 U462 ( .A(n427), .B(n751), .ZN(n656) );
  NAND2_X1 U463 ( .A1(n400), .A2(n399), .ZN(n398) );
  NOR2_X1 U464 ( .A1(n383), .A2(n381), .ZN(n404) );
  XNOR2_X2 U465 ( .A(n368), .B(n397), .ZN(n658) );
  NAND2_X1 U466 ( .A1(n398), .A2(n727), .ZN(n368) );
  NOR2_X1 U467 ( .A1(n705), .A2(n704), .ZN(n710) );
  XNOR2_X2 U468 ( .A(n369), .B(G131), .ZN(n496) );
  NAND2_X1 U469 ( .A1(n529), .A2(n762), .ZN(n383) );
  INV_X1 U470 ( .A(n656), .ZN(n372) );
  NAND2_X1 U471 ( .A1(n661), .A2(G478), .ZN(n374) );
  INV_X1 U472 ( .A(n598), .ZN(n596) );
  XNOR2_X2 U473 ( .A(n375), .B(n390), .ZN(n389) );
  NAND2_X1 U474 ( .A1(n598), .A2(n567), .ZN(n375) );
  XNOR2_X2 U475 ( .A(n377), .B(KEYINPUT35), .ZN(n654) );
  NAND2_X1 U476 ( .A1(n378), .A2(n522), .ZN(n377) );
  XNOR2_X1 U477 ( .A(n379), .B(KEYINPUT34), .ZN(n378) );
  NOR2_X2 U478 ( .A1(n721), .A2(n596), .ZN(n379) );
  XNOR2_X2 U479 ( .A(G143), .B(G128), .ZN(n505) );
  NAND2_X1 U480 ( .A1(n358), .A2(n386), .ZN(n385) );
  NAND2_X2 U481 ( .A1(n389), .A2(n388), .ZN(n590) );
  NAND2_X1 U482 ( .A1(n389), .A2(n363), .ZN(n577) );
  NAND2_X1 U483 ( .A1(n537), .A2(n487), .ZN(n392) );
  NAND2_X1 U484 ( .A1(n357), .A2(KEYINPUT87), .ZN(n581) );
  NAND2_X1 U485 ( .A1(n357), .A2(n583), .ZN(n585) );
  XNOR2_X2 U486 ( .A(n393), .B(n579), .ZN(n721) );
  XNOR2_X2 U487 ( .A(n396), .B(G146), .ZN(n476) );
  INV_X1 U488 ( .A(n566), .ZN(n560) );
  XNOR2_X2 U489 ( .A(n483), .B(n482), .ZN(n537) );
  AND2_X1 U490 ( .A1(n619), .A2(n414), .ZN(n725) );
  NAND2_X2 U491 ( .A1(n559), .A2(n558), .ZN(n752) );
  XNOR2_X1 U492 ( .A(n538), .B(KEYINPUT1), .ZN(n578) );
  XNOR2_X1 U493 ( .A(n403), .B(n550), .ZN(n559) );
  NAND2_X1 U494 ( .A1(n405), .A2(n404), .ZN(n403) );
  INV_X1 U495 ( .A(n614), .ZN(n406) );
  NAND2_X1 U496 ( .A1(n614), .A2(n413), .ZN(n412) );
  AND2_X1 U497 ( .A1(n613), .A2(KEYINPUT67), .ZN(n413) );
  INV_X1 U498 ( .A(n619), .ZN(n733) );
  INV_X1 U499 ( .A(n752), .ZN(n414) );
  XNOR2_X1 U500 ( .A(n537), .B(KEYINPUT38), .ZN(n705) );
  XNOR2_X1 U501 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U502 ( .A(n498), .B(n497), .Z(n416) );
  XNOR2_X1 U503 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n417) );
  XOR2_X1 U504 ( .A(n565), .B(KEYINPUT93), .Z(n418) );
  XNOR2_X1 U505 ( .A(n445), .B(G137), .ZN(n447) );
  XNOR2_X1 U506 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U507 ( .A(n499), .B(n416), .ZN(n500) );
  BUF_X1 U508 ( .A(n578), .Z(n692) );
  INV_X1 U509 ( .A(KEYINPUT63), .ZN(n627) );
  XOR2_X1 U510 ( .A(KEYINPUT48), .B(KEYINPUT72), .Z(n550) );
  XNOR2_X1 U511 ( .A(G140), .B(G137), .ZN(n458) );
  XOR2_X1 U512 ( .A(n492), .B(n458), .Z(n751) );
  XOR2_X1 U513 ( .A(KEYINPUT84), .B(KEYINPUT8), .Z(n420) );
  NAND2_X1 U514 ( .A1(G234), .A2(n753), .ZN(n419) );
  XNOR2_X1 U515 ( .A(n420), .B(n419), .ZN(n504) );
  NAND2_X1 U516 ( .A1(G221), .A2(n504), .ZN(n422) );
  XNOR2_X1 U517 ( .A(G119), .B(KEYINPUT23), .ZN(n421) );
  XNOR2_X1 U518 ( .A(n422), .B(n421), .ZN(n426) );
  XOR2_X1 U519 ( .A(KEYINPUT83), .B(KEYINPUT24), .Z(n424) );
  XNOR2_X1 U520 ( .A(n424), .B(n423), .ZN(n425) );
  INV_X1 U521 ( .A(G902), .ZN(n514) );
  NAND2_X1 U522 ( .A1(n656), .A2(n514), .ZN(n434) );
  XOR2_X1 U523 ( .A(KEYINPUT94), .B(KEYINPUT25), .Z(n430) );
  XNOR2_X1 U524 ( .A(G902), .B(KEYINPUT15), .ZN(n480) );
  NAND2_X1 U525 ( .A1(n480), .A2(G234), .ZN(n428) );
  XNOR2_X1 U526 ( .A(n428), .B(KEYINPUT20), .ZN(n440) );
  NAND2_X1 U527 ( .A1(G217), .A2(n440), .ZN(n429) );
  XNOR2_X1 U528 ( .A(n430), .B(n429), .ZN(n432) );
  INV_X1 U529 ( .A(KEYINPUT95), .ZN(n431) );
  XNOR2_X1 U530 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X2 U531 ( .A(n434), .B(n433), .ZN(n573) );
  NAND2_X1 U532 ( .A1(G234), .A2(G237), .ZN(n435) );
  XNOR2_X1 U533 ( .A(n435), .B(KEYINPUT14), .ZN(n436) );
  NAND2_X1 U534 ( .A1(G952), .A2(n436), .ZN(n719) );
  NOR2_X1 U535 ( .A1(G953), .A2(n719), .ZN(n564) );
  NAND2_X1 U536 ( .A1(G902), .A2(n436), .ZN(n561) );
  OR2_X1 U537 ( .A1(n753), .A2(n561), .ZN(n437) );
  XNOR2_X1 U538 ( .A(KEYINPUT104), .B(n437), .ZN(n438) );
  NOR2_X1 U539 ( .A1(G900), .A2(n438), .ZN(n439) );
  NOR2_X1 U540 ( .A1(n564), .A2(n439), .ZN(n540) );
  NOR2_X1 U541 ( .A1(n573), .A2(n540), .ZN(n443) );
  NAND2_X1 U542 ( .A1(n440), .A2(G221), .ZN(n442) );
  INV_X1 U543 ( .A(KEYINPUT21), .ZN(n441) );
  XNOR2_X1 U544 ( .A(n442), .B(n441), .ZN(n687) );
  NAND2_X1 U545 ( .A1(n443), .A2(n687), .ZN(n531) );
  XNOR2_X2 U546 ( .A(G113), .B(KEYINPUT75), .ZN(n444) );
  NAND2_X1 U547 ( .A1(n491), .A2(G210), .ZN(n446) );
  XNOR2_X1 U548 ( .A(n471), .B(n448), .ZN(n452) );
  XNOR2_X1 U549 ( .A(KEYINPUT70), .B(G101), .ZN(n450) );
  NAND2_X1 U550 ( .A1(n623), .A2(n514), .ZN(n454) );
  INV_X1 U551 ( .A(G472), .ZN(n453) );
  XNOR2_X2 U552 ( .A(n454), .B(n453), .ZN(n696) );
  XNOR2_X1 U553 ( .A(KEYINPUT106), .B(KEYINPUT28), .ZN(n455) );
  XNOR2_X1 U554 ( .A(n456), .B(n455), .ZN(n469) );
  NAND2_X1 U555 ( .A1(n753), .A2(G227), .ZN(n457) );
  XNOR2_X1 U556 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U557 ( .A(n461), .B(G104), .ZN(n741) );
  XNOR2_X1 U558 ( .A(n741), .B(KEYINPUT76), .ZN(n462) );
  NAND2_X1 U559 ( .A1(n663), .A2(n514), .ZN(n468) );
  XNOR2_X1 U560 ( .A(KEYINPUT74), .B(G469), .ZN(n466) );
  INV_X1 U561 ( .A(KEYINPUT73), .ZN(n465) );
  XNOR2_X1 U562 ( .A(n466), .B(n465), .ZN(n467) );
  NAND2_X1 U563 ( .A1(n469), .A2(n358), .ZN(n546) );
  XNOR2_X1 U564 ( .A(KEYINPUT16), .B(G122), .ZN(n470) );
  NAND2_X1 U565 ( .A1(n753), .A2(G224), .ZN(n472) );
  XNOR2_X1 U566 ( .A(n472), .B(KEYINPUT89), .ZN(n474) );
  XNOR2_X1 U567 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U568 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U569 ( .A(n740), .B(n477), .ZN(n479) );
  XNOR2_X1 U570 ( .A(n479), .B(n478), .ZN(n647) );
  INV_X1 U571 ( .A(n480), .ZN(n616) );
  OR2_X2 U572 ( .A1(n647), .A2(n616), .ZN(n483) );
  INV_X1 U573 ( .A(G237), .ZN(n481) );
  NAND2_X1 U574 ( .A1(n514), .A2(n481), .ZN(n484) );
  AND2_X1 U575 ( .A1(n484), .A2(G210), .ZN(n482) );
  NAND2_X1 U576 ( .A1(n484), .A2(G214), .ZN(n486) );
  INV_X1 U577 ( .A(KEYINPUT90), .ZN(n485) );
  XNOR2_X1 U578 ( .A(n486), .B(n485), .ZN(n704) );
  INV_X1 U579 ( .A(n704), .ZN(n487) );
  INV_X1 U580 ( .A(KEYINPUT78), .ZN(n488) );
  XOR2_X1 U581 ( .A(KEYINPUT47), .B(n682), .Z(n520) );
  XNOR2_X1 U582 ( .A(KEYINPUT13), .B(G475), .ZN(n503) );
  XOR2_X1 U583 ( .A(KEYINPUT97), .B(KEYINPUT12), .Z(n490) );
  XNOR2_X1 U584 ( .A(G122), .B(KEYINPUT11), .ZN(n489) );
  XNOR2_X1 U585 ( .A(n490), .B(n489), .ZN(n495) );
  NAND2_X1 U586 ( .A1(G214), .A2(n491), .ZN(n493) );
  XNOR2_X1 U587 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U588 ( .A(n495), .B(n494), .Z(n501) );
  XNOR2_X1 U589 ( .A(n496), .B(KEYINPUT98), .ZN(n499) );
  XOR2_X1 U590 ( .A(G104), .B(G140), .Z(n498) );
  XNOR2_X1 U591 ( .A(n501), .B(n500), .ZN(n642) );
  NOR2_X1 U592 ( .A1(G902), .A2(n642), .ZN(n502) );
  NAND2_X1 U593 ( .A1(G217), .A2(n504), .ZN(n507) );
  XNOR2_X1 U594 ( .A(n505), .B(KEYINPUT7), .ZN(n506) );
  XNOR2_X1 U595 ( .A(n507), .B(n506), .ZN(n513) );
  XOR2_X1 U596 ( .A(G122), .B(G107), .Z(n509) );
  XNOR2_X1 U597 ( .A(n509), .B(n508), .ZN(n511) );
  XOR2_X1 U598 ( .A(KEYINPUT9), .B(KEYINPUT99), .Z(n510) );
  XNOR2_X1 U599 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U600 ( .A(n513), .B(n512), .ZN(n659) );
  NAND2_X1 U601 ( .A1(n659), .A2(n514), .ZN(n516) );
  INV_X1 U602 ( .A(G478), .ZN(n515) );
  XNOR2_X1 U603 ( .A(n516), .B(n515), .ZN(n633) );
  NOR2_X1 U604 ( .A1(n632), .A2(n633), .ZN(n518) );
  XNOR2_X1 U605 ( .A(n518), .B(n517), .ZN(n551) );
  NAND2_X1 U606 ( .A1(n633), .A2(n632), .ZN(n669) );
  AND2_X1 U607 ( .A1(n551), .A2(n669), .ZN(n527) );
  NAND2_X1 U608 ( .A1(n682), .A2(n527), .ZN(n519) );
  NAND2_X1 U609 ( .A1(n520), .A2(n519), .ZN(n529) );
  INV_X1 U610 ( .A(n632), .ZN(n580) );
  NOR2_X1 U611 ( .A1(n633), .A2(n580), .ZN(n522) );
  NAND2_X1 U612 ( .A1(n522), .A2(n691), .ZN(n523) );
  INV_X1 U613 ( .A(n537), .ZN(n556) );
  NOR2_X1 U614 ( .A1(n523), .A2(n556), .ZN(n524) );
  INV_X1 U615 ( .A(KEYINPUT105), .ZN(n525) );
  XNOR2_X1 U616 ( .A(n526), .B(n525), .ZN(n761) );
  NAND2_X1 U617 ( .A1(KEYINPUT47), .A2(n527), .ZN(n528) );
  INV_X1 U618 ( .A(KEYINPUT6), .ZN(n530) );
  XNOR2_X1 U619 ( .A(n696), .B(n530), .ZN(n588) );
  NOR2_X1 U620 ( .A1(n531), .A2(n588), .ZN(n533) );
  NOR2_X1 U621 ( .A1(n704), .A2(n669), .ZN(n532) );
  NAND2_X1 U622 ( .A1(n533), .A2(n532), .ZN(n553) );
  XNOR2_X1 U623 ( .A(n534), .B(KEYINPUT36), .ZN(n535) );
  NAND2_X1 U624 ( .A1(n535), .A2(n692), .ZN(n536) );
  XNOR2_X1 U625 ( .A(n536), .B(KEYINPUT110), .ZN(n762) );
  INV_X1 U626 ( .A(n538), .ZN(n600) );
  XNOR2_X1 U627 ( .A(KEYINPUT107), .B(KEYINPUT40), .ZN(n542) );
  XNOR2_X1 U628 ( .A(n543), .B(n542), .ZN(n765) );
  XOR2_X1 U629 ( .A(KEYINPUT108), .B(KEYINPUT41), .Z(n545) );
  AND2_X1 U630 ( .A1(n633), .A2(n580), .ZN(n707) );
  NAND2_X1 U631 ( .A1(n707), .A2(n710), .ZN(n544) );
  XNOR2_X1 U632 ( .A(n545), .B(n544), .ZN(n720) );
  NOR2_X1 U633 ( .A1(n720), .A2(n546), .ZN(n548) );
  XNOR2_X1 U634 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n547) );
  XNOR2_X1 U635 ( .A(n548), .B(n547), .ZN(n764) );
  OR2_X1 U636 ( .A1(n552), .A2(n551), .ZN(n684) );
  NOR2_X1 U637 ( .A1(n553), .A2(n692), .ZN(n555) );
  INV_X1 U638 ( .A(KEYINPUT43), .ZN(n554) );
  XNOR2_X1 U639 ( .A(n555), .B(n554), .ZN(n557) );
  NAND2_X1 U640 ( .A1(n557), .A2(n556), .ZN(n629) );
  AND2_X1 U641 ( .A1(n684), .A2(n629), .ZN(n558) );
  XNOR2_X1 U642 ( .A(KEYINPUT91), .B(G898), .ZN(n736) );
  NAND2_X1 U643 ( .A1(G953), .A2(n736), .ZN(n743) );
  NOR2_X1 U644 ( .A1(n561), .A2(n743), .ZN(n562) );
  XNOR2_X1 U645 ( .A(n562), .B(KEYINPUT92), .ZN(n563) );
  OR2_X1 U646 ( .A1(n564), .A2(n563), .ZN(n565) );
  AND2_X1 U647 ( .A1(n707), .A2(n687), .ZN(n567) );
  INV_X1 U648 ( .A(KEYINPUT102), .ZN(n568) );
  XNOR2_X1 U649 ( .A(n590), .B(n568), .ZN(n571) );
  INV_X1 U650 ( .A(n573), .ZN(n569) );
  AND2_X1 U651 ( .A1(n569), .A2(n370), .ZN(n570) );
  NAND2_X1 U652 ( .A1(n571), .A2(n570), .ZN(n636) );
  INV_X1 U653 ( .A(KEYINPUT101), .ZN(n572) );
  XNOR2_X1 U654 ( .A(n573), .B(n572), .ZN(n688) );
  INV_X1 U655 ( .A(n688), .ZN(n574) );
  AND2_X1 U656 ( .A1(n574), .A2(n588), .ZN(n575) );
  XNOR2_X1 U657 ( .A(KEYINPUT68), .B(KEYINPUT32), .ZN(n576) );
  XNOR2_X1 U658 ( .A(n577), .B(n576), .ZN(n638) );
  AND2_X2 U659 ( .A1(n636), .A2(n638), .ZN(n584) );
  NAND2_X1 U660 ( .A1(n578), .A2(n691), .ZN(n593) );
  INV_X1 U661 ( .A(KEYINPUT33), .ZN(n579) );
  NAND2_X1 U662 ( .A1(n581), .A2(n582), .ZN(n587) );
  NOR2_X1 U663 ( .A1(KEYINPUT44), .A2(KEYINPUT87), .ZN(n583) );
  NAND2_X1 U664 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U665 ( .A1(n587), .A2(n586), .ZN(n607) );
  AND2_X1 U666 ( .A1(n654), .A2(KEYINPUT44), .ZN(n605) );
  INV_X1 U667 ( .A(n588), .ZN(n589) );
  NOR2_X1 U668 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U669 ( .A(n591), .B(KEYINPUT86), .ZN(n592) );
  NAND2_X1 U670 ( .A1(n592), .A2(n688), .ZN(n639) );
  INV_X1 U671 ( .A(n593), .ZN(n595) );
  INV_X1 U672 ( .A(n370), .ZN(n594) );
  NAND2_X1 U673 ( .A1(n595), .A2(n594), .ZN(n698) );
  NOR2_X1 U674 ( .A1(n596), .A2(n698), .ZN(n597) );
  XNOR2_X1 U675 ( .A(n597), .B(KEYINPUT31), .ZN(n634) );
  NAND2_X1 U676 ( .A1(n691), .A2(n370), .ZN(n599) );
  NOR2_X1 U677 ( .A1(n600), .A2(n599), .ZN(n601) );
  NAND2_X1 U678 ( .A1(n360), .A2(n601), .ZN(n668) );
  NAND2_X1 U679 ( .A1(n634), .A2(n668), .ZN(n602) );
  INV_X1 U680 ( .A(n527), .ZN(n709) );
  NAND2_X1 U681 ( .A1(n602), .A2(n709), .ZN(n603) );
  NAND2_X1 U682 ( .A1(n639), .A2(n603), .ZN(n604) );
  NOR2_X1 U683 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U684 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X2 U685 ( .A(n608), .B(n417), .ZN(n619) );
  NAND2_X1 U686 ( .A1(n609), .A2(n619), .ZN(n614) );
  INV_X1 U687 ( .A(KEYINPUT69), .ZN(n610) );
  NAND2_X1 U688 ( .A1(n610), .A2(KEYINPUT2), .ZN(n612) );
  NAND2_X1 U689 ( .A1(n616), .A2(KEYINPUT2), .ZN(n611) );
  NAND2_X1 U690 ( .A1(n611), .A2(KEYINPUT69), .ZN(n615) );
  AND2_X1 U691 ( .A1(n612), .A2(n615), .ZN(n613) );
  INV_X1 U692 ( .A(n615), .ZN(n617) );
  OR2_X1 U693 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U694 ( .A1(n658), .A2(G472), .ZN(n625) );
  XNOR2_X1 U695 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n621) );
  XNOR2_X1 U696 ( .A(KEYINPUT62), .B(KEYINPUT88), .ZN(n620) );
  XNOR2_X1 U697 ( .A(n621), .B(n620), .ZN(n622) );
  XNOR2_X1 U698 ( .A(n625), .B(n624), .ZN(n626) );
  NOR2_X2 U699 ( .A1(n626), .A2(n666), .ZN(n628) );
  XNOR2_X1 U700 ( .A(n628), .B(n627), .ZN(G57) );
  XNOR2_X1 U701 ( .A(n629), .B(G140), .ZN(G42) );
  XOR2_X1 U702 ( .A(G113), .B(KEYINPUT115), .Z(n631) );
  NOR2_X1 U703 ( .A1(n634), .A2(n669), .ZN(n630) );
  XOR2_X1 U704 ( .A(n631), .B(n630), .Z(G15) );
  OR2_X1 U705 ( .A1(n633), .A2(n632), .ZN(n671) );
  NOR2_X1 U706 ( .A1(n634), .A2(n671), .ZN(n635) );
  XOR2_X1 U707 ( .A(G116), .B(n635), .Z(G18) );
  BUF_X1 U708 ( .A(n636), .Z(n637) );
  XNOR2_X1 U709 ( .A(n637), .B(G110), .ZN(G12) );
  XNOR2_X1 U710 ( .A(n638), .B(G119), .ZN(G21) );
  XNOR2_X1 U711 ( .A(n639), .B(G101), .ZN(G3) );
  NAND2_X1 U712 ( .A1(n658), .A2(G475), .ZN(n644) );
  XNOR2_X1 U713 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n640) );
  XNOR2_X1 U714 ( .A(n640), .B(KEYINPUT59), .ZN(n641) );
  XNOR2_X1 U715 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U716 ( .A(n644), .B(n643), .ZN(n645) );
  NOR2_X2 U717 ( .A1(n645), .A2(n666), .ZN(n646) );
  XNOR2_X1 U718 ( .A(n646), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U719 ( .A1(n658), .A2(G210), .ZN(n651) );
  XNOR2_X1 U720 ( .A(KEYINPUT81), .B(KEYINPUT54), .ZN(n648) );
  XNOR2_X1 U721 ( .A(n648), .B(KEYINPUT55), .ZN(n649) );
  XNOR2_X1 U722 ( .A(n647), .B(n649), .ZN(n650) );
  XNOR2_X1 U723 ( .A(n651), .B(n650), .ZN(n652) );
  NOR2_X2 U724 ( .A1(n652), .A2(n666), .ZN(n653) );
  XNOR2_X1 U725 ( .A(n653), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U726 ( .A(n654), .B(G122), .Z(G24) );
  NAND2_X1 U727 ( .A1(n661), .A2(G217), .ZN(n655) );
  NOR2_X1 U728 ( .A1(n657), .A2(n666), .ZN(G66) );
  NOR2_X1 U729 ( .A1(n660), .A2(n666), .ZN(G63) );
  NAND2_X1 U730 ( .A1(n661), .A2(G469), .ZN(n665) );
  XNOR2_X1 U731 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n662) );
  XNOR2_X1 U732 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U733 ( .A(n665), .B(n664), .ZN(n667) );
  NOR2_X1 U734 ( .A1(n667), .A2(n666), .ZN(G54) );
  INV_X1 U735 ( .A(n668), .ZN(n672) );
  INV_X1 U736 ( .A(n669), .ZN(n681) );
  NAND2_X1 U737 ( .A1(n672), .A2(n681), .ZN(n670) );
  XNOR2_X1 U738 ( .A(n670), .B(G104), .ZN(G6) );
  XOR2_X1 U739 ( .A(KEYINPUT113), .B(KEYINPUT26), .Z(n674) );
  INV_X1 U740 ( .A(n671), .ZN(n677) );
  NAND2_X1 U741 ( .A1(n672), .A2(n677), .ZN(n673) );
  XNOR2_X1 U742 ( .A(n674), .B(n673), .ZN(n676) );
  XOR2_X1 U743 ( .A(G107), .B(KEYINPUT27), .Z(n675) );
  XNOR2_X1 U744 ( .A(n676), .B(n675), .ZN(G9) );
  XOR2_X1 U745 ( .A(KEYINPUT29), .B(KEYINPUT114), .Z(n679) );
  NAND2_X1 U746 ( .A1(n682), .A2(n677), .ZN(n678) );
  XNOR2_X1 U747 ( .A(n679), .B(n678), .ZN(n680) );
  XNOR2_X1 U748 ( .A(G128), .B(n680), .ZN(G30) );
  NAND2_X1 U749 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U750 ( .A(n683), .B(G146), .ZN(G48) );
  INV_X1 U751 ( .A(n684), .ZN(n685) );
  XOR2_X1 U752 ( .A(G134), .B(n685), .Z(n686) );
  XNOR2_X1 U753 ( .A(KEYINPUT116), .B(n686), .ZN(G36) );
  NOR2_X1 U754 ( .A1(n688), .A2(n687), .ZN(n690) );
  XNOR2_X1 U755 ( .A(KEYINPUT49), .B(KEYINPUT117), .ZN(n689) );
  XNOR2_X1 U756 ( .A(n690), .B(n689), .ZN(n695) );
  NOR2_X1 U757 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U758 ( .A(n693), .B(KEYINPUT50), .ZN(n694) );
  NOR2_X1 U759 ( .A1(n695), .A2(n694), .ZN(n697) );
  NAND2_X1 U760 ( .A1(n697), .A2(n370), .ZN(n699) );
  NAND2_X1 U761 ( .A1(n699), .A2(n698), .ZN(n702) );
  XOR2_X1 U762 ( .A(KEYINPUT51), .B(KEYINPUT119), .Z(n700) );
  XNOR2_X1 U763 ( .A(KEYINPUT118), .B(n700), .ZN(n701) );
  XNOR2_X1 U764 ( .A(n702), .B(n701), .ZN(n703) );
  NOR2_X1 U765 ( .A1(n720), .A2(n703), .ZN(n716) );
  NAND2_X1 U766 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U767 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U768 ( .A(n708), .B(KEYINPUT120), .ZN(n712) );
  NAND2_X1 U769 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U770 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U771 ( .A(KEYINPUT121), .B(n713), .ZN(n714) );
  NOR2_X1 U772 ( .A1(n714), .A2(n721), .ZN(n715) );
  NOR2_X1 U773 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U774 ( .A(n717), .B(KEYINPUT52), .ZN(n718) );
  NOR2_X1 U775 ( .A1(n719), .A2(n718), .ZN(n723) );
  NOR2_X1 U776 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U777 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U778 ( .A1(n724), .A2(n753), .ZN(n731) );
  NOR2_X1 U779 ( .A1(n725), .A2(KEYINPUT2), .ZN(n726) );
  XNOR2_X1 U780 ( .A(n726), .B(KEYINPUT79), .ZN(n728) );
  NAND2_X1 U781 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U782 ( .A(n729), .B(KEYINPUT85), .ZN(n730) );
  NOR2_X1 U783 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U784 ( .A(n732), .B(KEYINPUT53), .ZN(G75) );
  NOR2_X1 U785 ( .A1(n733), .A2(G953), .ZN(n739) );
  NAND2_X1 U786 ( .A1(G953), .A2(G224), .ZN(n734) );
  XOR2_X1 U787 ( .A(KEYINPUT61), .B(n734), .Z(n735) );
  NOR2_X1 U788 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U789 ( .A(n737), .B(KEYINPUT124), .ZN(n738) );
  NOR2_X1 U790 ( .A1(n739), .A2(n738), .ZN(n746) );
  XNOR2_X1 U791 ( .A(n741), .B(G101), .ZN(n742) );
  XNOR2_X1 U792 ( .A(n359), .B(n742), .ZN(n744) );
  NAND2_X1 U793 ( .A1(n744), .A2(n743), .ZN(n745) );
  XOR2_X1 U794 ( .A(n746), .B(n745), .Z(n747) );
  XNOR2_X1 U795 ( .A(KEYINPUT125), .B(n747), .ZN(G69) );
  XOR2_X1 U796 ( .A(n748), .B(n749), .Z(n750) );
  XNOR2_X1 U797 ( .A(n751), .B(n750), .ZN(n755) );
  XNOR2_X1 U798 ( .A(n755), .B(n752), .ZN(n754) );
  NAND2_X1 U799 ( .A1(n754), .A2(n753), .ZN(n760) );
  XNOR2_X1 U800 ( .A(G227), .B(n755), .ZN(n756) );
  NAND2_X1 U801 ( .A1(n756), .A2(G900), .ZN(n757) );
  XNOR2_X1 U802 ( .A(KEYINPUT126), .B(n757), .ZN(n758) );
  NAND2_X1 U803 ( .A1(n758), .A2(G953), .ZN(n759) );
  NAND2_X1 U804 ( .A1(n760), .A2(n759), .ZN(G72) );
  XOR2_X1 U805 ( .A(G143), .B(n761), .Z(G45) );
  XOR2_X1 U806 ( .A(n762), .B(G125), .Z(n763) );
  XNOR2_X1 U807 ( .A(KEYINPUT37), .B(n763), .ZN(G27) );
  XNOR2_X1 U808 ( .A(n764), .B(G137), .ZN(G39) );
  XNOR2_X1 U809 ( .A(n765), .B(G131), .ZN(G33) );
endmodule

