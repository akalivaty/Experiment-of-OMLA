//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1215, new_n1216, new_n1217, new_n1219,
    new_n1220, new_n1221, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1277, new_n1278, new_n1279;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G13), .ZN(new_n208));
  NAND3_X1  g0008(.A1(new_n208), .A2(G1), .A3(G20), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT64), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n202), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n212), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(KEYINPUT65), .B(G244), .ZN(new_n219));
  AND2_X1   g0019(.A1(new_n219), .A2(G77), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G107), .A2(G264), .ZN(new_n224));
  NAND4_X1  g0024(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G1), .ZN(new_n226));
  OAI22_X1  g0026(.A1(new_n220), .A2(new_n225), .B1(new_n226), .B2(new_n214), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT66), .Z(new_n228));
  INV_X1    g0028(.A(KEYINPUT1), .ZN(new_n229));
  OR2_X1    g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n228), .A2(new_n229), .ZN(new_n231));
  AND3_X1   g0031(.A1(new_n218), .A2(new_n230), .A3(new_n231), .ZN(G361));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(G226), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(new_n213), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NAND4_X1  g0055(.A1(new_n254), .A2(KEYINPUT7), .A3(new_n214), .A4(new_n255), .ZN(new_n256));
  AND2_X1   g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NOR3_X1   g0058(.A1(new_n257), .A2(new_n258), .A3(G20), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT7), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT74), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT74), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT7), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n256), .B1(new_n259), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G68), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT76), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n214), .A2(new_n253), .ZN(new_n268));
  INV_X1    g0068(.A(G159), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(G20), .A2(G33), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(KEYINPUT76), .A3(G159), .ZN(new_n272));
  XNOR2_X1  g0072(.A(G58), .B(G68), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n270), .A2(new_n272), .B1(new_n273), .B2(G20), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n266), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n251), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n254), .A2(new_n214), .A3(new_n255), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT74), .B(KEYINPUT7), .ZN(new_n279));
  OAI21_X1  g0079(.A(KEYINPUT75), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n257), .A2(new_n258), .ZN(new_n281));
  AOI21_X1  g0081(.A(KEYINPUT7), .B1(new_n281), .B2(new_n214), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT75), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n264), .A2(new_n281), .A3(new_n284), .A4(new_n214), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G68), .ZN(new_n286));
  OAI211_X1 g0086(.A(KEYINPUT16), .B(new_n274), .C1(new_n283), .C2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n226), .A2(G13), .A3(G20), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(new_n250), .ZN(new_n290));
  OR3_X1    g0090(.A1(new_n214), .A2(KEYINPUT70), .A3(G1), .ZN(new_n291));
  OAI21_X1  g0091(.A(KEYINPUT70), .B1(new_n214), .B2(G1), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(KEYINPUT8), .B(G58), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n290), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n289), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT78), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n296), .A2(KEYINPUT78), .A3(new_n297), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n277), .A2(new_n287), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G200), .ZN(new_n303));
  NAND2_X1  g0103(.A1(G33), .A2(G41), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n304), .A2(G1), .A3(G13), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n226), .B1(G41), .B2(G45), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n305), .A2(G232), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT79), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n307), .B(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n306), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n310), .A2(new_n305), .A3(G274), .ZN(new_n311));
  INV_X1    g0111(.A(G87), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n253), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(G223), .A2(G1698), .ZN(new_n314));
  INV_X1    g0114(.A(G226), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n314), .B1(new_n315), .B2(G1698), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n254), .A2(new_n255), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n313), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n311), .B1(new_n318), .B2(new_n305), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n303), .B1(new_n309), .B2(new_n319), .ZN(new_n320));
  XNOR2_X1  g0120(.A(new_n307), .B(KEYINPUT79), .ZN(new_n321));
  INV_X1    g0121(.A(G190), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n315), .A2(G1698), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(G223), .B2(G1698), .ZN(new_n324));
  OAI22_X1  g0124(.A1(new_n324), .A2(new_n281), .B1(new_n253), .B2(new_n312), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n321), .A2(new_n322), .A3(new_n311), .A4(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n320), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n302), .A2(KEYINPUT17), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G68), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n278), .A2(new_n279), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n331), .B1(new_n332), .B2(new_n256), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n270), .A2(new_n272), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n273), .A2(G20), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n276), .B1(new_n333), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n287), .A2(new_n250), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n300), .A2(new_n301), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n329), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT17), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n330), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT18), .ZN(new_n344));
  OAI21_X1  g0144(.A(G169), .B1(new_n309), .B2(new_n319), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n321), .A2(G179), .A3(new_n311), .A4(new_n327), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n344), .B1(new_n302), .B2(new_n348), .ZN(new_n349));
  AOI221_X4 g0149(.A(new_n344), .B1(new_n345), .B2(new_n346), .C1(new_n338), .C2(new_n339), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n349), .B1(new_n350), .B2(KEYINPUT80), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n338), .A2(new_n339), .B1(new_n345), .B2(new_n346), .ZN(new_n352));
  OR3_X1    g0152(.A1(new_n352), .A2(KEYINPUT80), .A3(KEYINPUT18), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n343), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT9), .ZN(new_n356));
  INV_X1    g0156(.A(G50), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n214), .B1(new_n201), .B2(new_n357), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n358), .B(KEYINPUT69), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n214), .A2(G33), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n295), .A2(new_n361), .B1(G150), .B2(new_n271), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n251), .B1(new_n359), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n290), .A2(new_n293), .A3(G50), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(G50), .B2(new_n288), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n356), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT71), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI211_X1 g0168(.A(KEYINPUT71), .B(new_n356), .C1(new_n363), .C2(new_n365), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT72), .ZN(new_n371));
  INV_X1    g0171(.A(G1698), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n317), .A2(G222), .A3(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n317), .A2(G223), .A3(G1698), .ZN(new_n374));
  INV_X1    g0174(.A(G77), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n373), .B(new_n374), .C1(new_n375), .C2(new_n317), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n326), .ZN(new_n377));
  AND3_X1   g0177(.A1(new_n310), .A2(new_n305), .A3(G274), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n326), .A2(new_n310), .ZN(new_n379));
  XOR2_X1   g0179(.A(KEYINPUT68), .B(G226), .Z(new_n380));
  AOI21_X1  g0180(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n371), .B1(new_n382), .B2(new_n322), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n377), .A2(KEYINPUT72), .A3(G190), .A4(new_n381), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n363), .A2(new_n365), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n386), .A2(KEYINPUT9), .B1(new_n382), .B2(G200), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n370), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT10), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT10), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n370), .A2(new_n385), .A3(new_n390), .A4(new_n387), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(G169), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n386), .B1(new_n393), .B2(new_n382), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(G179), .B2(new_n382), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n378), .B1(G238), .B2(new_n379), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n317), .A2(G232), .A3(G1698), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G33), .A2(G97), .ZN(new_n399));
  OAI211_X1 g0199(.A(G226), .B(new_n372), .C1(new_n257), .C2(new_n258), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n326), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT13), .ZN(new_n403));
  AND3_X1   g0203(.A1(new_n397), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n403), .B1(new_n397), .B2(new_n402), .ZN(new_n405));
  OAI21_X1  g0205(.A(G169), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT14), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n397), .A2(new_n402), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT13), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n397), .A2(new_n402), .A3(new_n403), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT14), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(new_n412), .A3(G169), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n409), .A2(G179), .A3(new_n410), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n407), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n289), .A2(new_n331), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n416), .B(KEYINPUT12), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n271), .A2(G50), .B1(G20), .B2(new_n331), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n375), .B2(new_n360), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n419), .A2(KEYINPUT11), .A3(new_n250), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n290), .A2(new_n293), .A3(G68), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n417), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT11), .B1(new_n419), .B2(new_n250), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n415), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n375), .B1(new_n291), .B2(new_n292), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n427), .A2(new_n290), .B1(new_n375), .B2(new_n289), .ZN(new_n428));
  OAI22_X1  g0228(.A1(new_n294), .A2(new_n268), .B1(new_n214), .B2(new_n375), .ZN(new_n429));
  XNOR2_X1  g0229(.A(KEYINPUT15), .B(G87), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n430), .A2(new_n360), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n250), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n317), .A2(G232), .A3(new_n372), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n317), .A2(G238), .A3(G1698), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n434), .B(new_n435), .C1(new_n205), .C2(new_n317), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n326), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n378), .B1(new_n219), .B2(new_n379), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n433), .B1(new_n440), .B2(G190), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(new_n303), .B2(new_n440), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n439), .A2(new_n393), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n443), .B(new_n433), .C1(G179), .C2(new_n439), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n426), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(G200), .B1(new_n404), .B2(new_n405), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n409), .A2(G190), .A3(new_n410), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n446), .A2(new_n447), .A3(new_n424), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT73), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n446), .A2(new_n447), .A3(KEYINPUT73), .A4(new_n424), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g0253(.A1(new_n355), .A2(new_n396), .A3(new_n445), .A4(new_n453), .ZN(new_n454));
  OAI211_X1 g0254(.A(G257), .B(G1698), .C1(new_n257), .C2(new_n258), .ZN(new_n455));
  OAI211_X1 g0255(.A(G250), .B(new_n372), .C1(new_n257), .C2(new_n258), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G33), .A2(G294), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n326), .ZN(new_n459));
  INV_X1    g0259(.A(G45), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n460), .A2(G1), .ZN(new_n461));
  XNOR2_X1  g0261(.A(KEYINPUT5), .B(G41), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n326), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G264), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n462), .A2(G274), .A3(new_n305), .A4(new_n461), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n459), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT86), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n466), .A2(new_n467), .A3(new_n303), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n467), .B1(new_n466), .B2(new_n303), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n466), .A2(KEYINPUT85), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n326), .A2(new_n458), .B1(new_n463), .B2(G264), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT85), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n472), .A2(new_n473), .A3(new_n465), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n322), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n470), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT24), .ZN(new_n478));
  OR2_X1    g0278(.A1(new_n478), .A2(KEYINPUT84), .ZN(new_n479));
  OAI21_X1  g0279(.A(KEYINPUT23), .B1(new_n214), .B2(G107), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT23), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n481), .A2(new_n205), .A3(G20), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n214), .A2(G33), .A3(G116), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n479), .A2(new_n480), .A3(new_n482), .A4(new_n483), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n214), .B(G87), .C1(new_n257), .C2(new_n258), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(KEYINPUT22), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT22), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n317), .A2(new_n487), .A3(new_n214), .A4(G87), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n484), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n478), .A2(KEYINPUT84), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  AOI211_X1 g0292(.A(new_n490), .B(new_n484), .C1(new_n486), .C2(new_n488), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n250), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n226), .A2(G33), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n288), .A2(new_n495), .A3(new_n213), .A4(new_n249), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n289), .A2(KEYINPUT25), .A3(new_n205), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT25), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(new_n288), .B2(G107), .ZN(new_n500));
  AOI22_X1  g0300(.A1(G107), .A2(new_n497), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  AND2_X1   g0301(.A1(new_n494), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n477), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g0303(.A(G250), .B(G1698), .C1(new_n257), .C2(new_n258), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G283), .ZN(new_n505));
  OAI211_X1 g0305(.A(G244), .B(new_n372), .C1(new_n257), .C2(new_n258), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT4), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n504), .B(new_n505), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n506), .A2(new_n507), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n326), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AND2_X1   g0310(.A1(KEYINPUT5), .A2(G41), .ZN(new_n511));
  NOR2_X1   g0311(.A1(KEYINPUT5), .A2(G41), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n461), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n513), .A2(G257), .A3(new_n305), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n465), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT81), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n514), .A2(KEYINPUT81), .A3(new_n465), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n510), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n393), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT6), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n521), .A2(new_n204), .A3(G107), .ZN(new_n522));
  XNOR2_X1  g0322(.A(G97), .B(G107), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n522), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  OAI22_X1  g0324(.A1(new_n524), .A2(new_n214), .B1(new_n375), .B2(new_n268), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n205), .B1(new_n332), .B2(new_n256), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n250), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n289), .A2(new_n204), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n497), .A2(G97), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n514), .A2(KEYINPUT81), .A3(new_n465), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT81), .B1(new_n514), .B2(new_n465), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(G179), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n533), .A2(new_n534), .A3(new_n510), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n520), .A2(new_n530), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n519), .A2(G200), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n529), .A2(new_n528), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n523), .A2(new_n521), .ZN(new_n539));
  INV_X1    g0339(.A(new_n522), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n541), .A2(G20), .B1(G77), .B2(new_n271), .ZN(new_n542));
  INV_X1    g0342(.A(new_n526), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n538), .B1(new_n544), .B2(new_n250), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n533), .A2(G190), .A3(new_n510), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n537), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n317), .A2(new_n214), .A3(G68), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT19), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n214), .B1(new_n399), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n550), .B1(G87), .B2(new_n206), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n549), .B1(new_n360), .B2(new_n204), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n548), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n553), .A2(new_n250), .B1(new_n289), .B2(new_n430), .ZN(new_n554));
  INV_X1    g0354(.A(new_n430), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n497), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(G244), .B(G1698), .C1(new_n257), .C2(new_n258), .ZN(new_n558));
  OAI211_X1 g0358(.A(G238), .B(new_n372), .C1(new_n257), .C2(new_n258), .ZN(new_n559));
  INV_X1    g0359(.A(G116), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n558), .B(new_n559), .C1(new_n253), .C2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n326), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n305), .A2(G274), .A3(new_n461), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n226), .A2(G45), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n305), .A2(G250), .A3(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n563), .A2(new_n565), .A3(KEYINPUT82), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(KEYINPUT82), .B1(new_n563), .B2(new_n565), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n562), .B(new_n534), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n568), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n570), .A2(new_n566), .B1(new_n326), .B2(new_n561), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n557), .B(new_n569), .C1(new_n571), .C2(G169), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n562), .B1(new_n567), .B2(new_n568), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(G200), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n562), .B(G190), .C1(new_n567), .C2(new_n568), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n497), .A2(G87), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n574), .A2(new_n554), .A3(new_n575), .A4(new_n576), .ZN(new_n577));
  AND4_X1   g0377(.A1(new_n536), .A2(new_n547), .A3(new_n572), .A4(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n513), .A2(G270), .A3(new_n305), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n465), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(G264), .B(G1698), .C1(new_n257), .C2(new_n258), .ZN(new_n582));
  OAI211_X1 g0382(.A(G257), .B(new_n372), .C1(new_n257), .C2(new_n258), .ZN(new_n583));
  INV_X1    g0383(.A(G303), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n582), .B(new_n583), .C1(new_n584), .C2(new_n317), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n326), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n505), .B(new_n214), .C1(G33), .C2(new_n204), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT20), .ZN(new_n589));
  AOI22_X1  g0389(.A1(KEYINPUT83), .A2(new_n589), .B1(new_n560), .B2(G20), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n590), .A3(new_n250), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n589), .A2(KEYINPUT83), .ZN(new_n592));
  OR2_X1    g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n288), .A2(new_n560), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n497), .B2(new_n560), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT83), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n591), .A2(new_n596), .A3(KEYINPUT20), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n593), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n587), .A2(new_n598), .A3(G169), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT21), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n598), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n581), .A2(new_n586), .A3(G190), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n580), .B1(new_n326), .B2(new_n585), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n602), .B(new_n603), .C1(new_n604), .C2(new_n303), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n587), .A2(new_n534), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n598), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n587), .A2(new_n598), .A3(KEYINPUT21), .A4(G169), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n601), .A2(new_n605), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n471), .A2(new_n474), .A3(G169), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n472), .A2(G179), .A3(new_n465), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n610), .A2(new_n611), .B1(new_n494), .B2(new_n501), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  AND4_X1   g0413(.A1(new_n454), .A2(new_n503), .A3(new_n578), .A4(new_n613), .ZN(G372));
  INV_X1    g0414(.A(new_n395), .ZN(new_n615));
  INV_X1    g0415(.A(new_n350), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n349), .ZN(new_n617));
  INV_X1    g0417(.A(new_n444), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n415), .A2(new_n425), .B1(new_n448), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n617), .B1(new_n619), .B2(new_n343), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT87), .ZN(new_n621));
  OR2_X1    g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n389), .A2(new_n391), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n623), .B1(new_n620), .B2(new_n621), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n615), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n601), .A2(new_n607), .A3(new_n608), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n578), .B(new_n503), .C1(new_n612), .C2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n572), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n554), .A2(new_n576), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n629), .B1(G200), .B2(new_n573), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n573), .A2(new_n393), .B1(new_n554), .B2(new_n556), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n630), .A2(new_n575), .B1(new_n631), .B2(new_n569), .ZN(new_n632));
  INV_X1    g0432(.A(new_n536), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(KEYINPUT26), .A3(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT26), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n577), .A2(new_n572), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n635), .B1(new_n636), .B2(new_n536), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n628), .B1(new_n634), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n627), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n454), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n625), .A2(new_n640), .ZN(G369));
  NAND3_X1  g0441(.A1(new_n226), .A2(new_n214), .A3(G13), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(new_n644), .A3(G213), .ZN(new_n645));
  INV_X1    g0445(.A(G343), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n602), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n626), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n650), .B1(new_n609), .B2(new_n649), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(G330), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n612), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n494), .A2(new_n501), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n657), .B1(new_n470), .B2(new_n476), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n502), .A2(new_n648), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n656), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n612), .A2(new_n648), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n655), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n626), .A2(new_n648), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n660), .A2(new_n666), .B1(new_n612), .B2(new_n648), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(new_n667), .ZN(G399));
  INV_X1    g0468(.A(G41), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n210), .A2(KEYINPUT88), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(KEYINPUT88), .B1(new_n210), .B2(new_n669), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(KEYINPUT89), .B1(new_n672), .B2(new_n217), .ZN(new_n673));
  INV_X1    g0473(.A(new_n672), .ZN(new_n674));
  NOR3_X1   g0474(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G1), .A3(new_n675), .ZN(new_n676));
  MUX2_X1   g0476(.A(KEYINPUT89), .B(new_n673), .S(new_n676), .Z(new_n677));
  XOR2_X1   g0477(.A(new_n677), .B(KEYINPUT28), .Z(new_n678));
  INV_X1    g0478(.A(KEYINPUT30), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n571), .A2(new_n533), .A3(new_n472), .A4(new_n510), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n604), .A2(G179), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n679), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n571), .A2(new_n472), .ZN(new_n683));
  INV_X1    g0483(.A(new_n519), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n683), .A2(new_n684), .A3(new_n606), .A4(KEYINPUT30), .ZN(new_n685));
  NOR3_X1   g0485(.A1(new_n571), .A2(new_n604), .A3(G179), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n686), .A2(new_n466), .A3(new_n519), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n682), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n647), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n578), .A2(new_n613), .A3(new_n503), .A4(new_n648), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n690), .B1(new_n691), .B2(KEYINPUT31), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n688), .A2(KEYINPUT31), .A3(new_n647), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT90), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT90), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n688), .A2(new_n695), .A3(KEYINPUT31), .A4(new_n647), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n692), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G330), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n647), .B1(new_n627), .B2(new_n638), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT29), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n700), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n678), .B1(new_n705), .B2(G1), .ZN(G364));
  NOR2_X1   g0506(.A1(new_n208), .A2(G20), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n226), .B1(new_n707), .B2(G45), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n672), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n210), .A2(new_n317), .ZN(new_n711));
  INV_X1    g0511(.A(G355), .ZN(new_n712));
  OAI22_X1  g0512(.A1(new_n711), .A2(new_n712), .B1(G116), .B2(new_n210), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n210), .A2(new_n281), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT91), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n216), .A2(G45), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n716), .B1(new_n247), .B2(G45), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n713), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(G13), .A2(G33), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(G20), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT92), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n213), .B1(G20), .B2(new_n393), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n710), .B1(new_n718), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n214), .A2(G179), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n728), .A2(new_n322), .A3(G200), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(new_n205), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n728), .A2(new_n322), .A3(new_n303), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n732), .A2(KEYINPUT32), .A3(G159), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT32), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(new_n731), .B2(new_n269), .ZN(new_n735));
  AOI211_X1 g0535(.A(new_n281), .B(new_n730), .C1(new_n733), .C2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n214), .A2(new_n534), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(new_n322), .A3(G200), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n728), .A2(G190), .A3(G200), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI22_X1  g0541(.A1(G68), .A2(new_n739), .B1(new_n741), .B2(G87), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n322), .A2(G179), .A3(G200), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n214), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(new_n204), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n737), .A2(G190), .A3(G200), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n745), .B1(G50), .B2(new_n747), .ZN(new_n748));
  AND3_X1   g0548(.A1(new_n736), .A2(new_n742), .A3(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n737), .A2(KEYINPUT93), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G200), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n737), .A2(KEYINPUT93), .ZN(new_n752));
  AND3_X1   g0552(.A1(new_n751), .A2(new_n322), .A3(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n751), .A2(G190), .A3(new_n752), .ZN(new_n755));
  XOR2_X1   g0555(.A(new_n755), .B(KEYINPUT94), .Z(new_n756));
  INV_X1    g0556(.A(G58), .ZN(new_n757));
  OAI221_X1 g0557(.A(new_n749), .B1(new_n375), .B2(new_n754), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n755), .ZN(new_n759));
  AOI22_X1  g0559(.A1(G322), .A2(new_n759), .B1(new_n753), .B2(G311), .ZN(new_n760));
  INV_X1    g0560(.A(G294), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n744), .A2(new_n761), .ZN(new_n762));
  AOI211_X1 g0562(.A(new_n317), .B(new_n762), .C1(G329), .C2(new_n732), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n740), .A2(new_n584), .ZN(new_n764));
  XOR2_X1   g0564(.A(KEYINPUT33), .B(G317), .Z(new_n765));
  INV_X1    g0565(.A(G283), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n738), .A2(new_n765), .B1(new_n729), .B2(new_n766), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n764), .B(new_n767), .C1(G326), .C2(new_n747), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n760), .A2(new_n763), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n758), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n727), .B1(new_n770), .B2(new_n724), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(new_n651), .B2(new_n722), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT95), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n651), .A2(G330), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n654), .A2(new_n710), .A3(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(G396));
  NOR2_X1   g0577(.A1(new_n444), .A2(new_n647), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n433), .A2(new_n647), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n442), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n778), .B1(new_n780), .B2(new_n444), .ZN(new_n781));
  OR2_X1    g0581(.A1(new_n701), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(KEYINPUT26), .B1(new_n632), .B2(new_n633), .ZN(new_n783));
  NOR3_X1   g0583(.A1(new_n636), .A2(new_n635), .A3(new_n536), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n572), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n612), .A2(new_n626), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n547), .A2(new_n536), .A3(new_n572), .A4(new_n577), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n786), .A2(new_n787), .A3(new_n658), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n648), .B(new_n781), .C1(new_n785), .C2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n782), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n710), .B1(new_n790), .B2(new_n699), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(new_n699), .B2(new_n790), .ZN(new_n792));
  INV_X1    g0592(.A(new_n724), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(new_n720), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n710), .B1(G77), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI22_X1  g0596(.A1(G294), .A2(new_n759), .B1(new_n753), .B2(G116), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n317), .B(new_n745), .C1(G311), .C2(new_n732), .ZN(new_n798));
  INV_X1    g0598(.A(new_n729), .ZN(new_n799));
  AOI22_X1  g0599(.A1(G283), .A2(new_n739), .B1(new_n799), .B2(G87), .ZN(new_n800));
  AOI22_X1  g0600(.A1(G303), .A2(new_n747), .B1(new_n741), .B2(G107), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n797), .A2(new_n798), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT96), .Z(new_n803));
  INV_X1    g0603(.A(G132), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n317), .B1(new_n731), .B2(new_n804), .C1(new_n331), .C2(new_n729), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n744), .A2(new_n757), .B1(new_n740), .B2(new_n357), .ZN(new_n806));
  AOI22_X1  g0606(.A1(G137), .A2(new_n747), .B1(new_n739), .B2(G150), .ZN(new_n807));
  INV_X1    g0607(.A(G143), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n807), .B1(new_n269), .B2(new_n754), .C1(new_n756), .C2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT34), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n805), .B(new_n806), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n803), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n796), .B1(new_n720), .B2(new_n781), .C1(new_n813), .C2(new_n793), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n792), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(G384));
  OR2_X1    g0616(.A1(new_n541), .A2(KEYINPUT35), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n541), .A2(KEYINPUT35), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n817), .A2(G116), .A3(new_n215), .A4(new_n818), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT36), .Z(new_n820));
  OAI211_X1 g0620(.A(new_n217), .B(G77), .C1(new_n757), .C2(new_n331), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n357), .A2(G68), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n226), .B(G13), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT39), .ZN(new_n825));
  AND3_X1   g0625(.A1(new_n329), .A2(new_n338), .A3(new_n339), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n645), .B1(new_n338), .B2(new_n339), .ZN(new_n827));
  NOR3_X1   g0627(.A1(new_n826), .A2(new_n352), .A3(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT37), .ZN(new_n829));
  OAI21_X1  g0629(.A(KEYINPUT98), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT99), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n828), .A2(new_n831), .A3(new_n829), .ZN(new_n832));
  INV_X1    g0632(.A(new_n352), .ZN(new_n833));
  INV_X1    g0633(.A(new_n827), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n833), .A2(new_n834), .A3(new_n340), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT98), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n835), .A2(new_n836), .A3(KEYINPUT37), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n833), .A2(new_n834), .A3(new_n829), .A4(new_n340), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(KEYINPUT99), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n830), .A2(new_n832), .A3(new_n837), .A4(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n617), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n827), .B1(new_n841), .B2(new_n343), .ZN(new_n842));
  AOI21_X1  g0642(.A(KEYINPUT38), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n278), .A2(new_n279), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n331), .B1(new_n844), .B2(new_n284), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n278), .A2(new_n260), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n846), .B(KEYINPUT75), .C1(new_n278), .C2(new_n279), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n336), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n251), .B1(new_n848), .B2(KEYINPUT16), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT97), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n276), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  AOI211_X1 g0651(.A(KEYINPUT97), .B(new_n336), .C1(new_n845), .C2(new_n847), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n849), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n298), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n348), .A2(new_n645), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n826), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n838), .B1(new_n857), .B2(new_n829), .ZN(new_n858));
  INV_X1    g0658(.A(new_n645), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  OAI211_X1 g0660(.A(KEYINPUT38), .B(new_n858), .C1(new_n354), .C2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n825), .B1(new_n843), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n426), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n648), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n858), .B1(new_n354), .B2(new_n860), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT38), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n869), .A2(KEYINPUT39), .A3(new_n861), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n863), .A2(new_n866), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n869), .A2(new_n861), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n424), .A2(new_n648), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n415), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n874), .B1(new_n452), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n448), .A2(new_n874), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n877), .B1(new_n415), .B2(new_n425), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n778), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n879), .B1(new_n789), .B2(new_n880), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n872), .A2(new_n881), .B1(new_n841), .B2(new_n645), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n871), .A2(KEYINPUT100), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT100), .B1(new_n871), .B2(new_n882), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n454), .B1(new_n704), .B2(new_n703), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n625), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n885), .B(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT40), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n840), .A2(new_n842), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n868), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n861), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n781), .B1(new_n876), .B2(new_n878), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n691), .A2(KEYINPUT31), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n689), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n693), .B(KEYINPUT101), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n893), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n889), .B1(new_n892), .B2(new_n897), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n872), .A2(new_n897), .A3(new_n889), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n895), .A2(new_n896), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n454), .A2(new_n901), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n900), .A2(new_n902), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n903), .A2(G330), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n888), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n226), .B2(new_n707), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n888), .A2(new_n905), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n824), .B1(new_n907), .B2(new_n908), .ZN(G367));
  INV_X1    g0709(.A(KEYINPUT105), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n547), .B(new_n536), .C1(new_n545), .C2(new_n648), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n536), .B2(new_n648), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n667), .A2(new_n912), .ZN(new_n913));
  OR2_X1    g0713(.A1(new_n913), .A2(KEYINPUT44), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n914), .A2(KEYINPUT104), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n914), .A2(KEYINPUT104), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n913), .A2(KEYINPUT44), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n667), .A2(new_n912), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n920), .A2(KEYINPUT103), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(KEYINPUT103), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n923), .A2(KEYINPUT45), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n923), .A2(KEYINPUT45), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n664), .B1(new_n919), .B2(new_n926), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n918), .B(new_n665), .C1(new_n924), .C2(new_n925), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n662), .B(new_n666), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(new_n654), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n705), .A2(new_n931), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n705), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n672), .B(KEYINPUT41), .Z(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n910), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  AOI211_X1 g0737(.A(KEYINPUT105), .B(new_n935), .C1(new_n933), .C2(new_n705), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n708), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n662), .A2(new_n666), .A3(new_n912), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n536), .B1(new_n911), .B2(new_n656), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n940), .A2(KEYINPUT42), .B1(new_n648), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(KEYINPUT42), .B2(new_n940), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n629), .A2(new_n647), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n632), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n572), .B2(new_n944), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(KEYINPUT43), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n943), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n946), .A2(KEYINPUT43), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n948), .B(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(KEYINPUT102), .B1(new_n664), .B2(new_n912), .ZN(new_n951));
  AND3_X1   g0751(.A1(new_n664), .A2(KEYINPUT102), .A3(new_n912), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n939), .B(new_n953), .C1(new_n951), .C2(new_n950), .ZN(new_n954));
  INV_X1    g0754(.A(G317), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n281), .B1(new_n731), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(KEYINPUT46), .B1(new_n741), .B2(G116), .ZN(new_n957));
  AOI211_X1 g0757(.A(new_n956), .B(new_n957), .C1(G311), .C2(new_n747), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n741), .A2(KEYINPUT46), .A3(G116), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n753), .A2(G283), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n729), .A2(new_n204), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n738), .A2(new_n761), .ZN(new_n962));
  INV_X1    g0762(.A(new_n744), .ZN(new_n963));
  AOI211_X1 g0763(.A(new_n961), .B(new_n962), .C1(G107), .C2(new_n963), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n958), .A2(new_n959), .A3(new_n960), .A4(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n756), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n965), .B1(G303), .B2(new_n966), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n738), .A2(new_n269), .B1(new_n746), .B2(new_n808), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n744), .A2(new_n331), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n729), .A2(new_n375), .ZN(new_n970));
  NOR3_X1   g0770(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(G137), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n317), .B1(new_n731), .B2(new_n973), .C1(new_n757), .C2(new_n740), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  AOI22_X1  g0775(.A1(G150), .A2(new_n759), .B1(new_n753), .B2(G50), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n967), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n977), .A2(KEYINPUT47), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(KEYINPUT47), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n978), .A2(new_n724), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n715), .A2(new_n240), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n981), .B(new_n725), .C1(new_n210), .C2(new_n430), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n710), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT106), .Z(new_n984));
  OAI211_X1 g0784(.A(new_n980), .B(new_n984), .C1(new_n722), .C2(new_n946), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n954), .A2(new_n985), .ZN(G387));
  NAND2_X1  g0786(.A1(new_n931), .A2(new_n709), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G311), .A2(new_n739), .B1(new_n747), .B2(G322), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n988), .B1(new_n584), .B2(new_n754), .C1(new_n756), .C2(new_n955), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT48), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n990), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n963), .A2(G283), .B1(new_n741), .B2(G294), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT49), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n996), .A2(KEYINPUT108), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(KEYINPUT108), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n729), .A2(new_n560), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n317), .B(new_n999), .C1(G326), .C2(new_n732), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n997), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(G50), .A2(new_n759), .B1(new_n753), .B2(G68), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n281), .B(new_n961), .C1(G150), .C2(new_n732), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(G159), .A2(new_n747), .B1(new_n741), .B2(G77), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n555), .A2(new_n963), .B1(new_n739), .B2(new_n295), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n793), .B1(new_n1001), .B2(new_n1006), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n711), .A2(new_n675), .B1(G107), .B2(new_n210), .ZN(new_n1008));
  XOR2_X1   g0808(.A(KEYINPUT107), .B(KEYINPUT50), .Z(new_n1009));
  OR3_X1    g0809(.A1(new_n1009), .A2(G50), .A3(new_n294), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1009), .B1(G50), .B2(new_n294), .ZN(new_n1011));
  AOI21_X1  g0811(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1010), .A2(new_n675), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  AND2_X1   g0813(.A1(new_n715), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n237), .A2(G45), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1008), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n710), .B1(new_n726), .B2(new_n1016), .C1(new_n662), .C2(new_n722), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n932), .A2(new_n672), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n705), .A2(new_n931), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n987), .B1(new_n1007), .B2(new_n1017), .C1(new_n1018), .C2(new_n1019), .ZN(G393));
  NAND2_X1  g0820(.A1(new_n929), .A2(new_n932), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n933), .A2(new_n672), .A3(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n929), .A2(new_n708), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n912), .A2(new_n722), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n715), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1025), .A2(new_n244), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n725), .B1(new_n204), .B2(new_n210), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n710), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(G150), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n755), .A2(new_n269), .B1(new_n1029), .B2(new_n746), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT51), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n744), .A2(new_n375), .B1(new_n738), .B2(new_n357), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n317), .B1(new_n731), .B2(new_n808), .C1(new_n312), .C2(new_n729), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n1032), .B(new_n1033), .C1(G68), .C2(new_n741), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1031), .B(new_n1034), .C1(new_n294), .C2(new_n754), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(G116), .A2(new_n963), .B1(new_n739), .B2(G303), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n754), .B2(new_n761), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT109), .Z(new_n1038));
  INV_X1    g0838(.A(G322), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n281), .B1(new_n731), .B2(new_n1039), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n730), .B(new_n1040), .C1(G283), .C2(new_n741), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n759), .A2(G311), .B1(G317), .B2(new_n747), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT52), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1035), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1028), .B1(new_n1045), .B2(new_n724), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1023), .B1(new_n1024), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1022), .A2(new_n1047), .ZN(G390));
  INV_X1    g0848(.A(KEYINPUT111), .ZN(new_n1049));
  OAI211_X1 g0849(.A(G330), .B(new_n781), .C1(new_n692), .C2(new_n697), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1050), .A2(new_n879), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n781), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n452), .A2(new_n875), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n873), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n878), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1052), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT101), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n693), .B(new_n1057), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1056), .B(G330), .C1(new_n692), .C2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT110), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1051), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n789), .A2(new_n880), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n879), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n866), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n892), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n863), .A2(new_n870), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1061), .B(new_n1065), .C1(new_n1066), .C2(new_n1064), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1059), .A2(KEYINPUT110), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1064), .B1(new_n863), .B2(new_n870), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n843), .A2(new_n862), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n1070), .A2(new_n866), .A3(new_n881), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1068), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1067), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n653), .B1(new_n895), .B2(new_n896), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n454), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n886), .A2(new_n1075), .A3(new_n625), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1050), .A2(new_n879), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n1059), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n1062), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n698), .A2(G330), .A3(new_n781), .A4(new_n1063), .ZN(new_n1080));
  OAI211_X1 g0880(.A(G330), .B(new_n781), .C1(new_n1058), .C2(new_n692), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n879), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n778), .B1(new_n701), .B2(new_n781), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1080), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1076), .B1(new_n1079), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1049), .B1(new_n1073), .B2(new_n1086), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1067), .A2(new_n1085), .A3(new_n1072), .A4(KEYINPUT111), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n674), .B1(new_n1073), .B2(new_n1086), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n710), .B1(new_n295), .B2(new_n794), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(G107), .A2(new_n739), .B1(new_n747), .B2(G283), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n754), .B2(new_n204), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT113), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n755), .A2(new_n560), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n281), .B1(new_n731), .B2(new_n761), .C1(new_n312), .C2(new_n740), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n744), .A2(new_n375), .B1(new_n729), .B2(new_n331), .ZN(new_n1098));
  NOR4_X1   g0898(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  OR2_X1    g0900(.A1(new_n1100), .A2(KEYINPUT114), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(KEYINPUT114), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(G159), .A2(new_n963), .B1(new_n747), .B2(G128), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(G137), .A2(new_n739), .B1(new_n732), .B2(G125), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1103), .B(new_n1104), .C1(new_n755), .C2(new_n804), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(KEYINPUT54), .B(G143), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n741), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT53), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n740), .B2(new_n1029), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n753), .A2(new_n1107), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n317), .B1(new_n729), .B2(new_n357), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1112), .B(KEYINPUT112), .Z(new_n1113));
  NAND2_X1  g0913(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1101), .B(new_n1102), .C1(new_n1105), .C2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1092), .B1(new_n1115), .B2(new_n724), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n1066), .B2(new_n720), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n1073), .B2(new_n708), .ZN(new_n1118));
  OR2_X1    g0918(.A1(new_n1091), .A2(new_n1118), .ZN(G378));
  INV_X1    g0919(.A(KEYINPUT57), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n897), .ZN(new_n1121));
  OAI21_X1  g0921(.A(KEYINPUT40), .B1(new_n1121), .B2(new_n1070), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n872), .A2(new_n897), .A3(new_n889), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n653), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n883), .B2(new_n884), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n871), .A2(new_n882), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT100), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n871), .A2(new_n882), .A3(KEYINPUT100), .ZN(new_n1129));
  OAI21_X1  g0929(.A(G330), .B1(new_n898), .B2(new_n899), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1125), .A2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n386), .A2(new_n645), .ZN(new_n1133));
  XOR2_X1   g0933(.A(new_n396), .B(new_n1133), .Z(new_n1134));
  INV_X1    g0934(.A(KEYINPUT118), .ZN(new_n1135));
  OR2_X1    g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  XOR2_X1   g0936(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1137));
  NAND2_X1  g0937(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1137), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1132), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1125), .A2(new_n1131), .A3(new_n1141), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1076), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1120), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1076), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1089), .A2(new_n1148), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n1125), .A2(new_n1131), .A3(new_n1141), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1141), .B1(new_n1125), .B2(new_n1131), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1149), .A2(new_n1152), .A3(KEYINPUT57), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1147), .A2(new_n1153), .A3(new_n672), .ZN(new_n1154));
  NOR3_X1   g0954(.A1(new_n1150), .A2(new_n1151), .A3(new_n708), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1141), .A2(new_n719), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n710), .B1(G50), .B2(new_n794), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(KEYINPUT117), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n738), .A2(new_n204), .B1(new_n740), .B2(new_n375), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n746), .A2(new_n560), .B1(new_n729), .B2(new_n757), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n669), .B(new_n281), .C1(new_n731), .C2(new_n766), .ZN(new_n1161));
  NOR4_X1   g0961(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .A4(new_n969), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1162), .B1(new_n205), .B2(new_n755), .C1(new_n430), .C2(new_n754), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT58), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n253), .A2(new_n669), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT115), .ZN(new_n1166));
  AOI21_X1  g0966(.A(G50), .B1(new_n281), .B2(new_n669), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1163), .A2(new_n1164), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1166), .B1(G124), .B2(new_n732), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n740), .A2(new_n1106), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT116), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(G150), .A2(new_n963), .B1(new_n747), .B2(G125), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1171), .B(new_n1172), .C1(new_n804), .C2(new_n738), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n754), .A2(new_n973), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1173), .B(new_n1174), .C1(G128), .C2(new_n759), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT59), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1169), .B1(new_n269), .B2(new_n729), .C1(new_n1175), .C2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1175), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1178), .A2(KEYINPUT59), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1168), .B1(new_n1164), .B2(new_n1163), .C1(new_n1177), .C2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1158), .B1(new_n1180), .B2(new_n724), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1156), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1155), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1154), .A2(new_n1184), .ZN(G375));
  NAND2_X1  g0985(.A1(new_n1079), .A2(new_n1084), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(new_n709), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n710), .B1(G68), .B2(new_n794), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT120), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n281), .B1(new_n732), .B2(G128), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n757), .B2(new_n729), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n744), .A2(new_n357), .B1(new_n738), .B2(new_n1106), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n746), .A2(new_n804), .B1(new_n740), .B2(new_n269), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n1194), .B1(new_n1029), .B2(new_n754), .C1(new_n756), .C2(new_n973), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n740), .A2(new_n204), .B1(new_n731), .B2(new_n584), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT121), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1197), .B1(new_n766), .B2(new_n755), .C1(new_n205), .C2(new_n754), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n555), .A2(new_n963), .B1(new_n739), .B2(G116), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n970), .A2(new_n317), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1199), .B(new_n1200), .C1(new_n761), .C2(new_n746), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1195), .B1(new_n1198), .B2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1189), .B1(new_n724), .B2(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT122), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n1063), .B2(new_n720), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1187), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  OR3_X1    g1007(.A1(new_n1186), .A2(KEYINPUT119), .A3(new_n1148), .ZN(new_n1208));
  OAI21_X1  g1008(.A(KEYINPUT119), .B1(new_n1186), .B2(new_n1148), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1086), .A2(new_n936), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1207), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  XOR2_X1   g1012(.A(new_n1212), .B(KEYINPUT123), .Z(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(G381));
  NOR4_X1   g1014(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1091), .A2(new_n1118), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1215), .A2(new_n1216), .A3(new_n1213), .ZN(new_n1217));
  OR3_X1    g1017(.A1(G387), .A2(G375), .A3(new_n1217), .ZN(G407));
  NAND2_X1  g1018(.A1(new_n646), .A2(G213), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1216), .A2(new_n1220), .ZN(new_n1221));
  OAI211_X1 g1021(.A(G407), .B(G213), .C1(G375), .C2(new_n1221), .ZN(G409));
  XNOR2_X1  g1022(.A(G393), .B(G396), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1223), .A2(new_n1022), .A3(new_n1047), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1223), .B1(new_n1022), .B2(new_n1047), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n954), .A2(new_n985), .A3(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1226), .B1(new_n954), .B2(new_n985), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(KEYINPUT124), .B1(new_n1155), .B2(new_n1183), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT124), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1232), .B(new_n1182), .C1(new_n1145), .C2(new_n708), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1149), .A2(new_n1152), .A3(new_n936), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1231), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n1216), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1154), .A2(G378), .A3(new_n1184), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1186), .A2(new_n1148), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n674), .B1(new_n1239), .B2(KEYINPUT60), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1086), .A2(KEYINPUT60), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1240), .B1(new_n1210), .B2(new_n1241), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n1242), .A2(G384), .A3(new_n1207), .ZN(new_n1243));
  AOI21_X1  g1043(.A(G384), .B1(new_n1242), .B2(new_n1207), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1238), .A2(new_n1219), .A3(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT63), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1220), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1249), .A2(KEYINPUT63), .A3(new_n1245), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1238), .A2(new_n1219), .ZN(new_n1251));
  INV_X1    g1051(.A(G2897), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1245), .B1(new_n1252), .B2(new_n1219), .ZN(new_n1253));
  OAI211_X1 g1053(.A(G2897), .B(new_n1220), .C1(new_n1243), .C2(new_n1244), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT61), .B1(new_n1251), .B2(new_n1256), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1230), .A2(new_n1248), .A3(new_n1250), .A4(new_n1257), .ZN(new_n1258));
  OR2_X1    g1058(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT61), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1260), .B1(new_n1249), .B2(new_n1255), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT62), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1246), .A2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1249), .A2(KEYINPUT62), .A3(new_n1245), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1261), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT125), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1259), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1264), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT62), .B1(new_n1249), .B2(new_n1245), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1266), .B(new_n1257), .C1(new_n1268), .C2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1258), .B1(new_n1267), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(KEYINPUT126), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT126), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1274), .B(new_n1258), .C1(new_n1267), .C2(new_n1271), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1273), .A2(new_n1275), .ZN(G405));
  XNOR2_X1  g1076(.A(G375), .B(G378), .ZN(new_n1277));
  OR3_X1    g1077(.A1(new_n1243), .A2(new_n1244), .A3(KEYINPUT127), .ZN(new_n1278));
  XNOR2_X1  g1078(.A(new_n1277), .B(new_n1278), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1259), .B(new_n1279), .ZN(G402));
endmodule


