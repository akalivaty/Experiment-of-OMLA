

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U547 ( .A(n702), .ZN(n724) );
  OR2_X1 U548 ( .A1(n708), .A2(n707), .ZN(n709) );
  BUF_X1 U549 ( .A(n690), .Z(n543) );
  XNOR2_X1 U550 ( .A(n527), .B(n526), .ZN(n690) );
  NAND2_X1 U551 ( .A1(n515), .A2(n785), .ZN(n697) );
  XNOR2_X1 U552 ( .A(n518), .B(KEYINPUT65), .ZN(n757) );
  NAND2_X1 U553 ( .A1(n521), .A2(n519), .ZN(n518) );
  NOR2_X1 U554 ( .A1(n716), .A2(n715), .ZN(n720) );
  XNOR2_X1 U555 ( .A(n714), .B(KEYINPUT99), .ZN(n715) );
  INV_X1 U556 ( .A(KEYINPUT100), .ZN(n711) );
  INV_X1 U557 ( .A(KEYINPUT32), .ZN(n522) );
  XNOR2_X1 U558 ( .A(n746), .B(KEYINPUT101), .ZN(n747) );
  OR2_X1 U559 ( .A1(n696), .A2(n517), .ZN(n516) );
  INV_X1 U560 ( .A(G40), .ZN(n517) );
  NOR2_X1 U561 ( .A1(G164), .A2(G1384), .ZN(n785) );
  INV_X1 U562 ( .A(n958), .ZN(n520) );
  NAND2_X1 U563 ( .A1(n528), .A2(G2105), .ZN(n527) );
  INV_X1 U564 ( .A(G2104), .ZN(n528) );
  OR2_X1 U565 ( .A1(n760), .A2(n530), .ZN(n529) );
  NOR2_X1 U566 ( .A1(G651), .A2(n623), .ZN(n648) );
  INV_X1 U567 ( .A(G2105), .ZN(n537) );
  XOR2_X1 U568 ( .A(n721), .B(KEYINPUT28), .Z(n513) );
  OR2_X1 U569 ( .A1(n516), .A2(n695), .ZN(n784) );
  NOR2_X1 U570 ( .A1(n695), .A2(n696), .ZN(G160) );
  INV_X1 U571 ( .A(n784), .ZN(n515) );
  NOR2_X1 U572 ( .A1(n822), .A2(n520), .ZN(n519) );
  NAND2_X1 U573 ( .A1(n816), .A2(n962), .ZN(n521) );
  XNOR2_X1 U574 ( .A(n523), .B(n522), .ZN(n755) );
  NAND2_X1 U575 ( .A1(n524), .A2(n745), .ZN(n523) );
  NAND2_X1 U576 ( .A1(n525), .A2(n738), .ZN(n524) );
  XNOR2_X1 U577 ( .A(n748), .B(KEYINPUT101), .ZN(n525) );
  NAND2_X1 U578 ( .A1(n690), .A2(G125), .ZN(n691) );
  INV_X1 U579 ( .A(KEYINPUT66), .ZN(n526) );
  NOR2_X1 U580 ( .A1(n761), .A2(n760), .ZN(n531) );
  NOR2_X1 U581 ( .A1(n761), .A2(n529), .ZN(n813) );
  INV_X1 U582 ( .A(n976), .ZN(n530) );
  NAND2_X1 U583 ( .A1(n531), .A2(n827), .ZN(n833) );
  BUF_X1 U584 ( .A(n702), .Z(n739) );
  OR2_X1 U585 ( .A1(n822), .A2(n821), .ZN(n532) );
  NOR2_X2 U586 ( .A1(n623), .A2(n557), .ZN(n645) );
  XNOR2_X1 U587 ( .A(n603), .B(KEYINPUT15), .ZN(n971) );
  NOR2_X1 U588 ( .A1(G2104), .A2(G2105), .ZN(n533) );
  XOR2_X1 U589 ( .A(KEYINPUT17), .B(n533), .Z(n547) );
  NAND2_X1 U590 ( .A1(n896), .A2(G138), .ZN(n536) );
  NAND2_X1 U591 ( .A1(n690), .A2(G126), .ZN(n534) );
  XOR2_X1 U592 ( .A(KEYINPUT91), .B(n534), .Z(n535) );
  NAND2_X1 U593 ( .A1(n536), .A2(n535), .ZN(n542) );
  AND2_X4 U594 ( .A1(n537), .A2(G2104), .ZN(n897) );
  NAND2_X1 U595 ( .A1(G102), .A2(n897), .ZN(n540) );
  NAND2_X1 U596 ( .A1(G2105), .A2(G2104), .ZN(n538) );
  XOR2_X2 U597 ( .A(KEYINPUT70), .B(n538), .Z(n891) );
  NAND2_X1 U598 ( .A1(G114), .A2(n891), .ZN(n539) );
  NAND2_X1 U599 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U600 ( .A1(n542), .A2(n541), .ZN(G164) );
  AND2_X1 U601 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U602 ( .A1(G123), .A2(n543), .ZN(n544) );
  XNOR2_X1 U603 ( .A(n544), .B(KEYINPUT18), .ZN(n546) );
  NAND2_X1 U604 ( .A1(G99), .A2(n897), .ZN(n545) );
  NAND2_X1 U605 ( .A1(n546), .A2(n545), .ZN(n551) );
  BUF_X1 U606 ( .A(n547), .Z(n896) );
  NAND2_X1 U607 ( .A1(G135), .A2(n896), .ZN(n549) );
  NAND2_X1 U608 ( .A1(G111), .A2(n891), .ZN(n548) );
  NAND2_X1 U609 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U610 ( .A1(n551), .A2(n550), .ZN(n940) );
  XNOR2_X1 U611 ( .A(n940), .B(G2096), .ZN(n552) );
  XNOR2_X1 U612 ( .A(n552), .B(KEYINPUT81), .ZN(n553) );
  OR2_X1 U613 ( .A1(G2100), .A2(n553), .ZN(G156) );
  INV_X1 U614 ( .A(G132), .ZN(G219) );
  INV_X1 U615 ( .A(G82), .ZN(G220) );
  INV_X1 U616 ( .A(G120), .ZN(G236) );
  INV_X1 U617 ( .A(G69), .ZN(G235) );
  INV_X1 U618 ( .A(G57), .ZN(G237) );
  INV_X1 U619 ( .A(G651), .ZN(n557) );
  NOR2_X1 U620 ( .A1(G543), .A2(n557), .ZN(n554) );
  XOR2_X1 U621 ( .A(KEYINPUT1), .B(n554), .Z(n647) );
  NAND2_X1 U622 ( .A1(G65), .A2(n647), .ZN(n556) );
  XOR2_X1 U623 ( .A(KEYINPUT0), .B(G543), .Z(n623) );
  NAND2_X1 U624 ( .A1(G53), .A2(n648), .ZN(n555) );
  NAND2_X1 U625 ( .A1(n556), .A2(n555), .ZN(n561) );
  NAND2_X1 U626 ( .A1(G78), .A2(n645), .ZN(n559) );
  NOR2_X1 U627 ( .A1(G651), .A2(G543), .ZN(n651) );
  NAND2_X1 U628 ( .A1(G91), .A2(n651), .ZN(n558) );
  NAND2_X1 U629 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X1 U630 ( .A1(n561), .A2(n560), .ZN(n719) );
  INV_X1 U631 ( .A(n719), .ZN(G299) );
  NAND2_X1 U632 ( .A1(n651), .A2(G90), .ZN(n562) );
  XOR2_X1 U633 ( .A(KEYINPUT75), .B(n562), .Z(n564) );
  NAND2_X1 U634 ( .A1(n645), .A2(G77), .ZN(n563) );
  NAND2_X1 U635 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U636 ( .A(n565), .B(KEYINPUT9), .ZN(n567) );
  NAND2_X1 U637 ( .A1(G64), .A2(n647), .ZN(n566) );
  NAND2_X1 U638 ( .A1(n567), .A2(n566), .ZN(n570) );
  NAND2_X1 U639 ( .A1(n648), .A2(G52), .ZN(n568) );
  XOR2_X1 U640 ( .A(KEYINPUT74), .B(n568), .Z(n569) );
  NOR2_X1 U641 ( .A1(n570), .A2(n569), .ZN(G171) );
  NAND2_X1 U642 ( .A1(G89), .A2(n651), .ZN(n571) );
  XOR2_X1 U643 ( .A(KEYINPUT4), .B(n571), .Z(n572) );
  XNOR2_X1 U644 ( .A(n572), .B(KEYINPUT79), .ZN(n574) );
  NAND2_X1 U645 ( .A1(G76), .A2(n645), .ZN(n573) );
  NAND2_X1 U646 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U647 ( .A(KEYINPUT5), .B(n575), .ZN(n581) );
  NAND2_X1 U648 ( .A1(G63), .A2(n647), .ZN(n577) );
  NAND2_X1 U649 ( .A1(G51), .A2(n648), .ZN(n576) );
  NAND2_X1 U650 ( .A1(n577), .A2(n576), .ZN(n579) );
  XOR2_X1 U651 ( .A(KEYINPUT6), .B(KEYINPUT80), .Z(n578) );
  XNOR2_X1 U652 ( .A(n579), .B(n578), .ZN(n580) );
  NAND2_X1 U653 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U654 ( .A(KEYINPUT7), .B(n582), .ZN(G168) );
  XOR2_X1 U655 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U656 ( .A1(G7), .A2(G661), .ZN(n583) );
  XNOR2_X1 U657 ( .A(n583), .B(KEYINPUT76), .ZN(n584) );
  XNOR2_X1 U658 ( .A(KEYINPUT10), .B(n584), .ZN(G223) );
  INV_X1 U659 ( .A(G223), .ZN(n838) );
  NAND2_X1 U660 ( .A1(n838), .A2(G567), .ZN(n585) );
  XOR2_X1 U661 ( .A(KEYINPUT11), .B(n585), .Z(G234) );
  NAND2_X1 U662 ( .A1(n647), .A2(G56), .ZN(n586) );
  XNOR2_X1 U663 ( .A(KEYINPUT14), .B(n586), .ZN(n592) );
  NAND2_X1 U664 ( .A1(n651), .A2(G81), .ZN(n587) );
  XNOR2_X1 U665 ( .A(n587), .B(KEYINPUT12), .ZN(n589) );
  NAND2_X1 U666 ( .A1(G68), .A2(n645), .ZN(n588) );
  NAND2_X1 U667 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U668 ( .A(KEYINPUT13), .B(n590), .ZN(n591) );
  NAND2_X1 U669 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U670 ( .A(n593), .B(KEYINPUT77), .ZN(n595) );
  NAND2_X1 U671 ( .A1(n648), .A2(G43), .ZN(n594) );
  NAND2_X1 U672 ( .A1(n595), .A2(n594), .ZN(n966) );
  INV_X1 U673 ( .A(G860), .ZN(n608) );
  OR2_X1 U674 ( .A1(n966), .A2(n608), .ZN(G153) );
  INV_X1 U675 ( .A(G171), .ZN(G301) );
  NAND2_X1 U676 ( .A1(G868), .A2(G301), .ZN(n605) );
  NAND2_X1 U677 ( .A1(G54), .A2(n648), .ZN(n602) );
  NAND2_X1 U678 ( .A1(G92), .A2(n651), .ZN(n597) );
  NAND2_X1 U679 ( .A1(G66), .A2(n647), .ZN(n596) );
  NAND2_X1 U680 ( .A1(n597), .A2(n596), .ZN(n600) );
  NAND2_X1 U681 ( .A1(n645), .A2(G79), .ZN(n598) );
  XOR2_X1 U682 ( .A(KEYINPUT78), .B(n598), .Z(n599) );
  NOR2_X1 U683 ( .A1(n600), .A2(n599), .ZN(n601) );
  NAND2_X1 U684 ( .A1(n602), .A2(n601), .ZN(n603) );
  INV_X1 U685 ( .A(n971), .ZN(n707) );
  INV_X1 U686 ( .A(G868), .ZN(n667) );
  NAND2_X1 U687 ( .A1(n707), .A2(n667), .ZN(n604) );
  NAND2_X1 U688 ( .A1(n605), .A2(n604), .ZN(G284) );
  NOR2_X1 U689 ( .A1(G286), .A2(n667), .ZN(n607) );
  NOR2_X1 U690 ( .A1(G868), .A2(G299), .ZN(n606) );
  NOR2_X1 U691 ( .A1(n607), .A2(n606), .ZN(G297) );
  NAND2_X1 U692 ( .A1(n608), .A2(G559), .ZN(n609) );
  NAND2_X1 U693 ( .A1(n609), .A2(n971), .ZN(n610) );
  XNOR2_X1 U694 ( .A(n610), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U695 ( .A1(G868), .A2(n966), .ZN(n613) );
  NAND2_X1 U696 ( .A1(n971), .A2(G868), .ZN(n611) );
  NOR2_X1 U697 ( .A1(G559), .A2(n611), .ZN(n612) );
  NOR2_X1 U698 ( .A1(n613), .A2(n612), .ZN(G282) );
  NAND2_X1 U699 ( .A1(G67), .A2(n647), .ZN(n615) );
  NAND2_X1 U700 ( .A1(G55), .A2(n648), .ZN(n614) );
  NAND2_X1 U701 ( .A1(n615), .A2(n614), .ZN(n619) );
  NAND2_X1 U702 ( .A1(G80), .A2(n645), .ZN(n617) );
  NAND2_X1 U703 ( .A1(G93), .A2(n651), .ZN(n616) );
  NAND2_X1 U704 ( .A1(n617), .A2(n616), .ZN(n618) );
  OR2_X1 U705 ( .A1(n619), .A2(n618), .ZN(n666) );
  NAND2_X1 U706 ( .A1(G559), .A2(n971), .ZN(n620) );
  XNOR2_X1 U707 ( .A(n620), .B(n966), .ZN(n664) );
  XNOR2_X1 U708 ( .A(KEYINPUT82), .B(n664), .ZN(n621) );
  NOR2_X1 U709 ( .A1(G860), .A2(n621), .ZN(n622) );
  XOR2_X1 U710 ( .A(n666), .B(n622), .Z(G145) );
  NAND2_X1 U711 ( .A1(G87), .A2(n623), .ZN(n624) );
  XNOR2_X1 U712 ( .A(n624), .B(KEYINPUT84), .ZN(n627) );
  NAND2_X1 U713 ( .A1(G74), .A2(G651), .ZN(n625) );
  XOR2_X1 U714 ( .A(KEYINPUT83), .B(n625), .Z(n626) );
  NAND2_X1 U715 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U716 ( .A1(n647), .A2(n628), .ZN(n630) );
  NAND2_X1 U717 ( .A1(n648), .A2(G49), .ZN(n629) );
  NAND2_X1 U718 ( .A1(n630), .A2(n629), .ZN(G288) );
  NAND2_X1 U719 ( .A1(G75), .A2(n645), .ZN(n632) );
  NAND2_X1 U720 ( .A1(G88), .A2(n651), .ZN(n631) );
  NAND2_X1 U721 ( .A1(n632), .A2(n631), .ZN(n636) );
  NAND2_X1 U722 ( .A1(G62), .A2(n647), .ZN(n634) );
  NAND2_X1 U723 ( .A1(G50), .A2(n648), .ZN(n633) );
  NAND2_X1 U724 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U725 ( .A1(n636), .A2(n635), .ZN(G166) );
  NAND2_X1 U726 ( .A1(G86), .A2(n651), .ZN(n638) );
  NAND2_X1 U727 ( .A1(G61), .A2(n647), .ZN(n637) );
  NAND2_X1 U728 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U729 ( .A1(n645), .A2(G73), .ZN(n639) );
  XOR2_X1 U730 ( .A(KEYINPUT2), .B(n639), .Z(n640) );
  NOR2_X1 U731 ( .A1(n641), .A2(n640), .ZN(n642) );
  XOR2_X1 U732 ( .A(KEYINPUT85), .B(n642), .Z(n644) );
  NAND2_X1 U733 ( .A1(n648), .A2(G48), .ZN(n643) );
  NAND2_X1 U734 ( .A1(n644), .A2(n643), .ZN(G305) );
  NAND2_X1 U735 ( .A1(n645), .A2(G72), .ZN(n646) );
  XNOR2_X1 U736 ( .A(KEYINPUT72), .B(n646), .ZN(n656) );
  NAND2_X1 U737 ( .A1(G60), .A2(n647), .ZN(n650) );
  NAND2_X1 U738 ( .A1(G47), .A2(n648), .ZN(n649) );
  NAND2_X1 U739 ( .A1(n650), .A2(n649), .ZN(n654) );
  NAND2_X1 U740 ( .A1(G85), .A2(n651), .ZN(n652) );
  XNOR2_X1 U741 ( .A(KEYINPUT71), .B(n652), .ZN(n653) );
  NOR2_X1 U742 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U743 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U744 ( .A(KEYINPUT73), .B(n657), .Z(G290) );
  XNOR2_X1 U745 ( .A(KEYINPUT86), .B(KEYINPUT19), .ZN(n658) );
  XOR2_X1 U746 ( .A(n658), .B(n666), .Z(n659) );
  XNOR2_X1 U747 ( .A(n659), .B(G288), .ZN(n662) );
  XNOR2_X1 U748 ( .A(n719), .B(G166), .ZN(n660) );
  XNOR2_X1 U749 ( .A(n660), .B(G305), .ZN(n661) );
  XNOR2_X1 U750 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U751 ( .A(n663), .B(G290), .ZN(n911) );
  XNOR2_X1 U752 ( .A(n664), .B(n911), .ZN(n665) );
  NAND2_X1 U753 ( .A1(n665), .A2(G868), .ZN(n669) );
  NAND2_X1 U754 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U755 ( .A1(n669), .A2(n668), .ZN(G295) );
  NAND2_X1 U756 ( .A1(G2084), .A2(G2078), .ZN(n670) );
  XNOR2_X1 U757 ( .A(n670), .B(KEYINPUT20), .ZN(n671) );
  XNOR2_X1 U758 ( .A(n671), .B(KEYINPUT87), .ZN(n672) );
  NAND2_X1 U759 ( .A1(n672), .A2(G2090), .ZN(n673) );
  XNOR2_X1 U760 ( .A(KEYINPUT21), .B(n673), .ZN(n674) );
  NAND2_X1 U761 ( .A1(n674), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U762 ( .A(KEYINPUT88), .B(G44), .ZN(n675) );
  XNOR2_X1 U763 ( .A(n675), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U764 ( .A1(G235), .A2(G236), .ZN(n676) );
  XNOR2_X1 U765 ( .A(n676), .B(KEYINPUT89), .ZN(n677) );
  NOR2_X1 U766 ( .A1(G237), .A2(n677), .ZN(n678) );
  XNOR2_X1 U767 ( .A(KEYINPUT90), .B(n678), .ZN(n679) );
  NAND2_X1 U768 ( .A1(n679), .A2(G108), .ZN(n843) );
  NAND2_X1 U769 ( .A1(n843), .A2(G567), .ZN(n684) );
  NOR2_X1 U770 ( .A1(G220), .A2(G219), .ZN(n680) );
  XOR2_X1 U771 ( .A(KEYINPUT22), .B(n680), .Z(n681) );
  NOR2_X1 U772 ( .A1(G218), .A2(n681), .ZN(n682) );
  NAND2_X1 U773 ( .A1(G96), .A2(n682), .ZN(n844) );
  NAND2_X1 U774 ( .A1(n844), .A2(G2106), .ZN(n683) );
  NAND2_X1 U775 ( .A1(n684), .A2(n683), .ZN(n845) );
  NAND2_X1 U776 ( .A1(G483), .A2(G661), .ZN(n685) );
  NOR2_X1 U777 ( .A1(n845), .A2(n685), .ZN(n842) );
  NAND2_X1 U778 ( .A1(n842), .A2(G36), .ZN(G176) );
  INV_X1 U779 ( .A(G166), .ZN(G303) );
  NAND2_X1 U780 ( .A1(G137), .A2(n896), .ZN(n687) );
  NAND2_X1 U781 ( .A1(G113), .A2(n891), .ZN(n686) );
  NAND2_X1 U782 ( .A1(n687), .A2(n686), .ZN(n696) );
  NAND2_X1 U783 ( .A1(G101), .A2(n897), .ZN(n688) );
  XNOR2_X1 U784 ( .A(n688), .B(KEYINPUT68), .ZN(n689) );
  XNOR2_X1 U785 ( .A(n689), .B(KEYINPUT23), .ZN(n693) );
  XNOR2_X1 U786 ( .A(KEYINPUT67), .B(n691), .ZN(n692) );
  NOR2_X1 U787 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U788 ( .A(n694), .B(KEYINPUT69), .ZN(n695) );
  XNOR2_X2 U789 ( .A(n697), .B(KEYINPUT64), .ZN(n702) );
  NAND2_X1 U790 ( .A1(n724), .A2(G1996), .ZN(n698) );
  XNOR2_X1 U791 ( .A(n698), .B(KEYINPUT26), .ZN(n701) );
  AND2_X1 U792 ( .A1(n702), .A2(G1341), .ZN(n699) );
  NOR2_X1 U793 ( .A1(n699), .A2(n966), .ZN(n700) );
  AND2_X1 U794 ( .A1(n701), .A2(n700), .ZN(n706) );
  NOR2_X1 U795 ( .A1(G2067), .A2(n702), .ZN(n704) );
  NOR2_X1 U796 ( .A1(G1348), .A2(n724), .ZN(n703) );
  NOR2_X1 U797 ( .A1(n704), .A2(n703), .ZN(n708) );
  NAND2_X1 U798 ( .A1(n707), .A2(n708), .ZN(n705) );
  NAND2_X1 U799 ( .A1(n706), .A2(n705), .ZN(n710) );
  NAND2_X1 U800 ( .A1(n710), .A2(n709), .ZN(n712) );
  XNOR2_X1 U801 ( .A(n712), .B(n711), .ZN(n718) );
  NAND2_X1 U802 ( .A1(G2072), .A2(n724), .ZN(n713) );
  XNOR2_X1 U803 ( .A(KEYINPUT27), .B(n713), .ZN(n716) );
  NAND2_X1 U804 ( .A1(n702), .A2(G1956), .ZN(n714) );
  NAND2_X1 U805 ( .A1(n720), .A2(n719), .ZN(n717) );
  NAND2_X1 U806 ( .A1(n718), .A2(n717), .ZN(n722) );
  NOR2_X1 U807 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U808 ( .A1(n722), .A2(n513), .ZN(n723) );
  XNOR2_X1 U809 ( .A(n723), .B(KEYINPUT29), .ZN(n728) );
  XOR2_X1 U810 ( .A(G2078), .B(KEYINPUT25), .Z(n986) );
  NOR2_X1 U811 ( .A1(n739), .A2(n986), .ZN(n726) );
  NOR2_X1 U812 ( .A1(G1961), .A2(n724), .ZN(n725) );
  NOR2_X1 U813 ( .A1(n726), .A2(n725), .ZN(n732) );
  NOR2_X1 U814 ( .A1(G301), .A2(n732), .ZN(n727) );
  NOR2_X1 U815 ( .A1(n728), .A2(n727), .ZN(n737) );
  NAND2_X1 U816 ( .A1(n702), .A2(G8), .ZN(n822) );
  NOR2_X1 U817 ( .A1(G1966), .A2(n822), .ZN(n750) );
  NOR2_X1 U818 ( .A1(n739), .A2(G2084), .ZN(n751) );
  NOR2_X1 U819 ( .A1(n750), .A2(n751), .ZN(n729) );
  NAND2_X1 U820 ( .A1(G8), .A2(n729), .ZN(n730) );
  XNOR2_X1 U821 ( .A(KEYINPUT30), .B(n730), .ZN(n731) );
  NOR2_X1 U822 ( .A1(G168), .A2(n731), .ZN(n734) );
  AND2_X1 U823 ( .A1(G301), .A2(n732), .ZN(n733) );
  NOR2_X1 U824 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U825 ( .A(n735), .B(KEYINPUT31), .ZN(n736) );
  NOR2_X2 U826 ( .A1(n737), .A2(n736), .ZN(n748) );
  AND2_X1 U827 ( .A1(G286), .A2(G8), .ZN(n738) );
  INV_X1 U828 ( .A(G8), .ZN(n744) );
  NOR2_X1 U829 ( .A1(n739), .A2(G2090), .ZN(n741) );
  NOR2_X1 U830 ( .A1(G1971), .A2(n822), .ZN(n740) );
  NOR2_X1 U831 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U832 ( .A1(n742), .A2(G303), .ZN(n743) );
  OR2_X1 U833 ( .A1(n744), .A2(n743), .ZN(n745) );
  INV_X1 U834 ( .A(KEYINPUT102), .ZN(n746) );
  XNOR2_X1 U835 ( .A(n748), .B(n747), .ZN(n749) );
  NOR2_X1 U836 ( .A1(n750), .A2(n749), .ZN(n753) );
  NAND2_X1 U837 ( .A1(G8), .A2(n751), .ZN(n752) );
  NAND2_X1 U838 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U839 ( .A1(n755), .A2(n754), .ZN(n816) );
  NOR2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n758) );
  NOR2_X1 U841 ( .A1(G1971), .A2(G303), .ZN(n756) );
  NOR2_X1 U842 ( .A1(n758), .A2(n756), .ZN(n962) );
  NAND2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n958) );
  NOR2_X1 U844 ( .A1(KEYINPUT33), .A2(n757), .ZN(n761) );
  NAND2_X1 U845 ( .A1(n758), .A2(KEYINPUT33), .ZN(n759) );
  NOR2_X1 U846 ( .A1(n822), .A2(n759), .ZN(n760) );
  XOR2_X1 U847 ( .A(G1981), .B(G305), .Z(n976) );
  INV_X1 U848 ( .A(KEYINPUT103), .ZN(n811) );
  XNOR2_X1 U849 ( .A(KEYINPUT92), .B(KEYINPUT34), .ZN(n765) );
  NAND2_X1 U850 ( .A1(G140), .A2(n896), .ZN(n763) );
  NAND2_X1 U851 ( .A1(G104), .A2(n897), .ZN(n762) );
  NAND2_X1 U852 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U853 ( .A(n765), .B(n764), .ZN(n771) );
  NAND2_X1 U854 ( .A1(G116), .A2(n891), .ZN(n766) );
  XOR2_X1 U855 ( .A(KEYINPUT93), .B(n766), .Z(n768) );
  NAND2_X1 U856 ( .A1(G128), .A2(n543), .ZN(n767) );
  NAND2_X1 U857 ( .A1(n768), .A2(n767), .ZN(n769) );
  XOR2_X1 U858 ( .A(KEYINPUT35), .B(n769), .Z(n770) );
  NOR2_X1 U859 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U860 ( .A(KEYINPUT36), .B(n772), .ZN(n905) );
  XNOR2_X1 U861 ( .A(KEYINPUT37), .B(G2067), .ZN(n799) );
  NAND2_X1 U862 ( .A1(n905), .A2(n799), .ZN(n938) );
  NAND2_X1 U863 ( .A1(G119), .A2(n543), .ZN(n774) );
  NAND2_X1 U864 ( .A1(G107), .A2(n891), .ZN(n773) );
  NAND2_X1 U865 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U866 ( .A(KEYINPUT94), .B(n775), .ZN(n780) );
  NAND2_X1 U867 ( .A1(G131), .A2(n896), .ZN(n777) );
  NAND2_X1 U868 ( .A1(G95), .A2(n897), .ZN(n776) );
  NAND2_X1 U869 ( .A1(n777), .A2(n776), .ZN(n778) );
  XOR2_X1 U870 ( .A(KEYINPUT95), .B(n778), .Z(n779) );
  NOR2_X1 U871 ( .A1(n780), .A2(n779), .ZN(n781) );
  XOR2_X1 U872 ( .A(KEYINPUT96), .B(n781), .Z(n888) );
  OR2_X1 U873 ( .A1(G1991), .A2(n888), .ZN(n937) );
  NOR2_X1 U874 ( .A1(G1986), .A2(G290), .ZN(n782) );
  XOR2_X1 U875 ( .A(n782), .B(KEYINPUT106), .Z(n783) );
  NAND2_X1 U876 ( .A1(n937), .A2(n783), .ZN(n795) );
  NOR2_X1 U877 ( .A1(n785), .A2(n784), .ZN(n806) );
  NAND2_X1 U878 ( .A1(G1991), .A2(n888), .ZN(n794) );
  NAND2_X1 U879 ( .A1(n896), .A2(G141), .ZN(n787) );
  NAND2_X1 U880 ( .A1(G129), .A2(n543), .ZN(n786) );
  NAND2_X1 U881 ( .A1(n787), .A2(n786), .ZN(n790) );
  NAND2_X1 U882 ( .A1(n897), .A2(G105), .ZN(n788) );
  XOR2_X1 U883 ( .A(KEYINPUT38), .B(n788), .Z(n789) );
  NOR2_X1 U884 ( .A1(n790), .A2(n789), .ZN(n792) );
  NAND2_X1 U885 ( .A1(G117), .A2(n891), .ZN(n791) );
  NAND2_X1 U886 ( .A1(n792), .A2(n791), .ZN(n884) );
  NAND2_X1 U887 ( .A1(G1996), .A2(n884), .ZN(n793) );
  NAND2_X1 U888 ( .A1(n794), .A2(n793), .ZN(n948) );
  NAND2_X1 U889 ( .A1(n806), .A2(n948), .ZN(n803) );
  NAND2_X1 U890 ( .A1(n795), .A2(n803), .ZN(n797) );
  NOR2_X1 U891 ( .A1(n884), .A2(G1996), .ZN(n796) );
  XNOR2_X1 U892 ( .A(n796), .B(KEYINPUT105), .ZN(n945) );
  NAND2_X1 U893 ( .A1(n797), .A2(n945), .ZN(n798) );
  XOR2_X1 U894 ( .A(KEYINPUT39), .B(n798), .Z(n800) );
  NOR2_X1 U895 ( .A1(n905), .A2(n799), .ZN(n936) );
  NAND2_X1 U896 ( .A1(n806), .A2(n936), .ZN(n804) );
  NAND2_X1 U897 ( .A1(n800), .A2(n804), .ZN(n801) );
  NAND2_X1 U898 ( .A1(n938), .A2(n801), .ZN(n802) );
  NAND2_X1 U899 ( .A1(n802), .A2(n806), .ZN(n824) );
  INV_X1 U900 ( .A(n824), .ZN(n810) );
  NAND2_X1 U901 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U902 ( .A(KEYINPUT97), .B(n805), .Z(n808) );
  XNOR2_X1 U903 ( .A(G1986), .B(G290), .ZN(n968) );
  AND2_X1 U904 ( .A1(n968), .A2(n806), .ZN(n807) );
  NOR2_X1 U905 ( .A1(n808), .A2(n807), .ZN(n809) );
  OR2_X1 U906 ( .A1(n810), .A2(n809), .ZN(n829) );
  AND2_X1 U907 ( .A1(n811), .A2(n829), .ZN(n812) );
  NAND2_X1 U908 ( .A1(n813), .A2(n812), .ZN(n835) );
  NOR2_X1 U909 ( .A1(G2090), .A2(G303), .ZN(n814) );
  NAND2_X1 U910 ( .A1(G8), .A2(n814), .ZN(n815) );
  NAND2_X1 U911 ( .A1(n816), .A2(n815), .ZN(n817) );
  NAND2_X1 U912 ( .A1(n817), .A2(n822), .ZN(n818) );
  XNOR2_X1 U913 ( .A(n818), .B(KEYINPUT104), .ZN(n823) );
  NOR2_X1 U914 ( .A1(G1981), .A2(G305), .ZN(n819) );
  XOR2_X1 U915 ( .A(n819), .B(KEYINPUT24), .Z(n820) );
  XNOR2_X1 U916 ( .A(KEYINPUT98), .B(n820), .ZN(n821) );
  AND2_X1 U917 ( .A1(n823), .A2(n532), .ZN(n825) );
  NAND2_X1 U918 ( .A1(n825), .A2(n824), .ZN(n828) );
  INV_X1 U919 ( .A(n828), .ZN(n826) );
  AND2_X1 U920 ( .A1(n976), .A2(n826), .ZN(n827) );
  NOR2_X1 U921 ( .A1(n828), .A2(KEYINPUT103), .ZN(n831) );
  INV_X1 U922 ( .A(n829), .ZN(n830) );
  NOR2_X1 U923 ( .A1(n831), .A2(n830), .ZN(n832) );
  NAND2_X1 U924 ( .A1(n833), .A2(n832), .ZN(n834) );
  NAND2_X1 U925 ( .A1(n835), .A2(n834), .ZN(n837) );
  XOR2_X1 U926 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n836) );
  XNOR2_X1 U927 ( .A(n837), .B(n836), .ZN(G329) );
  NAND2_X1 U928 ( .A1(n838), .A2(G2106), .ZN(n839) );
  XNOR2_X1 U929 ( .A(n839), .B(KEYINPUT108), .ZN(G217) );
  AND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n840) );
  NAND2_X1 U931 ( .A1(G661), .A2(n840), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n841) );
  NAND2_X1 U933 ( .A1(n842), .A2(n841), .ZN(G188) );
  NOR2_X1 U934 ( .A1(n844), .A2(n843), .ZN(G325) );
  XNOR2_X1 U935 ( .A(KEYINPUT109), .B(G325), .ZN(G261) );
  INV_X1 U937 ( .A(G108), .ZN(G238) );
  INV_X1 U938 ( .A(G96), .ZN(G221) );
  INV_X1 U939 ( .A(n845), .ZN(G319) );
  XNOR2_X1 U940 ( .A(G1981), .B(KEYINPUT112), .ZN(n855) );
  XOR2_X1 U941 ( .A(G1971), .B(G1956), .Z(n847) );
  XNOR2_X1 U942 ( .A(G1986), .B(G1966), .ZN(n846) );
  XNOR2_X1 U943 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U944 ( .A(G1976), .B(G1961), .Z(n849) );
  XNOR2_X1 U945 ( .A(G1996), .B(G1991), .ZN(n848) );
  XNOR2_X1 U946 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U947 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U948 ( .A(G2474), .B(KEYINPUT41), .ZN(n852) );
  XNOR2_X1 U949 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U950 ( .A(n855), .B(n854), .ZN(G229) );
  XOR2_X1 U951 ( .A(KEYINPUT111), .B(KEYINPUT110), .Z(n857) );
  XNOR2_X1 U952 ( .A(G2678), .B(KEYINPUT43), .ZN(n856) );
  XNOR2_X1 U953 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U954 ( .A(KEYINPUT42), .B(G2090), .Z(n859) );
  XNOR2_X1 U955 ( .A(G2067), .B(G2072), .ZN(n858) );
  XNOR2_X1 U956 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U957 ( .A(n861), .B(n860), .Z(n863) );
  XNOR2_X1 U958 ( .A(G2096), .B(G2100), .ZN(n862) );
  XNOR2_X1 U959 ( .A(n863), .B(n862), .ZN(n865) );
  XOR2_X1 U960 ( .A(G2084), .B(G2078), .Z(n864) );
  XNOR2_X1 U961 ( .A(n865), .B(n864), .ZN(G227) );
  NAND2_X1 U962 ( .A1(G100), .A2(n897), .ZN(n867) );
  NAND2_X1 U963 ( .A1(G112), .A2(n891), .ZN(n866) );
  NAND2_X1 U964 ( .A1(n867), .A2(n866), .ZN(n873) );
  NAND2_X1 U965 ( .A1(G124), .A2(n543), .ZN(n868) );
  XNOR2_X1 U966 ( .A(n868), .B(KEYINPUT44), .ZN(n870) );
  NAND2_X1 U967 ( .A1(G136), .A2(n896), .ZN(n869) );
  NAND2_X1 U968 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U969 ( .A(KEYINPUT113), .B(n871), .Z(n872) );
  NOR2_X1 U970 ( .A1(n873), .A2(n872), .ZN(G162) );
  NAND2_X1 U971 ( .A1(G139), .A2(n896), .ZN(n875) );
  NAND2_X1 U972 ( .A1(G103), .A2(n897), .ZN(n874) );
  NAND2_X1 U973 ( .A1(n875), .A2(n874), .ZN(n880) );
  NAND2_X1 U974 ( .A1(G127), .A2(n543), .ZN(n877) );
  NAND2_X1 U975 ( .A1(G115), .A2(n891), .ZN(n876) );
  NAND2_X1 U976 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U977 ( .A(KEYINPUT47), .B(n878), .Z(n879) );
  NOR2_X1 U978 ( .A1(n880), .A2(n879), .ZN(n931) );
  XOR2_X1 U979 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n882) );
  XNOR2_X1 U980 ( .A(KEYINPUT117), .B(KEYINPUT116), .ZN(n881) );
  XNOR2_X1 U981 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U982 ( .A(n931), .B(n883), .ZN(n886) );
  XNOR2_X1 U983 ( .A(n884), .B(G162), .ZN(n885) );
  XNOR2_X1 U984 ( .A(n886), .B(n885), .ZN(n887) );
  XOR2_X1 U985 ( .A(n887), .B(n940), .Z(n890) );
  XNOR2_X1 U986 ( .A(G164), .B(n888), .ZN(n889) );
  XNOR2_X1 U987 ( .A(n890), .B(n889), .ZN(n907) );
  NAND2_X1 U988 ( .A1(G118), .A2(n891), .ZN(n892) );
  XNOR2_X1 U989 ( .A(n892), .B(KEYINPUT114), .ZN(n894) );
  NAND2_X1 U990 ( .A1(G130), .A2(n543), .ZN(n893) );
  NAND2_X1 U991 ( .A1(n894), .A2(n893), .ZN(n895) );
  XNOR2_X1 U992 ( .A(n895), .B(KEYINPUT115), .ZN(n902) );
  NAND2_X1 U993 ( .A1(G142), .A2(n896), .ZN(n899) );
  NAND2_X1 U994 ( .A1(G106), .A2(n897), .ZN(n898) );
  NAND2_X1 U995 ( .A1(n899), .A2(n898), .ZN(n900) );
  XNOR2_X1 U996 ( .A(KEYINPUT45), .B(n900), .ZN(n901) );
  NAND2_X1 U997 ( .A1(n902), .A2(n901), .ZN(n903) );
  XNOR2_X1 U998 ( .A(n903), .B(G160), .ZN(n904) );
  XNOR2_X1 U999 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1000 ( .A(n907), .B(n906), .ZN(n908) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n908), .ZN(G395) );
  XOR2_X1 U1002 ( .A(KEYINPUT118), .B(G286), .Z(n910) );
  XNOR2_X1 U1003 ( .A(G171), .B(n971), .ZN(n909) );
  XNOR2_X1 U1004 ( .A(n910), .B(n909), .ZN(n913) );
  XNOR2_X1 U1005 ( .A(n966), .B(n911), .ZN(n912) );
  XNOR2_X1 U1006 ( .A(n913), .B(n912), .ZN(n914) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n914), .ZN(G397) );
  XOR2_X1 U1008 ( .A(G2451), .B(G2430), .Z(n916) );
  XNOR2_X1 U1009 ( .A(G2438), .B(G2443), .ZN(n915) );
  XNOR2_X1 U1010 ( .A(n916), .B(n915), .ZN(n922) );
  XOR2_X1 U1011 ( .A(G2435), .B(G2454), .Z(n918) );
  XNOR2_X1 U1012 ( .A(G1348), .B(G1341), .ZN(n917) );
  XNOR2_X1 U1013 ( .A(n918), .B(n917), .ZN(n920) );
  XOR2_X1 U1014 ( .A(G2446), .B(G2427), .Z(n919) );
  XNOR2_X1 U1015 ( .A(n920), .B(n919), .ZN(n921) );
  XOR2_X1 U1016 ( .A(n922), .B(n921), .Z(n923) );
  NAND2_X1 U1017 ( .A1(G14), .A2(n923), .ZN(n930) );
  NAND2_X1 U1018 ( .A1(G319), .A2(n930), .ZN(n927) );
  NOR2_X1 U1019 ( .A1(G229), .A2(G227), .ZN(n924) );
  XOR2_X1 U1020 ( .A(KEYINPUT49), .B(n924), .Z(n925) );
  XNOR2_X1 U1021 ( .A(n925), .B(KEYINPUT119), .ZN(n926) );
  NOR2_X1 U1022 ( .A1(n927), .A2(n926), .ZN(n929) );
  NOR2_X1 U1023 ( .A1(G395), .A2(G397), .ZN(n928) );
  NAND2_X1 U1024 ( .A1(n929), .A2(n928), .ZN(G225) );
  INV_X1 U1025 ( .A(G225), .ZN(G308) );
  INV_X1 U1026 ( .A(n930), .ZN(G401) );
  XOR2_X1 U1027 ( .A(G2072), .B(n931), .Z(n933) );
  XOR2_X1 U1028 ( .A(G164), .B(G2078), .Z(n932) );
  NOR2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1030 ( .A(KEYINPUT50), .B(n934), .Z(n935) );
  NOR2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n942) );
  NAND2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1034 ( .A1(n942), .A2(n941), .ZN(n952) );
  XNOR2_X1 U1035 ( .A(G2090), .B(G162), .ZN(n943) );
  XNOR2_X1 U1036 ( .A(n943), .B(KEYINPUT120), .ZN(n944) );
  NAND2_X1 U1037 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1038 ( .A(n946), .B(KEYINPUT51), .ZN(n950) );
  XOR2_X1 U1039 ( .A(G160), .B(G2084), .Z(n947) );
  NOR2_X1 U1040 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1041 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1042 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1043 ( .A(KEYINPUT52), .B(n953), .ZN(n955) );
  INV_X1 U1044 ( .A(KEYINPUT55), .ZN(n954) );
  NAND2_X1 U1045 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1046 ( .A1(n956), .A2(G29), .ZN(n1032) );
  XNOR2_X1 U1047 ( .A(KEYINPUT56), .B(G16), .ZN(n982) );
  NAND2_X1 U1048 ( .A1(G1971), .A2(G303), .ZN(n957) );
  NAND2_X1 U1049 ( .A1(n958), .A2(n957), .ZN(n960) );
  XNOR2_X1 U1050 ( .A(G1961), .B(G301), .ZN(n959) );
  NOR2_X1 U1051 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1052 ( .A1(n962), .A2(n961), .ZN(n965) );
  XOR2_X1 U1053 ( .A(G1956), .B(G299), .Z(n963) );
  XNOR2_X1 U1054 ( .A(KEYINPUT123), .B(n963), .ZN(n964) );
  NOR2_X1 U1055 ( .A1(n965), .A2(n964), .ZN(n970) );
  XNOR2_X1 U1056 ( .A(G1341), .B(n966), .ZN(n967) );
  NOR2_X1 U1057 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1058 ( .A1(n970), .A2(n969), .ZN(n974) );
  XOR2_X1 U1059 ( .A(n971), .B(G1348), .Z(n972) );
  XNOR2_X1 U1060 ( .A(KEYINPUT122), .B(n972), .ZN(n973) );
  NOR2_X1 U1061 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1062 ( .A(KEYINPUT124), .B(n975), .ZN(n980) );
  XNOR2_X1 U1063 ( .A(G1966), .B(G168), .ZN(n977) );
  NAND2_X1 U1064 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1065 ( .A(KEYINPUT57), .B(n978), .ZN(n979) );
  NAND2_X1 U1066 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1067 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1068 ( .A(n983), .B(KEYINPUT125), .ZN(n1029) );
  XNOR2_X1 U1069 ( .A(G2067), .B(G26), .ZN(n985) );
  XNOR2_X1 U1070 ( .A(G2072), .B(G33), .ZN(n984) );
  NOR2_X1 U1071 ( .A1(n985), .A2(n984), .ZN(n990) );
  XNOR2_X1 U1072 ( .A(G1996), .B(G32), .ZN(n988) );
  XNOR2_X1 U1073 ( .A(G27), .B(n986), .ZN(n987) );
  NOR2_X1 U1074 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1075 ( .A1(n990), .A2(n989), .ZN(n994) );
  XOR2_X1 U1076 ( .A(G25), .B(G1991), .Z(n991) );
  NAND2_X1 U1077 ( .A1(n991), .A2(G28), .ZN(n992) );
  XOR2_X1 U1078 ( .A(KEYINPUT121), .B(n992), .Z(n993) );
  NOR2_X1 U1079 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1080 ( .A(KEYINPUT53), .B(n995), .Z(n998) );
  XOR2_X1 U1081 ( .A(G34), .B(KEYINPUT54), .Z(n996) );
  XNOR2_X1 U1082 ( .A(G2084), .B(n996), .ZN(n997) );
  NAND2_X1 U1083 ( .A1(n998), .A2(n997), .ZN(n1000) );
  XNOR2_X1 U1084 ( .A(G35), .B(G2090), .ZN(n999) );
  NOR2_X1 U1085 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1086 ( .A(KEYINPUT55), .B(n1001), .Z(n1002) );
  NOR2_X1 U1087 ( .A1(G29), .A2(n1002), .ZN(n1026) );
  XNOR2_X1 U1088 ( .A(G1971), .B(G22), .ZN(n1004) );
  XNOR2_X1 U1089 ( .A(G1976), .B(G23), .ZN(n1003) );
  NOR2_X1 U1090 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1091 ( .A(KEYINPUT126), .B(n1005), .Z(n1007) );
  XNOR2_X1 U1092 ( .A(G1986), .B(G24), .ZN(n1006) );
  NOR2_X1 U1093 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1094 ( .A(KEYINPUT58), .B(n1008), .ZN(n1012) );
  XNOR2_X1 U1095 ( .A(G1966), .B(G21), .ZN(n1010) );
  XNOR2_X1 U1096 ( .A(G5), .B(G1961), .ZN(n1009) );
  NOR2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1022) );
  XOR2_X1 U1099 ( .A(G1348), .B(KEYINPUT59), .Z(n1013) );
  XNOR2_X1 U1100 ( .A(G4), .B(n1013), .ZN(n1015) );
  XNOR2_X1 U1101 ( .A(G20), .B(G1956), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1019) );
  XNOR2_X1 U1103 ( .A(G1981), .B(G6), .ZN(n1017) );
  XNOR2_X1 U1104 ( .A(G19), .B(G1341), .ZN(n1016) );
  NOR2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(KEYINPUT60), .B(n1020), .ZN(n1021) );
  NOR2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1109 ( .A(KEYINPUT61), .B(n1023), .Z(n1024) );
  NOR2_X1 U1110 ( .A1(G16), .A2(n1024), .ZN(n1025) );
  NOR2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1112 ( .A1(G11), .A2(n1027), .ZN(n1028) );
  NOR2_X1 U1113 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1114 ( .A(KEYINPUT127), .B(n1030), .Z(n1031) );
  NAND2_X1 U1115 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XOR2_X1 U1116 ( .A(KEYINPUT62), .B(n1033), .Z(G311) );
  INV_X1 U1117 ( .A(G311), .ZN(G150) );
endmodule

