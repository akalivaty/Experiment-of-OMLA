//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 0 0 1 0 1 1 0 1 0 1 0 1 0 0 0 1 0 0 1 0 0 1 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1265, new_n1266, new_n1267,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT0), .Z(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n209), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n203), .A2(G50), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n214), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G116), .A2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G50), .ZN(new_n221));
  INV_X1    g0021(.A(G226), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(G77), .B2(G244), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n225), .A2(new_n226), .A3(KEYINPUT66), .ZN(new_n227));
  INV_X1    g0027(.A(G238), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT65), .B(G68), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n224), .B(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(KEYINPUT66), .B1(new_n225), .B2(new_n226), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n211), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(KEYINPUT1), .ZN(new_n233));
  OR2_X1    g0033(.A1(new_n232), .A2(KEYINPUT1), .ZN(new_n234));
  NAND3_X1  g0034(.A1(new_n219), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n235), .B(KEYINPUT67), .Z(G361));
  XOR2_X1   g0036(.A(G238), .B(G244), .Z(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G226), .B(G232), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT69), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n250), .B(new_n251), .Z(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n215), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  OAI21_X1  g0056(.A(KEYINPUT70), .B1(new_n256), .B2(G20), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT70), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(new_n209), .A3(G33), .ZN(new_n259));
  AND2_X1   g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT8), .B(G58), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n263));
  INV_X1    g0063(.A(G150), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n263), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n255), .B1(new_n262), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G13), .ZN(new_n269));
  NOR3_X1   g0069(.A1(new_n269), .A2(new_n209), .A3(G1), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(new_n255), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n221), .B1(new_n208), .B2(G20), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n271), .A2(new_n272), .B1(new_n221), .B2(new_n270), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n268), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g0074(.A(new_n274), .B(KEYINPUT73), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT9), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT73), .ZN(new_n277));
  XNOR2_X1  g0077(.A(new_n274), .B(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT9), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT3), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n256), .ZN(new_n282));
  NAND2_X1  g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  AOI21_X1  g0083(.A(G1698), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G222), .ZN(new_n285));
  INV_X1    g0085(.A(G77), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n282), .A2(new_n283), .ZN(new_n287));
  INV_X1    g0087(.A(G223), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(G1698), .ZN(new_n289));
  OAI221_X1 g0089(.A(new_n285), .B1(new_n286), .B2(new_n287), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G41), .ZN(new_n293));
  INV_X1    g0093(.A(G45), .ZN(new_n294));
  AOI21_X1  g0094(.A(G1), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(G33), .A2(G41), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n296), .A2(G1), .A3(G13), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n295), .A2(new_n297), .A3(G274), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n291), .A2(new_n295), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n299), .B1(G226), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n292), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G200), .ZN(new_n303));
  INV_X1    g0103(.A(new_n302), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n304), .A2(G190), .B1(KEYINPUT74), .B2(KEYINPUT10), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n276), .A2(new_n280), .A3(new_n303), .A4(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(KEYINPUT74), .A2(KEYINPUT10), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n306), .B(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n274), .B1(new_n304), .B2(G169), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n302), .A2(G179), .ZN(new_n311));
  OR2_X1    g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n257), .A2(new_n259), .ZN(new_n313));
  INV_X1    g0113(.A(G87), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT15), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT15), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G87), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n313), .A2(new_n318), .B1(G20), .B2(G77), .ZN(new_n319));
  XNOR2_X1  g0119(.A(new_n261), .B(KEYINPUT71), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n319), .B1(new_n320), .B2(new_n266), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n255), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n271), .A2(KEYINPUT72), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n208), .A2(G20), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT72), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(new_n270), .B2(new_n255), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n323), .A2(G77), .A3(new_n324), .A4(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n269), .A2(G1), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G20), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n322), .B(new_n327), .C1(G77), .C2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G1698), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n287), .A2(G232), .A3(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G107), .ZN(new_n333));
  OAI221_X1 g0133(.A(new_n332), .B1(new_n333), .B2(new_n287), .C1(new_n289), .C2(new_n228), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n291), .ZN(new_n335));
  INV_X1    g0135(.A(G179), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n299), .B1(G244), .B2(new_n300), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n335), .A2(new_n337), .ZN(new_n339));
  INV_X1    g0139(.A(G169), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AND3_X1   g0141(.A1(new_n330), .A2(new_n338), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n339), .A2(G200), .ZN(new_n343));
  INV_X1    g0143(.A(G190), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n345), .A2(new_n330), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n342), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n309), .A2(new_n312), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n271), .ZN(new_n349));
  INV_X1    g0149(.A(new_n261), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n324), .ZN(new_n351));
  OAI22_X1  g0151(.A1(new_n349), .A2(new_n351), .B1(new_n329), .B2(new_n350), .ZN(new_n352));
  INV_X1    g0152(.A(new_n255), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT78), .ZN(new_n354));
  INV_X1    g0154(.A(G159), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n266), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n203), .B1(new_n229), .B2(new_n201), .ZN(new_n357));
  AOI211_X1 g0157(.A(new_n354), .B(new_n356), .C1(new_n357), .C2(G20), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n202), .A2(KEYINPUT65), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT65), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(G68), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n201), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n203), .ZN(new_n363));
  OAI21_X1  g0163(.A(G20), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n356), .ZN(new_n365));
  AOI21_X1  g0165(.A(KEYINPUT78), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n358), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT16), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT7), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n287), .B2(G20), .ZN(new_n370));
  AND2_X1   g0170(.A1(KEYINPUT3), .A2(G33), .ZN(new_n371));
  NOR2_X1   g0171(.A1(KEYINPUT3), .A2(G33), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n373), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n368), .B1(new_n375), .B2(G68), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n353), .B1(new_n367), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n360), .A2(G68), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n202), .A2(KEYINPUT65), .ZN(new_n379));
  OAI21_X1  g0179(.A(G58), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n209), .B1(new_n380), .B2(new_n203), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n354), .B1(new_n381), .B2(new_n356), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n364), .A2(KEYINPUT78), .A3(new_n365), .ZN(new_n383));
  INV_X1    g0183(.A(new_n229), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n375), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n382), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n368), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n352), .B1(new_n377), .B2(new_n387), .ZN(new_n388));
  OAI211_X1 g0188(.A(G223), .B(new_n331), .C1(new_n371), .C2(new_n372), .ZN(new_n389));
  OAI211_X1 g0189(.A(G226), .B(G1698), .C1(new_n371), .C2(new_n372), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n389), .B(new_n390), .C1(new_n256), .C2(new_n314), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n291), .ZN(new_n392));
  INV_X1    g0192(.A(G274), .ZN(new_n393));
  INV_X1    g0193(.A(new_n215), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n393), .B1(new_n394), .B2(new_n296), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n300), .A2(G232), .B1(new_n395), .B2(new_n295), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n392), .A2(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n397), .A2(new_n336), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n340), .B1(new_n392), .B2(new_n396), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT18), .B1(new_n388), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(G200), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n397), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(G190), .B2(new_n397), .ZN(new_n404));
  INV_X1    g0204(.A(new_n352), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT16), .B1(new_n367), .B2(new_n385), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n376), .A2(new_n382), .A3(new_n383), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n255), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n404), .B(new_n405), .C1(new_n406), .C2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT17), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n405), .B1(new_n406), .B2(new_n408), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT18), .ZN(new_n413));
  OR2_X1    g0213(.A1(new_n398), .A2(new_n399), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n377), .A2(new_n387), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n416), .A2(KEYINPUT17), .A3(new_n405), .A4(new_n404), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n401), .A2(new_n411), .A3(new_n415), .A4(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n229), .A2(G20), .ZN(new_n419));
  OAI221_X1 g0219(.A(new_n419), .B1(new_n221), .B2(new_n266), .C1(new_n260), .C2(new_n286), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n255), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT76), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT11), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT76), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n419), .B1(new_n221), .B2(new_n266), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n260), .A2(new_n286), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n424), .B(new_n255), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n422), .A2(new_n423), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n427), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n424), .B1(new_n420), .B2(new_n255), .ZN(new_n430));
  OAI21_X1  g0230(.A(KEYINPUT11), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n323), .A2(G68), .A3(new_n324), .A4(new_n326), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT12), .B1(new_n270), .B2(new_n202), .ZN(new_n433));
  INV_X1    g0233(.A(new_n419), .ZN(new_n434));
  AND2_X1   g0234(.A1(new_n328), .A2(KEYINPUT12), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n428), .A2(new_n431), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(KEYINPUT77), .A2(G169), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n284), .A2(G226), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n287), .A2(G232), .A3(G1698), .ZN(new_n441));
  NAND2_X1  g0241(.A1(G33), .A2(G97), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n291), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT13), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT75), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n298), .A2(new_n446), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n299), .A2(KEYINPUT75), .B1(new_n300), .B2(G238), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n444), .A2(new_n445), .A3(new_n447), .A4(new_n448), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n284), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n297), .B1(new_n450), .B2(new_n441), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n300), .A2(G238), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n395), .A2(KEYINPUT75), .A3(new_n295), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n452), .A2(new_n453), .A3(new_n447), .ZN(new_n454));
  OAI21_X1  g0254(.A(KEYINPUT13), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n439), .B1(new_n449), .B2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT14), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n449), .A2(new_n455), .A3(G179), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n460), .B1(new_n456), .B2(new_n457), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n438), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n449), .A2(new_n455), .A3(G190), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n402), .B1(new_n449), .B2(new_n455), .ZN(new_n464));
  OR3_X1    g0264(.A1(new_n438), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n348), .A2(new_n418), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(G116), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n254), .A2(new_n215), .B1(G20), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G33), .A2(G283), .ZN(new_n471));
  INV_X1    g0271(.A(G97), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n471), .B(new_n209), .C1(G33), .C2(new_n472), .ZN(new_n473));
  AND3_X1   g0273(.A1(new_n470), .A2(KEYINPUT20), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT20), .B1(new_n470), .B2(new_n473), .ZN(new_n475));
  OR2_X1    g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n256), .A2(G1), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n477), .A2(new_n469), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n323), .A2(new_n326), .A3(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(KEYINPUT84), .B1(new_n329), .B2(G116), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT84), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n270), .A2(new_n481), .A3(new_n469), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n476), .A2(new_n479), .A3(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT85), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n476), .A2(KEYINPUT85), .A3(new_n479), .A4(new_n483), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g0288(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n489));
  OAI21_X1  g0289(.A(KEYINPUT80), .B1(new_n489), .B2(G41), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT80), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT5), .ZN(new_n492));
  AND2_X1   g0292(.A1(new_n492), .A2(KEYINPUT79), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n492), .A2(KEYINPUT79), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n491), .B(new_n293), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n208), .A2(G45), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n496), .B1(new_n492), .B2(G41), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n490), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n498), .A2(G270), .A3(new_n297), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n490), .A2(new_n495), .A3(new_n395), .A4(new_n497), .ZN(new_n500));
  OAI211_X1 g0300(.A(G264), .B(G1698), .C1(new_n371), .C2(new_n372), .ZN(new_n501));
  OAI211_X1 g0301(.A(G257), .B(new_n331), .C1(new_n371), .C2(new_n372), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n282), .A2(G303), .A3(new_n283), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n291), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n499), .A2(new_n500), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G190), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n488), .B(new_n507), .C1(new_n402), .C2(new_n506), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n486), .A2(new_n487), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n505), .A2(new_n500), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n340), .B1(new_n510), .B2(new_n499), .ZN(new_n511));
  AOI21_X1  g0311(.A(KEYINPUT21), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n499), .A2(new_n500), .A3(new_n505), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n514), .A2(KEYINPUT21), .A3(G169), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n510), .A2(G179), .A3(new_n499), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT86), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n517), .A2(new_n518), .A3(new_n509), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n518), .B1(new_n517), .B2(new_n509), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n508), .B(new_n513), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT6), .ZN(new_n522));
  NOR3_X1   g0322(.A1(new_n522), .A2(new_n472), .A3(G107), .ZN(new_n523));
  XNOR2_X1  g0323(.A(G97), .B(G107), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n523), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  OAI22_X1  g0325(.A1(new_n525), .A2(new_n209), .B1(new_n286), .B2(new_n266), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n333), .B1(new_n370), .B2(new_n374), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n255), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n329), .A2(G97), .ZN(new_n529));
  NOR3_X1   g0329(.A1(new_n270), .A2(new_n255), .A3(new_n477), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n529), .B1(new_n530), .B2(G97), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n498), .A2(G257), .A3(new_n297), .ZN(new_n533));
  OAI211_X1 g0333(.A(G250), .B(G1698), .C1(new_n371), .C2(new_n372), .ZN(new_n534));
  OAI211_X1 g0334(.A(G244), .B(new_n331), .C1(new_n371), .C2(new_n372), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT4), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n471), .B(new_n534), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(KEYINPUT4), .B1(new_n284), .B2(G244), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n291), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n533), .A2(new_n539), .A3(new_n500), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n532), .B1(G200), .B2(new_n540), .ZN(new_n541));
  OR2_X1    g0341(.A1(new_n540), .A2(new_n344), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n533), .A2(new_n539), .A3(new_n336), .A4(new_n500), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n540), .A2(new_n340), .B1(new_n528), .B2(new_n531), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n541), .A2(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NOR3_X1   g0345(.A1(new_n256), .A2(new_n469), .A3(G20), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT23), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(new_n209), .B2(G107), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n333), .A2(KEYINPUT23), .A3(G20), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n546), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n209), .B(G87), .C1(new_n371), .C2(new_n372), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n551), .A2(KEYINPUT22), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n551), .A2(KEYINPUT22), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n550), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n554), .A2(KEYINPUT24), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT24), .ZN(new_n556));
  XNOR2_X1  g0356(.A(new_n551), .B(KEYINPUT22), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n556), .B1(new_n557), .B2(new_n550), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n255), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT25), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n329), .B2(G107), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n270), .A2(KEYINPUT25), .A3(new_n333), .ZN(new_n562));
  AOI22_X1  g0362(.A1(G107), .A2(new_n530), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n287), .A2(G257), .A3(G1698), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n287), .A2(G250), .A3(new_n331), .ZN(new_n566));
  XNOR2_X1  g0366(.A(KEYINPUT87), .B(G294), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n565), .B(new_n566), .C1(new_n256), .C2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n291), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n498), .A2(G264), .A3(new_n297), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n569), .A2(new_n570), .A3(G179), .A4(new_n500), .ZN(new_n571));
  OR2_X1    g0371(.A1(new_n571), .A2(KEYINPUT88), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n569), .A2(new_n570), .A3(new_n500), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n573), .A2(G169), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n571), .A2(KEYINPUT88), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n564), .B(new_n572), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n496), .A2(G274), .ZN(new_n577));
  AOI21_X1  g0377(.A(G250), .B1(new_n208), .B2(G45), .ZN(new_n578));
  NOR3_X1   g0378(.A1(new_n577), .A2(new_n291), .A3(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(G244), .B(G1698), .C1(new_n371), .C2(new_n372), .ZN(new_n580));
  OAI211_X1 g0380(.A(G238), .B(new_n331), .C1(new_n371), .C2(new_n372), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n580), .B(new_n581), .C1(new_n256), .C2(new_n469), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n579), .B1(new_n582), .B2(new_n291), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n583), .A2(new_n344), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n583), .A2(G200), .ZN(new_n585));
  OR2_X1    g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT19), .B1(new_n313), .B2(G97), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT19), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n209), .B1(new_n442), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n314), .A2(new_n472), .A3(new_n333), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n209), .B(G68), .C1(new_n371), .C2(new_n372), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n255), .B1(new_n587), .B2(new_n593), .ZN(new_n594));
  XNOR2_X1  g0394(.A(KEYINPUT15), .B(G87), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n270), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(KEYINPUT81), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT81), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n594), .A2(new_n599), .A3(new_n596), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n598), .A2(new_n600), .B1(G87), .B2(new_n530), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT82), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n318), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n595), .A2(KEYINPUT82), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT83), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(new_n606), .A3(new_n530), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n603), .A2(new_n604), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n353), .B(new_n329), .C1(G1), .C2(new_n256), .ZN(new_n609));
  OAI21_X1  g0409(.A(KEYINPUT83), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n594), .A2(new_n599), .A3(new_n596), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n599), .B1(new_n594), .B2(new_n596), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n583), .A2(G179), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(new_n340), .B2(new_n583), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n586), .A2(new_n601), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n573), .A2(G200), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n569), .A2(new_n570), .A3(G190), .A4(new_n500), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n559), .A2(new_n618), .A3(new_n563), .A4(new_n619), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n545), .A2(new_n576), .A3(new_n617), .A4(new_n620), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n468), .A2(new_n521), .A3(new_n621), .ZN(G372));
  NAND2_X1  g0422(.A1(new_n614), .A2(new_n616), .ZN(new_n623));
  OAI22_X1  g0423(.A1(new_n612), .A2(new_n613), .B1(new_n314), .B2(new_n609), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n584), .A2(new_n585), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n620), .B(new_n623), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n532), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n540), .A2(G200), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n542), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n544), .A2(new_n543), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n626), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n574), .A2(new_n575), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n554), .A2(KEYINPUT24), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n557), .A2(new_n556), .A3(new_n550), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n353), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n563), .ZN(new_n637));
  OAI22_X1  g0437(.A1(new_n636), .A2(new_n637), .B1(new_n571), .B2(KEYINPUT88), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n517), .A2(new_n509), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n513), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n632), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n623), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT26), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n607), .A2(new_n610), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n645), .B1(new_n598), .B2(new_n600), .ZN(new_n646));
  INV_X1    g0446(.A(new_n616), .ZN(new_n647));
  OAI22_X1  g0447(.A1(new_n646), .A2(new_n647), .B1(new_n624), .B2(new_n625), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n644), .B1(new_n648), .B2(new_n630), .ZN(new_n649));
  INV_X1    g0449(.A(new_n630), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n617), .A2(KEYINPUT26), .A3(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n643), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n642), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n467), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n312), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n401), .A2(new_n415), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n456), .A2(new_n457), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n658), .A2(new_n458), .A3(new_n460), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n342), .B1(new_n659), .B2(new_n438), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n465), .A2(new_n411), .A3(new_n417), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n657), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n655), .B1(new_n662), .B2(new_n309), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n654), .A2(new_n663), .ZN(G369));
  NAND2_X1  g0464(.A1(new_n328), .A2(new_n209), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(G213), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(G343), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n488), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n641), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n521), .B2(new_n672), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n674), .A2(G330), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n639), .A2(new_n670), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n670), .B1(new_n636), .B2(new_n637), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n620), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n676), .B1(new_n639), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n513), .B1(new_n519), .B2(new_n520), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n639), .A2(new_n678), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(new_n682), .A3(new_n671), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n639), .A2(new_n671), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n680), .A2(new_n686), .ZN(G399));
  NAND2_X1  g0487(.A1(new_n212), .A2(new_n293), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(new_n208), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n590), .A2(G116), .ZN(new_n691));
  AOI22_X1  g0491(.A1(new_n690), .A2(new_n691), .B1(new_n218), .B2(new_n689), .ZN(new_n692));
  XOR2_X1   g0492(.A(new_n692), .B(KEYINPUT28), .Z(new_n693));
  NAND3_X1  g0493(.A1(new_n569), .A2(new_n570), .A3(new_n583), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(KEYINPUT90), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT90), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n569), .A2(new_n570), .A3(new_n583), .A4(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n516), .A2(new_n540), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT30), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n698), .A2(new_n699), .A3(KEYINPUT30), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n583), .A2(G179), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n573), .A2(new_n540), .A3(new_n514), .A4(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  XOR2_X1   g0506(.A(KEYINPUT89), .B(KEYINPUT31), .Z(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n706), .A2(new_n670), .A3(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n705), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n710), .B1(new_n700), .B2(new_n701), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n671), .B1(new_n711), .B2(new_n703), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n709), .B1(KEYINPUT31), .B2(new_n712), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n521), .A2(new_n621), .A3(new_n670), .ZN(new_n714));
  OAI21_X1  g0514(.A(G330), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT91), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n513), .B(new_n576), .C1(new_n519), .C2(new_n520), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n632), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n652), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n717), .B1(new_n720), .B2(new_n671), .ZN(new_n721));
  AOI211_X1 g0521(.A(KEYINPUT91), .B(new_n670), .C1(new_n719), .C2(new_n652), .ZN(new_n722));
  OAI21_X1  g0522(.A(KEYINPUT29), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n670), .B1(new_n642), .B2(new_n652), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(KEYINPUT29), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n716), .B1(new_n723), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n693), .B1(new_n727), .B2(G1), .ZN(G364));
  NOR3_X1   g0528(.A1(new_n269), .A2(new_n294), .A3(G20), .ZN(new_n729));
  OR2_X1    g0529(.A1(new_n729), .A2(KEYINPUT92), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(KEYINPUT92), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n690), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n675), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(G330), .B2(new_n674), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n215), .B1(G20), .B2(new_n340), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT97), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(new_n209), .B2(G190), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n344), .A2(KEYINPUT97), .A3(G20), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n402), .A2(G179), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(G283), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(G303), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n743), .A2(G20), .A3(G190), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n209), .A2(new_n336), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n750), .A2(G190), .A3(G200), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(G311), .ZN(new_n753));
  OAI221_X1 g0553(.A(new_n373), .B1(new_n747), .B2(new_n748), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n741), .A2(new_n742), .A3(new_n336), .A4(new_n402), .ZN(new_n755));
  XOR2_X1   g0555(.A(new_n755), .B(KEYINPUT100), .Z(new_n756));
  AOI211_X1 g0556(.A(new_n746), .B(new_n754), .C1(G329), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n749), .A2(G200), .ZN(new_n758));
  OR2_X1    g0558(.A1(new_n758), .A2(KEYINPUT96), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(KEYINPUT96), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n759), .A2(new_n344), .A3(new_n760), .ZN(new_n761));
  XOR2_X1   g0561(.A(KEYINPUT33), .B(G317), .Z(new_n762));
  INV_X1    g0562(.A(G322), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n750), .A2(new_n344), .A3(G200), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n761), .A2(new_n762), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT101), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n344), .A2(G179), .A3(G200), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n209), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n567), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n759), .A2(G190), .A3(new_n760), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n770), .B1(new_n772), .B2(G326), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n773), .A2(KEYINPUT99), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(KEYINPUT99), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n757), .A2(new_n767), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n769), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G97), .ZN(new_n778));
  OAI221_X1 g0578(.A(new_n778), .B1(new_n333), .B2(new_n744), .C1(new_n761), .C2(new_n202), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(G50), .B2(new_n772), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n755), .A2(new_n355), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT32), .ZN(new_n782));
  AOI22_X1  g0582(.A1(G58), .A2(new_n764), .B1(new_n751), .B2(G77), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(KEYINPUT95), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n748), .A2(new_n314), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n373), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n784), .B1(KEYINPUT98), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(KEYINPUT98), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n788), .B1(KEYINPUT95), .B2(new_n783), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n780), .A2(new_n782), .A3(new_n787), .A4(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n739), .B1(new_n776), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G13), .A2(G33), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(G20), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n738), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n795), .B(KEYINPUT94), .Z(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n217), .A2(G45), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n212), .A2(new_n373), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n798), .B(new_n799), .C1(new_n249), .C2(G45), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n212), .A2(new_n287), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n801), .A2(new_n206), .B1(G116), .B2(new_n212), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT93), .Z(new_n803));
  OR2_X1    g0603(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n734), .B(new_n791), .C1(new_n797), .C2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n794), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n805), .B1(new_n674), .B2(new_n806), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n737), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(G396));
  NAND2_X1  g0609(.A1(new_n342), .A2(new_n671), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n346), .A2(new_n343), .B1(new_n330), .B2(new_n670), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n810), .B1(new_n811), .B2(new_n342), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n724), .B(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n735), .B1(new_n814), .B2(new_n715), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n715), .B2(new_n814), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n738), .A2(new_n792), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n734), .B1(new_n286), .B2(new_n817), .ZN(new_n818));
  AOI22_X1  g0618(.A1(G143), .A2(new_n764), .B1(new_n751), .B2(G159), .ZN(new_n819));
  INV_X1    g0619(.A(G137), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n819), .B1(new_n761), .B2(new_n264), .C1(new_n820), .C2(new_n771), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT34), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n744), .A2(new_n202), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n287), .B1(new_n748), .B2(new_n221), .C1(new_n769), .C2(new_n201), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n823), .B(new_n824), .C1(new_n756), .C2(G132), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n756), .A2(G311), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G116), .A2(new_n751), .B1(new_n764), .B2(G294), .ZN(new_n827));
  INV_X1    g0627(.A(new_n744), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(G87), .ZN(new_n829));
  INV_X1    g0629(.A(new_n748), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n287), .B1(new_n830), .B2(G107), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n827), .A2(new_n778), .A3(new_n829), .A4(new_n831), .ZN(new_n832));
  XOR2_X1   g0632(.A(KEYINPUT102), .B(G283), .Z(new_n833));
  OAI22_X1  g0633(.A1(new_n747), .A2(new_n771), .B1(new_n761), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n822), .A2(new_n825), .B1(new_n826), .B2(new_n835), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n818), .B1(new_n739), .B2(new_n836), .C1(new_n813), .C2(new_n793), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n816), .A2(new_n837), .ZN(G384));
  INV_X1    g0638(.A(new_n525), .ZN(new_n839));
  OR2_X1    g0639(.A1(new_n839), .A2(KEYINPUT35), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(KEYINPUT35), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n840), .A2(G116), .A3(new_n216), .A4(new_n841), .ZN(new_n842));
  XOR2_X1   g0642(.A(new_n842), .B(KEYINPUT36), .Z(new_n843));
  NAND3_X1  g0643(.A1(new_n380), .A2(new_n218), .A3(G77), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n221), .A2(G68), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n208), .B(G13), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n375), .A2(G68), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT16), .B1(new_n367), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n405), .B1(new_n849), .B2(new_n408), .ZN(new_n850));
  INV_X1    g0650(.A(new_n668), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n418), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n406), .A2(new_n408), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n854), .A2(new_n352), .B1(new_n414), .B2(new_n851), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n409), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT37), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n850), .B1(new_n414), .B2(new_n851), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n857), .B1(new_n388), .B2(new_n404), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n856), .A2(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n853), .A2(new_n860), .A3(KEYINPUT38), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT39), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT38), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n416), .A2(new_n405), .B1(new_n400), .B2(new_n668), .ZN(new_n865));
  OAI21_X1  g0665(.A(KEYINPUT37), .B1(new_n865), .B2(KEYINPUT103), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n856), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n855), .A2(KEYINPUT103), .A3(KEYINPUT37), .A4(new_n409), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n388), .A2(new_n668), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n418), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT104), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT104), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n418), .A2(new_n873), .A3(new_n870), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n869), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n863), .B1(new_n864), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n853), .A2(new_n860), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n864), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n862), .B1(new_n878), .B2(new_n861), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT105), .B1(new_n876), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n861), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT38), .B1(new_n853), .B2(new_n860), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT39), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT105), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n867), .A2(new_n868), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n873), .B1(new_n418), .B2(new_n870), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT38), .B1(new_n887), .B2(new_n874), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n883), .B(new_n884), .C1(new_n888), .C2(new_n863), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n880), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n659), .A2(new_n438), .A3(new_n671), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  OR2_X1    g0693(.A1(new_n811), .A2(new_n342), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n724), .A2(new_n894), .B1(new_n342), .B2(new_n671), .ZN(new_n895));
  NOR3_X1   g0695(.A1(new_n438), .A2(new_n463), .A3(new_n464), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n438), .B(new_n670), .C1(new_n659), .C2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n438), .A2(new_n670), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n462), .A2(new_n465), .A3(new_n898), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n895), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n878), .A2(new_n861), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n901), .A2(new_n902), .B1(new_n656), .B2(new_n668), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n893), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n723), .A2(new_n467), .A3(new_n726), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n663), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n904), .B(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n875), .A2(new_n864), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n861), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n812), .B1(new_n897), .B2(new_n899), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n706), .A2(KEYINPUT31), .A3(new_n670), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n708), .B2(new_n712), .ZN(new_n912));
  OAI211_X1 g0712(.A(KEYINPUT40), .B(new_n910), .C1(new_n912), .C2(new_n714), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n626), .A2(new_n639), .A3(new_n631), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n511), .A2(KEYINPUT21), .B1(new_n506), .B2(G179), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT86), .B1(new_n916), .B2(new_n488), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n517), .A2(new_n518), .A3(new_n509), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n512), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n915), .A2(new_n919), .A3(new_n508), .A4(new_n671), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n706), .A2(new_n670), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n707), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n920), .A2(new_n911), .A3(new_n922), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n923), .B(new_n910), .C1(new_n881), .C2(new_n882), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT40), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n909), .A2(new_n914), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n926), .A2(new_n467), .A3(new_n923), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(G330), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n926), .B1(new_n467), .B2(new_n923), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n907), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(G1), .B1(new_n269), .B2(G20), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n907), .A2(new_n930), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n847), .B1(new_n933), .B2(new_n934), .ZN(G367));
  INV_X1    g0735(.A(KEYINPUT106), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n617), .B1(new_n601), .B2(new_n671), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n643), .A2(new_n624), .A3(new_n670), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n919), .A2(new_n670), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n629), .B(new_n630), .C1(new_n627), .C2(new_n671), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n650), .A2(new_n670), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n940), .A2(KEYINPUT42), .A3(new_n682), .A4(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT42), .ZN(new_n945));
  INV_X1    g0745(.A(new_n943), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n945), .B1(new_n683), .B2(new_n946), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n630), .B1(new_n941), .B2(new_n576), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n949), .A2(new_n671), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n936), .B(new_n939), .C1(new_n948), .C2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n939), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n944), .A2(new_n947), .B1(new_n671), .B2(new_n949), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n952), .B1(new_n953), .B2(KEYINPUT106), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT43), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  AND3_X1   g0756(.A1(new_n951), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(KEYINPUT43), .B1(new_n951), .B2(new_n954), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n957), .A2(new_n958), .B1(new_n680), .B2(new_n946), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n680), .A2(new_n946), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n951), .A2(new_n954), .A3(new_n956), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n951), .A2(new_n954), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n960), .B(new_n961), .C1(new_n962), .C2(KEYINPUT43), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n959), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n688), .B(KEYINPUT41), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n674), .A2(G330), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n966), .B(new_n683), .C1(new_n679), .C2(new_n940), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n683), .B1(new_n940), .B2(new_n679), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n675), .A2(new_n968), .ZN(new_n969));
  AOI221_X4 g0769(.A(new_n716), .B1(new_n967), .B2(new_n969), .C1(new_n723), .C2(new_n726), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n683), .A2(new_n684), .A3(new_n943), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT45), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n683), .A2(KEYINPUT45), .A3(new_n684), .A4(new_n943), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n686), .B2(new_n943), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n685), .A2(new_n946), .A3(new_n976), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n975), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n680), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(KEYINPUT108), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT108), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n980), .A2(new_n984), .A3(new_n981), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n975), .A2(new_n978), .A3(new_n680), .A4(new_n979), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n970), .A2(new_n983), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n965), .B1(new_n987), .B2(new_n727), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n732), .A2(new_n208), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n964), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n797), .B1(new_n212), .B2(new_n595), .ZN(new_n992));
  AND3_X1   g0792(.A1(new_n244), .A2(new_n212), .A3(new_n373), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n735), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n744), .A2(new_n286), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n287), .B1(new_n201), .B2(new_n748), .C1(new_n752), .C2(new_n221), .ZN(new_n996));
  INV_X1    g0796(.A(new_n755), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n995), .B(new_n996), .C1(G137), .C2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n777), .A2(G68), .ZN(new_n999));
  INV_X1    g0799(.A(G143), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n999), .B1(new_n264), .B2(new_n765), .C1(new_n771), .C2(new_n1000), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n998), .B1(KEYINPUT109), .B2(new_n1001), .C1(new_n355), .C2(new_n761), .ZN(new_n1002));
  AND2_X1   g0802(.A1(new_n1001), .A2(KEYINPUT109), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n373), .B1(new_n765), .B2(new_n747), .C1(new_n752), .C2(new_n833), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(G317), .B2(new_n997), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n472), .B2(new_n744), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n748), .A2(new_n469), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1007), .A2(KEYINPUT46), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n1007), .A2(KEYINPUT46), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n1008), .B(new_n1009), .C1(G107), .C2(new_n777), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1010), .B1(new_n753), .B2(new_n771), .C1(new_n567), .C2(new_n761), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n1002), .A2(new_n1003), .B1(new_n1006), .B2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n1013));
  XNOR2_X1  g0813(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n994), .B1(new_n1014), .B2(new_n738), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n952), .A2(new_n794), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n991), .A2(new_n1017), .ZN(G387));
  INV_X1    g0818(.A(KEYINPUT29), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n545), .A2(new_n617), .A3(new_n620), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(new_n919), .B2(new_n576), .ZN(new_n1021));
  NOR3_X1   g0821(.A1(new_n648), .A2(new_n644), .A3(new_n630), .ZN(new_n1022));
  AOI21_X1  g0822(.A(KEYINPUT26), .B1(new_n617), .B2(new_n650), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n623), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n671), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(KEYINPUT91), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n720), .A2(new_n717), .A3(new_n671), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1019), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n715), .B1(new_n1028), .B2(new_n725), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n967), .A2(new_n969), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n727), .A2(new_n1030), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1032), .A2(new_n1033), .A3(new_n689), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n679), .A2(new_n806), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n801), .A2(new_n691), .B1(G107), .B2(new_n212), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n320), .A2(G50), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT50), .ZN(new_n1038));
  AOI21_X1  g0838(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1038), .A2(new_n691), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n799), .B1(new_n241), .B2(G45), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1036), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n735), .B1(new_n1042), .B2(new_n796), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n608), .A2(new_n769), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n287), .B1(new_n752), .B2(new_n202), .C1(new_n221), .C2(new_n765), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1044), .B(new_n1045), .C1(G97), .C2(new_n828), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n761), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(G159), .A2(new_n772), .B1(new_n1047), .B2(new_n350), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n830), .A2(G77), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n264), .B2(new_n755), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT111), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1046), .A2(new_n1048), .A3(new_n1051), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n769), .A2(new_n833), .B1(new_n748), .B2(new_n567), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G303), .A2(new_n751), .B1(new_n764), .B2(G317), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1054), .B1(new_n761), .B2(new_n753), .C1(new_n763), .C2(new_n771), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT48), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1053), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n1056), .B2(new_n1055), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT49), .Z(new_n1059));
  AOI21_X1  g0859(.A(new_n287), .B1(new_n997), .B2(G326), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n469), .B2(new_n744), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1052), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1043), .B1(new_n1062), .B2(new_n738), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n1030), .A2(new_n990), .B1(new_n1035), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1034), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT112), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1034), .A2(KEYINPUT112), .A3(new_n1064), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(new_n1068), .ZN(G393));
  AND2_X1   g0869(.A1(new_n982), .A2(new_n986), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n987), .B(new_n689), .C1(new_n970), .C2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n982), .A2(new_n986), .A3(new_n990), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n252), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n797), .B1(new_n472), .B2(new_n212), .C1(new_n1073), .C2(new_n799), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT113), .ZN(new_n1075));
  OR2_X1    g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1076), .A2(new_n735), .A3(new_n1077), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n772), .A2(G317), .B1(G311), .B2(new_n764), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT52), .ZN(new_n1080));
  INV_X1    g0880(.A(G294), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n373), .B1(new_n748), .B2(new_n833), .C1(new_n752), .C2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(G116), .B2(new_n777), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(G322), .A2(new_n997), .B1(new_n828), .B2(G107), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1083), .B(new_n1084), .C1(new_n747), .C2(new_n761), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n771), .A2(new_n264), .B1(new_n355), .B2(new_n765), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT51), .Z(new_n1087));
  OAI21_X1  g0887(.A(new_n287), .B1(new_n748), .B2(new_n229), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n769), .A2(new_n286), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n1088), .B(new_n1089), .C1(G87), .C2(new_n828), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n320), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1091), .A2(new_n751), .B1(new_n997), .B2(G143), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1090), .B(new_n1092), .C1(new_n221), .C2(new_n761), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n1080), .A2(new_n1085), .B1(new_n1087), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1078), .B1(new_n738), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n943), .B2(new_n806), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1072), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(KEYINPUT114), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT114), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1072), .A2(new_n1099), .A3(new_n1096), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1071), .A2(new_n1101), .ZN(G390));
  NAND3_X1  g0902(.A1(new_n1026), .A2(new_n1027), .A3(new_n810), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n894), .ZN(new_n1104));
  OAI211_X1 g0904(.A(G330), .B(new_n910), .C1(new_n713), .C2(new_n714), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT115), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT31), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n921), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n920), .A2(new_n709), .A3(new_n1109), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1110), .A2(KEYINPUT115), .A3(G330), .A4(new_n910), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1107), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n923), .A2(G330), .A3(new_n813), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n900), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1104), .A2(new_n1112), .A3(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n900), .B1(new_n715), .B2(new_n812), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n923), .A2(G330), .A3(new_n910), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n895), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1115), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n467), .A2(G330), .A3(new_n923), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n905), .A2(new_n663), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n891), .B1(new_n895), .B2(new_n900), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n880), .A2(new_n889), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n892), .B1(new_n908), .B2(new_n861), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n1104), .B2(new_n900), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n1126), .A2(new_n1128), .A3(new_n1112), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1117), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1124), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1117), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1126), .A2(new_n1128), .A3(new_n1112), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1103), .A2(new_n894), .B1(new_n900), .B2(new_n1113), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n1136), .A2(new_n1112), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n905), .A2(new_n663), .A3(new_n1122), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1134), .A2(new_n1135), .A3(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1131), .A2(new_n1140), .A3(new_n689), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n734), .B1(new_n261), .B2(new_n817), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(KEYINPUT54), .B(G143), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n752), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(G132), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n287), .B1(new_n765), .B2(new_n1145), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n1144), .B(new_n1146), .C1(G159), .C2(new_n777), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n756), .A2(G125), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n830), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT53), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n748), .B2(new_n264), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1149), .A2(new_n1151), .B1(G50), .B2(new_n828), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(G128), .A2(new_n772), .B1(new_n1047), .B2(G137), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1147), .A2(new_n1148), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT116), .ZN(new_n1155));
  OR2_X1    g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n765), .A2(new_n469), .B1(new_n752), .B2(new_n472), .ZN(new_n1157));
  NOR4_X1   g0957(.A1(new_n1157), .A2(new_n1089), .A3(new_n785), .A4(new_n287), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n823), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n756), .A2(G294), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G107), .A2(new_n1047), .B1(new_n772), .B2(G283), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n1156), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1142), .B1(new_n739), .B2(new_n1164), .C1(new_n890), .C2(new_n793), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT117), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1165), .B(new_n1166), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n990), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1141), .A2(new_n1167), .A3(new_n1169), .ZN(G378));
  AOI21_X1  g0970(.A(new_n1138), .B1(new_n1168), .B2(new_n1121), .ZN(new_n1171));
  OR2_X1    g0971(.A1(new_n306), .A2(new_n307), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n306), .A2(new_n307), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1172), .A2(new_n1173), .A3(new_n312), .ZN(new_n1174));
  XOR2_X1   g0974(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1175), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n309), .A2(new_n312), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n278), .A2(new_n851), .ZN(new_n1180));
  XOR2_X1   g0980(.A(new_n1180), .B(KEYINPUT119), .Z(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1176), .A2(new_n1178), .A3(new_n1181), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n926), .B2(G330), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n914), .B1(new_n888), .B2(new_n881), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n924), .A2(new_n925), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1187), .A2(new_n1185), .A3(new_n1188), .A4(G330), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n891), .B1(new_n880), .B2(new_n889), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n903), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n1186), .A2(new_n1190), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1187), .A2(new_n1188), .A3(G330), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1185), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n893), .A2(new_n1196), .A3(new_n903), .A4(new_n1189), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1193), .A2(new_n1197), .A3(KEYINPUT57), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1193), .A2(new_n1197), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(new_n1123), .B2(new_n1140), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n689), .B1(new_n1171), .B2(new_n1198), .C1(new_n1200), .C2(KEYINPUT57), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1193), .A2(new_n1197), .A3(new_n990), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n817), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n735), .B1(G50), .B2(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n287), .A2(G41), .ZN(new_n1205));
  AOI211_X1 g1005(.A(G50), .B(new_n1205), .C1(new_n256), .C2(new_n293), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(G97), .A2(new_n1047), .B1(new_n772), .B2(G116), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n764), .A2(G107), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1208), .A2(new_n999), .A3(new_n1049), .A4(new_n1205), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n605), .B2(new_n751), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n756), .A2(G283), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n744), .A2(new_n201), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT118), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1207), .A2(new_n1210), .A3(new_n1211), .A4(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT58), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1206), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n764), .A2(G128), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n748), .B2(new_n1143), .C1(new_n752), .C2(new_n820), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(G150), .B2(new_n777), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1219), .B1(new_n1145), .B2(new_n761), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(G125), .B2(new_n772), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1222), .A2(KEYINPUT59), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n256), .B(new_n293), .C1(new_n744), .C2(new_n355), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(G124), .B2(new_n997), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT59), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1225), .B1(new_n1221), .B2(new_n1226), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1216), .B1(new_n1215), .B2(new_n1214), .C1(new_n1223), .C2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1204), .B1(new_n1228), .B2(new_n738), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n1195), .B2(new_n793), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1202), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1201), .A2(new_n1232), .ZN(G375));
  NAND2_X1  g1033(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n965), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1234), .A2(new_n1124), .A3(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n900), .A2(new_n792), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n735), .B1(G68), .B2(new_n1203), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(new_n1238), .B(KEYINPUT120), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n771), .A2(new_n1145), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n373), .B1(new_n830), .B2(G159), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1241), .B1(new_n765), .B2(new_n820), .C1(new_n264), .C2(new_n752), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n1240), .B(new_n1242), .C1(G50), .C2(new_n777), .ZN(new_n1243));
  OR2_X1    g1043(.A1(new_n761), .A2(new_n1143), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n756), .A2(G128), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1243), .A2(new_n1213), .A3(new_n1244), .A4(new_n1245), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n756), .A2(G303), .B1(G97), .B2(new_n830), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(KEYINPUT121), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n469), .A2(new_n761), .B1(new_n771), .B2(new_n1081), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n287), .B1(new_n751), .B2(G107), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(new_n745), .B2(new_n765), .ZN(new_n1251));
  OR4_X1    g1051(.A1(new_n995), .A2(new_n1249), .A3(new_n1044), .A4(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1246), .B1(new_n1248), .B2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1239), .B1(new_n1253), .B2(new_n738), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n1121), .A2(new_n990), .B1(new_n1237), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1236), .A2(new_n1255), .ZN(G381));
  INV_X1    g1056(.A(G375), .ZN(new_n1257));
  INV_X1    g1057(.A(G378), .ZN(new_n1258));
  INV_X1    g1058(.A(G390), .ZN(new_n1259));
  INV_X1    g1059(.A(G384), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1067), .A2(new_n808), .A3(new_n1068), .ZN(new_n1262));
  NOR4_X1   g1062(.A1(new_n1261), .A2(G387), .A3(G381), .A4(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1257), .A2(new_n1258), .A3(new_n1263), .ZN(G407));
  NAND2_X1  g1064(.A1(new_n669), .A2(G213), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1257), .A2(new_n1258), .A3(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(G407), .A2(new_n1267), .A3(G213), .ZN(G409));
  NAND4_X1  g1068(.A1(new_n1138), .A2(new_n1115), .A3(KEYINPUT60), .A4(new_n1120), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1124), .A2(new_n689), .A3(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(KEYINPUT60), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1255), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n1260), .ZN(new_n1273));
  OAI211_X1 g1073(.A(G384), .B(new_n1255), .C1(new_n1270), .C2(new_n1271), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(KEYINPUT123), .ZN(new_n1277));
  INV_X1    g1077(.A(G2897), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1265), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT123), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1280), .B1(new_n1275), .B2(new_n1281), .ZN(new_n1282));
  AOI211_X1 g1082(.A(KEYINPUT123), .B(new_n1279), .C1(new_n1273), .C2(new_n1274), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1277), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1231), .A2(KEYINPUT122), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1140), .A2(new_n1123), .ZN(new_n1287));
  AND2_X1   g1087(.A1(new_n1193), .A2(new_n1197), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1287), .A2(new_n1235), .A3(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT122), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1202), .A2(new_n1290), .A3(new_n1230), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1286), .A2(new_n1289), .A3(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(new_n1258), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n689), .B1(new_n1171), .B2(new_n1198), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT57), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1295));
  OAI211_X1 g1095(.A(G378), .B(new_n1232), .C1(new_n1294), .C2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1293), .A2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1265), .ZN(new_n1298));
  AOI21_X1  g1098(.A(KEYINPUT61), .B1(new_n1285), .B2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT63), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1300), .B1(new_n1298), .B2(new_n1275), .ZN(new_n1301));
  AND3_X1   g1101(.A1(new_n991), .A2(new_n1017), .A3(G390), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(KEYINPUT126), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1259), .A2(KEYINPUT125), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT125), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(G390), .A2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1304), .A2(G387), .A3(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n991), .A2(new_n1017), .A3(G390), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT126), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1068), .ZN(new_n1311));
  AOI21_X1  g1111(.A(KEYINPUT112), .B1(new_n1034), .B2(new_n1064), .ZN(new_n1312));
  OAI21_X1  g1112(.A(G396), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1262), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1303), .A2(new_n1307), .A3(new_n1310), .A4(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n959), .A2(new_n963), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n985), .A2(new_n986), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n984), .B1(new_n980), .B2(new_n981), .ZN(new_n1318));
  NOR3_X1   g1118(.A1(new_n1317), .A2(new_n1033), .A3(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1235), .B1(new_n1319), .B2(new_n1029), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1316), .B1(new_n1320), .B2(new_n989), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1017), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1259), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(new_n1308), .ZN(new_n1324));
  AND2_X1   g1124(.A1(new_n1313), .A2(new_n1262), .ZN(new_n1325));
  AOI21_X1  g1125(.A(KEYINPUT124), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT124), .ZN(new_n1327));
  AOI211_X1 g1127(.A(new_n1327), .B(new_n1314), .C1(new_n1323), .C2(new_n1308), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1315), .B1(new_n1326), .B2(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1266), .B1(new_n1293), .B2(new_n1296), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1330), .A2(KEYINPUT63), .A3(new_n1276), .ZN(new_n1331));
  NAND4_X1  g1131(.A1(new_n1299), .A2(new_n1301), .A3(new_n1329), .A4(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT62), .ZN(new_n1333));
  AND3_X1   g1133(.A1(new_n1330), .A2(new_n1333), .A3(new_n1276), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT61), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1335), .B1(new_n1330), .B2(new_n1284), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1333), .B1(new_n1330), .B2(new_n1276), .ZN(new_n1337));
  NOR3_X1   g1137(.A1(new_n1334), .A2(new_n1336), .A3(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT127), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1329), .A2(new_n1339), .ZN(new_n1340));
  OAI211_X1 g1140(.A(KEYINPUT127), .B(new_n1315), .C1(new_n1326), .C2(new_n1328), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1332), .B1(new_n1338), .B2(new_n1342), .ZN(G405));
  NAND2_X1  g1143(.A1(G375), .A2(new_n1258), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1344), .A2(new_n1275), .A3(new_n1296), .ZN(new_n1345));
  AOI21_X1  g1145(.A(G378), .B1(new_n1201), .B2(new_n1232), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1296), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1276), .B1(new_n1346), .B2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1345), .A2(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(new_n1341), .ZN(new_n1350));
  AOI21_X1  g1150(.A(G390), .B1(new_n991), .B2(new_n1017), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1325), .B1(new_n1302), .B2(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1352), .A2(new_n1327), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1324), .A2(KEYINPUT124), .A3(new_n1325), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1353), .A2(new_n1354), .ZN(new_n1355));
  AOI21_X1  g1155(.A(KEYINPUT127), .B1(new_n1355), .B2(new_n1315), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1349), .B1(new_n1350), .B2(new_n1356), .ZN(new_n1357));
  NAND4_X1  g1157(.A1(new_n1340), .A2(new_n1341), .A3(new_n1348), .A4(new_n1345), .ZN(new_n1358));
  AND2_X1   g1158(.A1(new_n1357), .A2(new_n1358), .ZN(G402));
endmodule


