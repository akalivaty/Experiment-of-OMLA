

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X2 U557 ( .A1(n701), .A2(n692), .ZN(n693) );
  XNOR2_X1 U558 ( .A(KEYINPUT17), .B(n525), .ZN(n899) );
  OR2_X1 U559 ( .A1(n663), .A2(n789), .ZN(n662) );
  NAND2_X1 U560 ( .A1(n764), .A2(n611), .ZN(n641) );
  XOR2_X1 U561 ( .A(KEYINPUT14), .B(n638), .Z(n522) );
  AND2_X1 U562 ( .A1(G8), .A2(n734), .ZN(n523) );
  INV_X1 U563 ( .A(G8), .ZN(n690) );
  OR2_X1 U564 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U565 ( .A1(n696), .A2(n695), .ZN(n697) );
  OR2_X1 U566 ( .A1(n706), .A2(n705), .ZN(n716) );
  INV_X1 U567 ( .A(n985), .ZN(n723) );
  NAND2_X1 U568 ( .A1(n724), .A2(n723), .ZN(n725) );
  OR2_X1 U569 ( .A1(n735), .A2(n523), .ZN(n737) );
  NAND2_X1 U570 ( .A1(G8), .A2(n708), .ZN(n736) );
  XNOR2_X1 U571 ( .A(n631), .B(KEYINPUT74), .ZN(n632) );
  XNOR2_X1 U572 ( .A(n633), .B(n632), .ZN(n635) );
  INV_X1 U573 ( .A(G651), .ZN(n539) );
  NOR2_X1 U574 ( .A1(n639), .A2(n522), .ZN(n640) );
  NOR2_X1 U575 ( .A1(G2105), .A2(n530), .ZN(n898) );
  XNOR2_X1 U576 ( .A(KEYINPUT70), .B(n536), .ZN(n813) );
  NOR2_X1 U577 ( .A1(G2104), .A2(G2105), .ZN(n524) );
  XOR2_X1 U578 ( .A(KEYINPUT66), .B(n524), .Z(n525) );
  NAND2_X1 U579 ( .A1(G138), .A2(n899), .ZN(n528) );
  INV_X1 U580 ( .A(G2104), .ZN(n530) );
  NAND2_X1 U581 ( .A1(G102), .A2(n898), .ZN(n526) );
  XOR2_X1 U582 ( .A(KEYINPUT89), .B(n526), .Z(n527) );
  NAND2_X1 U583 ( .A1(n528), .A2(n527), .ZN(n534) );
  INV_X1 U584 ( .A(G2105), .ZN(n529) );
  NOR2_X1 U585 ( .A1(G2104), .A2(n529), .ZN(n903) );
  NAND2_X1 U586 ( .A1(G126), .A2(n903), .ZN(n532) );
  NOR2_X1 U587 ( .A1(n530), .A2(n529), .ZN(n904) );
  NAND2_X1 U588 ( .A1(G114), .A2(n904), .ZN(n531) );
  NAND2_X1 U589 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U590 ( .A1(n534), .A2(n533), .ZN(G164) );
  XOR2_X1 U591 ( .A(G543), .B(KEYINPUT0), .Z(n579) );
  NOR2_X1 U592 ( .A1(G651), .A2(n579), .ZN(n809) );
  NAND2_X1 U593 ( .A1(G48), .A2(n809), .ZN(n538) );
  NOR2_X1 U594 ( .A1(G543), .A2(n539), .ZN(n535) );
  XOR2_X1 U595 ( .A(KEYINPUT1), .B(n535), .Z(n536) );
  NAND2_X1 U596 ( .A1(G61), .A2(n813), .ZN(n537) );
  NAND2_X1 U597 ( .A1(n538), .A2(n537), .ZN(n543) );
  OR2_X1 U598 ( .A1(n539), .A2(n579), .ZN(n540) );
  XNOR2_X1 U599 ( .A(KEYINPUT69), .B(n540), .ZN(n806) );
  NAND2_X1 U600 ( .A1(n806), .A2(G73), .ZN(n541) );
  XOR2_X1 U601 ( .A(KEYINPUT2), .B(n541), .Z(n542) );
  NOR2_X1 U602 ( .A1(n543), .A2(n542), .ZN(n546) );
  NOR2_X1 U603 ( .A1(G651), .A2(G543), .ZN(n544) );
  XOR2_X2 U604 ( .A(KEYINPUT65), .B(n544), .Z(n805) );
  NAND2_X1 U605 ( .A1(n805), .A2(G86), .ZN(n545) );
  NAND2_X1 U606 ( .A1(n546), .A2(n545), .ZN(G305) );
  NAND2_X1 U607 ( .A1(G90), .A2(n805), .ZN(n548) );
  NAND2_X1 U608 ( .A1(G77), .A2(n806), .ZN(n547) );
  NAND2_X1 U609 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U610 ( .A(KEYINPUT9), .B(n549), .ZN(n554) );
  NAND2_X1 U611 ( .A1(G52), .A2(n809), .ZN(n551) );
  NAND2_X1 U612 ( .A1(G64), .A2(n813), .ZN(n550) );
  NAND2_X1 U613 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U614 ( .A(KEYINPUT72), .B(n552), .Z(n553) );
  NAND2_X1 U615 ( .A1(n554), .A2(n553), .ZN(G301) );
  NAND2_X1 U616 ( .A1(n809), .A2(G51), .ZN(n555) );
  XNOR2_X1 U617 ( .A(n555), .B(KEYINPUT80), .ZN(n557) );
  NAND2_X1 U618 ( .A1(G63), .A2(n813), .ZN(n556) );
  NAND2_X1 U619 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U620 ( .A(KEYINPUT6), .B(n558), .ZN(n567) );
  NAND2_X1 U621 ( .A1(G76), .A2(n806), .ZN(n563) );
  XOR2_X1 U622 ( .A(KEYINPUT4), .B(KEYINPUT78), .Z(n560) );
  NAND2_X1 U623 ( .A1(G89), .A2(n805), .ZN(n559) );
  XNOR2_X1 U624 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U625 ( .A(KEYINPUT77), .B(n561), .ZN(n562) );
  NAND2_X1 U626 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U627 ( .A(n564), .B(KEYINPUT5), .ZN(n565) );
  XNOR2_X1 U628 ( .A(n565), .B(KEYINPUT79), .ZN(n566) );
  NOR2_X1 U629 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U630 ( .A(KEYINPUT7), .B(n568), .Z(G168) );
  XOR2_X1 U631 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U632 ( .A1(G88), .A2(n805), .ZN(n570) );
  NAND2_X1 U633 ( .A1(G75), .A2(n806), .ZN(n569) );
  NAND2_X1 U634 ( .A1(n570), .A2(n569), .ZN(n574) );
  NAND2_X1 U635 ( .A1(G50), .A2(n809), .ZN(n572) );
  NAND2_X1 U636 ( .A1(G62), .A2(n813), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U638 ( .A1(n574), .A2(n573), .ZN(G166) );
  INV_X1 U639 ( .A(G166), .ZN(G303) );
  NAND2_X1 U640 ( .A1(G49), .A2(n809), .ZN(n576) );
  NAND2_X1 U641 ( .A1(G74), .A2(G651), .ZN(n575) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U643 ( .A1(n813), .A2(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n578), .B(KEYINPUT84), .ZN(n581) );
  NAND2_X1 U645 ( .A1(G87), .A2(n579), .ZN(n580) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(G288) );
  NAND2_X1 U647 ( .A1(n805), .A2(G85), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n582), .B(KEYINPUT68), .ZN(n584) );
  NAND2_X1 U649 ( .A1(G72), .A2(n806), .ZN(n583) );
  NAND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(n587) );
  NAND2_X1 U651 ( .A1(G47), .A2(n809), .ZN(n585) );
  XNOR2_X1 U652 ( .A(KEYINPUT71), .B(n585), .ZN(n586) );
  NOR2_X1 U653 ( .A1(n587), .A2(n586), .ZN(n589) );
  NAND2_X1 U654 ( .A1(G60), .A2(n813), .ZN(n588) );
  NAND2_X1 U655 ( .A1(n589), .A2(n588), .ZN(G290) );
  NAND2_X1 U656 ( .A1(G131), .A2(n899), .ZN(n592) );
  NAND2_X1 U657 ( .A1(G107), .A2(n904), .ZN(n590) );
  XOR2_X1 U658 ( .A(KEYINPUT93), .B(n590), .Z(n591) );
  NAND2_X1 U659 ( .A1(n592), .A2(n591), .ZN(n596) );
  NAND2_X1 U660 ( .A1(G95), .A2(n898), .ZN(n594) );
  NAND2_X1 U661 ( .A1(G119), .A2(n903), .ZN(n593) );
  NAND2_X1 U662 ( .A1(n594), .A2(n593), .ZN(n595) );
  OR2_X1 U663 ( .A1(n596), .A2(n595), .ZN(n895) );
  AND2_X1 U664 ( .A1(n895), .A2(G1991), .ZN(n605) );
  NAND2_X1 U665 ( .A1(n904), .A2(G117), .ZN(n598) );
  NAND2_X1 U666 ( .A1(G141), .A2(n899), .ZN(n597) );
  NAND2_X1 U667 ( .A1(n598), .A2(n597), .ZN(n601) );
  NAND2_X1 U668 ( .A1(n898), .A2(G105), .ZN(n599) );
  XOR2_X1 U669 ( .A(KEYINPUT38), .B(n599), .Z(n600) );
  NOR2_X1 U670 ( .A1(n601), .A2(n600), .ZN(n603) );
  NAND2_X1 U671 ( .A1(n903), .A2(G129), .ZN(n602) );
  NAND2_X1 U672 ( .A1(n603), .A2(n602), .ZN(n880) );
  AND2_X1 U673 ( .A1(n880), .A2(G1996), .ZN(n604) );
  NOR2_X1 U674 ( .A1(n605), .A2(n604), .ZN(n947) );
  NOR2_X1 U675 ( .A1(G164), .A2(G1384), .ZN(n642) );
  NAND2_X1 U676 ( .A1(G137), .A2(n899), .ZN(n607) );
  NAND2_X1 U677 ( .A1(n904), .A2(G113), .ZN(n606) );
  NAND2_X1 U678 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U679 ( .A(n608), .B(KEYINPUT67), .ZN(n764) );
  NAND2_X1 U680 ( .A1(G101), .A2(n898), .ZN(n609) );
  XOR2_X1 U681 ( .A(KEYINPUT23), .B(n609), .Z(n765) );
  AND2_X1 U682 ( .A1(G40), .A2(n765), .ZN(n610) );
  NAND2_X1 U683 ( .A1(G125), .A2(n903), .ZN(n763) );
  AND2_X1 U684 ( .A1(n610), .A2(n763), .ZN(n611) );
  NOR2_X1 U685 ( .A1(n642), .A2(n641), .ZN(n758) );
  INV_X1 U686 ( .A(n758), .ZN(n612) );
  NOR2_X1 U687 ( .A1(n947), .A2(n612), .ZN(n750) );
  INV_X1 U688 ( .A(n750), .ZN(n626) );
  XNOR2_X1 U689 ( .A(G2067), .B(KEYINPUT37), .ZN(n756) );
  XNOR2_X1 U690 ( .A(KEYINPUT36), .B(KEYINPUT92), .ZN(n624) );
  NAND2_X1 U691 ( .A1(n904), .A2(G116), .ZN(n613) );
  XOR2_X1 U692 ( .A(KEYINPUT91), .B(n613), .Z(n615) );
  NAND2_X1 U693 ( .A1(n903), .A2(G128), .ZN(n614) );
  NAND2_X1 U694 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U695 ( .A(KEYINPUT35), .B(n616), .ZN(n622) );
  NAND2_X1 U696 ( .A1(G104), .A2(n898), .ZN(n618) );
  NAND2_X1 U697 ( .A1(G140), .A2(n899), .ZN(n617) );
  NAND2_X1 U698 ( .A1(n618), .A2(n617), .ZN(n620) );
  XOR2_X1 U699 ( .A(KEYINPUT34), .B(KEYINPUT90), .Z(n619) );
  XNOR2_X1 U700 ( .A(n620), .B(n619), .ZN(n621) );
  NAND2_X1 U701 ( .A1(n622), .A2(n621), .ZN(n623) );
  XOR2_X1 U702 ( .A(n624), .B(n623), .Z(n912) );
  NOR2_X1 U703 ( .A1(n756), .A2(n912), .ZN(n754) );
  NAND2_X1 U704 ( .A1(n758), .A2(n754), .ZN(n625) );
  NAND2_X1 U705 ( .A1(n626), .A2(n625), .ZN(n743) );
  INV_X1 U706 ( .A(n641), .ZN(n627) );
  NAND2_X2 U707 ( .A1(n642), .A2(n627), .ZN(n708) );
  NOR2_X1 U708 ( .A1(G1981), .A2(G305), .ZN(n628) );
  XOR2_X1 U709 ( .A(n628), .B(KEYINPUT24), .Z(n629) );
  NOR2_X1 U710 ( .A1(n736), .A2(n629), .ZN(n741) );
  NOR2_X1 U711 ( .A1(G2084), .A2(n708), .ZN(n691) );
  NAND2_X1 U712 ( .A1(G8), .A2(n691), .ZN(n630) );
  XNOR2_X1 U713 ( .A(KEYINPUT94), .B(n630), .ZN(n703) );
  NOR2_X1 U714 ( .A1(G1966), .A2(n736), .ZN(n701) );
  NAND2_X1 U715 ( .A1(G81), .A2(n805), .ZN(n633) );
  XOR2_X1 U716 ( .A(KEYINPUT12), .B(KEYINPUT75), .Z(n631) );
  NAND2_X1 U717 ( .A1(n806), .A2(G68), .ZN(n634) );
  NAND2_X1 U718 ( .A1(n635), .A2(n634), .ZN(n637) );
  INV_X1 U719 ( .A(KEYINPUT13), .ZN(n636) );
  XNOR2_X1 U720 ( .A(n637), .B(n636), .ZN(n639) );
  NAND2_X1 U721 ( .A1(G56), .A2(n813), .ZN(n638) );
  XNOR2_X1 U722 ( .A(n640), .B(KEYINPUT76), .ZN(n782) );
  NAND2_X1 U723 ( .A1(n809), .A2(G43), .ZN(n781) );
  NAND2_X1 U724 ( .A1(n782), .A2(n781), .ZN(n649) );
  INV_X1 U725 ( .A(G1996), .ZN(n958) );
  NOR2_X1 U726 ( .A1(n641), .A2(n958), .ZN(n643) );
  AND2_X1 U727 ( .A1(n643), .A2(n642), .ZN(n645) );
  XOR2_X1 U728 ( .A(KEYINPUT26), .B(KEYINPUT96), .Z(n644) );
  XNOR2_X1 U729 ( .A(n645), .B(n644), .ZN(n647) );
  NAND2_X1 U730 ( .A1(n708), .A2(G1341), .ZN(n646) );
  NAND2_X1 U731 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U732 ( .A1(n649), .A2(n648), .ZN(n651) );
  INV_X1 U733 ( .A(KEYINPUT64), .ZN(n650) );
  XNOR2_X1 U734 ( .A(n651), .B(n650), .ZN(n663) );
  NAND2_X1 U735 ( .A1(G54), .A2(n809), .ZN(n653) );
  NAND2_X1 U736 ( .A1(G66), .A2(n813), .ZN(n652) );
  NAND2_X1 U737 ( .A1(n653), .A2(n652), .ZN(n657) );
  NAND2_X1 U738 ( .A1(G92), .A2(n805), .ZN(n655) );
  NAND2_X1 U739 ( .A1(G79), .A2(n806), .ZN(n654) );
  NAND2_X1 U740 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U741 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U742 ( .A(n658), .B(KEYINPUT15), .ZN(n789) );
  INV_X1 U743 ( .A(n708), .ZN(n683) );
  NOR2_X1 U744 ( .A1(n683), .A2(G1348), .ZN(n660) );
  NOR2_X1 U745 ( .A1(G2067), .A2(n708), .ZN(n659) );
  NOR2_X1 U746 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U747 ( .A1(n662), .A2(n661), .ZN(n665) );
  NAND2_X1 U748 ( .A1(n663), .A2(n789), .ZN(n664) );
  NAND2_X1 U749 ( .A1(n665), .A2(n664), .ZN(n676) );
  NAND2_X1 U750 ( .A1(G53), .A2(n809), .ZN(n667) );
  NAND2_X1 U751 ( .A1(G65), .A2(n813), .ZN(n666) );
  NAND2_X1 U752 ( .A1(n667), .A2(n666), .ZN(n671) );
  NAND2_X1 U753 ( .A1(G91), .A2(n805), .ZN(n669) );
  NAND2_X1 U754 ( .A1(G78), .A2(n806), .ZN(n668) );
  NAND2_X1 U755 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U756 ( .A1(n671), .A2(n670), .ZN(n990) );
  NAND2_X1 U757 ( .A1(n683), .A2(G2072), .ZN(n672) );
  XNOR2_X1 U758 ( .A(n672), .B(KEYINPUT27), .ZN(n674) );
  INV_X1 U759 ( .A(G1956), .ZN(n1016) );
  NOR2_X1 U760 ( .A1(n1016), .A2(n683), .ZN(n673) );
  NOR2_X1 U761 ( .A1(n674), .A2(n673), .ZN(n677) );
  NAND2_X1 U762 ( .A1(n990), .A2(n677), .ZN(n675) );
  NAND2_X1 U763 ( .A1(n676), .A2(n675), .ZN(n681) );
  NOR2_X1 U764 ( .A1(n990), .A2(n677), .ZN(n679) );
  XNOR2_X1 U765 ( .A(KEYINPUT95), .B(KEYINPUT28), .ZN(n678) );
  XNOR2_X1 U766 ( .A(n679), .B(n678), .ZN(n680) );
  NAND2_X1 U767 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U768 ( .A(n682), .B(KEYINPUT29), .ZN(n687) );
  NAND2_X1 U769 ( .A1(G1961), .A2(n708), .ZN(n685) );
  XOR2_X1 U770 ( .A(KEYINPUT25), .B(G2078), .Z(n959) );
  NAND2_X1 U771 ( .A1(n683), .A2(n959), .ZN(n684) );
  NAND2_X1 U772 ( .A1(n685), .A2(n684), .ZN(n688) );
  NOR2_X1 U773 ( .A1(G301), .A2(n688), .ZN(n686) );
  NOR2_X1 U774 ( .A1(n687), .A2(n686), .ZN(n700) );
  NAND2_X1 U775 ( .A1(G301), .A2(n688), .ZN(n689) );
  XNOR2_X1 U776 ( .A(n689), .B(KEYINPUT97), .ZN(n696) );
  XNOR2_X1 U777 ( .A(KEYINPUT30), .B(n693), .ZN(n694) );
  NOR2_X1 U778 ( .A1(n694), .A2(G168), .ZN(n695) );
  XNOR2_X1 U779 ( .A(KEYINPUT98), .B(n697), .ZN(n698) );
  XNOR2_X1 U780 ( .A(KEYINPUT31), .B(n698), .ZN(n699) );
  NOR2_X1 U781 ( .A1(n700), .A2(n699), .ZN(n706) );
  NOR2_X1 U782 ( .A1(n701), .A2(n706), .ZN(n702) );
  NAND2_X1 U783 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U784 ( .A(KEYINPUT99), .B(n704), .ZN(n719) );
  NAND2_X1 U785 ( .A1(G286), .A2(G8), .ZN(n705) );
  NOR2_X1 U786 ( .A1(G1971), .A2(n736), .ZN(n707) );
  XNOR2_X1 U787 ( .A(n707), .B(KEYINPUT100), .ZN(n710) );
  NOR2_X1 U788 ( .A1(n708), .A2(G2090), .ZN(n709) );
  NOR2_X1 U789 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U790 ( .A(n711), .B(KEYINPUT101), .ZN(n712) );
  NOR2_X1 U791 ( .A1(G166), .A2(n712), .ZN(n713) );
  XOR2_X1 U792 ( .A(KEYINPUT102), .B(n713), .Z(n714) );
  OR2_X1 U793 ( .A1(n690), .A2(n714), .ZN(n715) );
  NAND2_X1 U794 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U795 ( .A(KEYINPUT32), .B(n717), .ZN(n718) );
  NOR2_X1 U796 ( .A1(n719), .A2(n718), .ZN(n735) );
  NOR2_X1 U797 ( .A1(G1971), .A2(G303), .ZN(n720) );
  XNOR2_X1 U798 ( .A(n720), .B(KEYINPUT103), .ZN(n722) );
  INV_X1 U799 ( .A(KEYINPUT33), .ZN(n721) );
  AND2_X1 U800 ( .A1(n722), .A2(n721), .ZN(n724) );
  NOR2_X1 U801 ( .A1(G1976), .A2(G288), .ZN(n985) );
  OR2_X1 U802 ( .A1(n735), .A2(n725), .ZN(n733) );
  NAND2_X1 U803 ( .A1(G1976), .A2(G288), .ZN(n982) );
  INV_X1 U804 ( .A(n982), .ZN(n726) );
  NOR2_X1 U805 ( .A1(n726), .A2(n736), .ZN(n727) );
  NOR2_X1 U806 ( .A1(KEYINPUT33), .A2(n727), .ZN(n730) );
  NAND2_X1 U807 ( .A1(n985), .A2(KEYINPUT33), .ZN(n728) );
  NOR2_X1 U808 ( .A1(n728), .A2(n736), .ZN(n729) );
  NOR2_X1 U809 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U810 ( .A(G1981), .B(G305), .Z(n986) );
  AND2_X1 U811 ( .A1(n731), .A2(n986), .ZN(n732) );
  NAND2_X1 U812 ( .A1(n733), .A2(n732), .ZN(n739) );
  NOR2_X1 U813 ( .A1(G2090), .A2(G303), .ZN(n734) );
  NAND2_X1 U814 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U815 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U816 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U817 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U818 ( .A(n744), .B(KEYINPUT104), .ZN(n746) );
  XNOR2_X1 U819 ( .A(G1986), .B(G290), .ZN(n996) );
  NAND2_X1 U820 ( .A1(n996), .A2(n758), .ZN(n745) );
  NAND2_X1 U821 ( .A1(n746), .A2(n745), .ZN(n761) );
  NOR2_X1 U822 ( .A1(G1996), .A2(n880), .ZN(n942) );
  NOR2_X1 U823 ( .A1(G1986), .A2(G290), .ZN(n748) );
  NOR2_X1 U824 ( .A1(G1991), .A2(n895), .ZN(n747) );
  XOR2_X1 U825 ( .A(KEYINPUT105), .B(n747), .Z(n948) );
  NOR2_X1 U826 ( .A1(n748), .A2(n948), .ZN(n749) );
  NOR2_X1 U827 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U828 ( .A(n751), .B(KEYINPUT106), .ZN(n752) );
  NOR2_X1 U829 ( .A1(n942), .A2(n752), .ZN(n753) );
  XNOR2_X1 U830 ( .A(n753), .B(KEYINPUT39), .ZN(n755) );
  INV_X1 U831 ( .A(n754), .ZN(n930) );
  NAND2_X1 U832 ( .A1(n755), .A2(n930), .ZN(n757) );
  NAND2_X1 U833 ( .A1(n912), .A2(n756), .ZN(n936) );
  NAND2_X1 U834 ( .A1(n757), .A2(n936), .ZN(n759) );
  NAND2_X1 U835 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U836 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U837 ( .A(n762), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U838 ( .A1(n764), .A2(n763), .ZN(n766) );
  AND2_X1 U839 ( .A1(n766), .A2(n765), .ZN(G160) );
  XNOR2_X1 U840 ( .A(G2454), .B(G2443), .ZN(n776) );
  XOR2_X1 U841 ( .A(G2430), .B(KEYINPUT108), .Z(n768) );
  XNOR2_X1 U842 ( .A(G2446), .B(KEYINPUT107), .ZN(n767) );
  XNOR2_X1 U843 ( .A(n768), .B(n767), .ZN(n772) );
  XOR2_X1 U844 ( .A(G2451), .B(G2427), .Z(n770) );
  XNOR2_X1 U845 ( .A(G1348), .B(G1341), .ZN(n769) );
  XNOR2_X1 U846 ( .A(n770), .B(n769), .ZN(n771) );
  XOR2_X1 U847 ( .A(n772), .B(n771), .Z(n774) );
  XNOR2_X1 U848 ( .A(G2435), .B(G2438), .ZN(n773) );
  XNOR2_X1 U849 ( .A(n774), .B(n773), .ZN(n775) );
  XNOR2_X1 U850 ( .A(n776), .B(n775), .ZN(n777) );
  AND2_X1 U851 ( .A1(n777), .A2(G14), .ZN(G401) );
  AND2_X1 U852 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U853 ( .A(G132), .ZN(G219) );
  INV_X1 U854 ( .A(G82), .ZN(G220) );
  INV_X1 U855 ( .A(G57), .ZN(G237) );
  INV_X1 U856 ( .A(G108), .ZN(G238) );
  INV_X1 U857 ( .A(G120), .ZN(G236) );
  NAND2_X1 U858 ( .A1(G7), .A2(G661), .ZN(n778) );
  XNOR2_X1 U859 ( .A(n778), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U860 ( .A(G223), .ZN(n846) );
  NAND2_X1 U861 ( .A1(n846), .A2(G567), .ZN(n779) );
  XNOR2_X1 U862 ( .A(n779), .B(KEYINPUT73), .ZN(n780) );
  XNOR2_X1 U863 ( .A(KEYINPUT11), .B(n780), .ZN(G234) );
  AND2_X1 U864 ( .A1(n782), .A2(n781), .ZN(n792) );
  NAND2_X1 U865 ( .A1(n792), .A2(G860), .ZN(G153) );
  NAND2_X1 U866 ( .A1(G868), .A2(G301), .ZN(n784) );
  INV_X1 U867 ( .A(G868), .ZN(n827) );
  NAND2_X1 U868 ( .A1(n789), .A2(n827), .ZN(n783) );
  NAND2_X1 U869 ( .A1(n784), .A2(n783), .ZN(G284) );
  INV_X1 U870 ( .A(n990), .ZN(G299) );
  NOR2_X1 U871 ( .A1(G286), .A2(n827), .ZN(n786) );
  NOR2_X1 U872 ( .A1(G868), .A2(G299), .ZN(n785) );
  NOR2_X1 U873 ( .A1(n786), .A2(n785), .ZN(G297) );
  INV_X1 U874 ( .A(G559), .ZN(n787) );
  NOR2_X1 U875 ( .A1(G860), .A2(n787), .ZN(n788) );
  XNOR2_X1 U876 ( .A(KEYINPUT81), .B(n788), .ZN(n790) );
  INV_X1 U877 ( .A(n789), .ZN(n981) );
  NAND2_X1 U878 ( .A1(n790), .A2(n981), .ZN(n791) );
  XNOR2_X1 U879 ( .A(n791), .B(KEYINPUT16), .ZN(G148) );
  INV_X1 U880 ( .A(n792), .ZN(n999) );
  NOR2_X1 U881 ( .A1(G868), .A2(n999), .ZN(n795) );
  NAND2_X1 U882 ( .A1(G868), .A2(n981), .ZN(n793) );
  NOR2_X1 U883 ( .A1(G559), .A2(n793), .ZN(n794) );
  NOR2_X1 U884 ( .A1(n795), .A2(n794), .ZN(G282) );
  NAND2_X1 U885 ( .A1(n903), .A2(G123), .ZN(n796) );
  XNOR2_X1 U886 ( .A(n796), .B(KEYINPUT18), .ZN(n798) );
  NAND2_X1 U887 ( .A1(G111), .A2(n904), .ZN(n797) );
  NAND2_X1 U888 ( .A1(n798), .A2(n797), .ZN(n802) );
  NAND2_X1 U889 ( .A1(G99), .A2(n898), .ZN(n800) );
  NAND2_X1 U890 ( .A1(G135), .A2(n899), .ZN(n799) );
  NAND2_X1 U891 ( .A1(n800), .A2(n799), .ZN(n801) );
  NOR2_X1 U892 ( .A1(n802), .A2(n801), .ZN(n945) );
  XOR2_X1 U893 ( .A(n945), .B(G2096), .Z(n803) );
  NOR2_X1 U894 ( .A1(G2100), .A2(n803), .ZN(n804) );
  XOR2_X1 U895 ( .A(KEYINPUT82), .B(n804), .Z(G156) );
  NAND2_X1 U896 ( .A1(G93), .A2(n805), .ZN(n808) );
  NAND2_X1 U897 ( .A1(G80), .A2(n806), .ZN(n807) );
  NAND2_X1 U898 ( .A1(n808), .A2(n807), .ZN(n812) );
  NAND2_X1 U899 ( .A1(G55), .A2(n809), .ZN(n810) );
  XNOR2_X1 U900 ( .A(KEYINPUT83), .B(n810), .ZN(n811) );
  NOR2_X1 U901 ( .A1(n812), .A2(n811), .ZN(n815) );
  NAND2_X1 U902 ( .A1(G67), .A2(n813), .ZN(n814) );
  NAND2_X1 U903 ( .A1(n815), .A2(n814), .ZN(n828) );
  NAND2_X1 U904 ( .A1(n981), .A2(G559), .ZN(n825) );
  XNOR2_X1 U905 ( .A(n999), .B(n825), .ZN(n816) );
  NOR2_X1 U906 ( .A1(G860), .A2(n816), .ZN(n817) );
  XOR2_X1 U907 ( .A(n828), .B(n817), .Z(G145) );
  XOR2_X1 U908 ( .A(KEYINPUT19), .B(KEYINPUT85), .Z(n818) );
  XNOR2_X1 U909 ( .A(G288), .B(n818), .ZN(n819) );
  XNOR2_X1 U910 ( .A(G166), .B(n819), .ZN(n821) );
  XNOR2_X1 U911 ( .A(G290), .B(n990), .ZN(n820) );
  XNOR2_X1 U912 ( .A(n821), .B(n820), .ZN(n822) );
  XNOR2_X1 U913 ( .A(n822), .B(G305), .ZN(n823) );
  XNOR2_X1 U914 ( .A(n823), .B(n828), .ZN(n824) );
  XNOR2_X1 U915 ( .A(n824), .B(n999), .ZN(n917) );
  XOR2_X1 U916 ( .A(n917), .B(n825), .Z(n826) );
  NAND2_X1 U917 ( .A1(G868), .A2(n826), .ZN(n830) );
  NAND2_X1 U918 ( .A1(n828), .A2(n827), .ZN(n829) );
  NAND2_X1 U919 ( .A1(n830), .A2(n829), .ZN(G295) );
  NAND2_X1 U920 ( .A1(G2084), .A2(G2078), .ZN(n832) );
  XOR2_X1 U921 ( .A(KEYINPUT20), .B(KEYINPUT86), .Z(n831) );
  XNOR2_X1 U922 ( .A(n832), .B(n831), .ZN(n833) );
  NAND2_X1 U923 ( .A1(G2090), .A2(n833), .ZN(n834) );
  XNOR2_X1 U924 ( .A(KEYINPUT21), .B(n834), .ZN(n835) );
  NAND2_X1 U925 ( .A1(n835), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U926 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U927 ( .A1(G483), .A2(G661), .ZN(n844) );
  NOR2_X1 U928 ( .A1(G236), .A2(G238), .ZN(n836) );
  NAND2_X1 U929 ( .A1(G69), .A2(n836), .ZN(n837) );
  NOR2_X1 U930 ( .A1(n837), .A2(G237), .ZN(n838) );
  XNOR2_X1 U931 ( .A(n838), .B(KEYINPUT87), .ZN(n927) );
  NAND2_X1 U932 ( .A1(n927), .A2(G567), .ZN(n843) );
  NOR2_X1 U933 ( .A1(G220), .A2(G219), .ZN(n839) );
  XOR2_X1 U934 ( .A(KEYINPUT22), .B(n839), .Z(n840) );
  NOR2_X1 U935 ( .A1(G218), .A2(n840), .ZN(n841) );
  NAND2_X1 U936 ( .A1(G96), .A2(n841), .ZN(n928) );
  NAND2_X1 U937 ( .A1(n928), .A2(G2106), .ZN(n842) );
  NAND2_X1 U938 ( .A1(n843), .A2(n842), .ZN(n929) );
  NOR2_X1 U939 ( .A1(n844), .A2(n929), .ZN(n845) );
  XNOR2_X1 U940 ( .A(n845), .B(KEYINPUT88), .ZN(n851) );
  NAND2_X1 U941 ( .A1(G36), .A2(n851), .ZN(G176) );
  NAND2_X1 U942 ( .A1(G2106), .A2(n846), .ZN(G217) );
  NAND2_X1 U943 ( .A1(G15), .A2(G2), .ZN(n848) );
  INV_X1 U944 ( .A(G661), .ZN(n847) );
  NOR2_X1 U945 ( .A1(n848), .A2(n847), .ZN(n849) );
  XNOR2_X1 U946 ( .A(n849), .B(KEYINPUT109), .ZN(G259) );
  NAND2_X1 U947 ( .A1(G3), .A2(G1), .ZN(n850) );
  NAND2_X1 U948 ( .A1(n851), .A2(n850), .ZN(G188) );
  XOR2_X1 U949 ( .A(G1976), .B(G1956), .Z(n853) );
  XNOR2_X1 U950 ( .A(G1996), .B(G1991), .ZN(n852) );
  XNOR2_X1 U951 ( .A(n853), .B(n852), .ZN(n863) );
  XOR2_X1 U952 ( .A(KEYINPUT112), .B(KEYINPUT111), .Z(n855) );
  XNOR2_X1 U953 ( .A(G1986), .B(G2474), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U955 ( .A(G1981), .B(G1971), .Z(n857) );
  XNOR2_X1 U956 ( .A(G1966), .B(G1961), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U958 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U959 ( .A(KEYINPUT41), .B(KEYINPUT113), .ZN(n860) );
  XNOR2_X1 U960 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U961 ( .A(n863), .B(n862), .Z(G229) );
  XOR2_X1 U962 ( .A(G2096), .B(KEYINPUT43), .Z(n865) );
  XNOR2_X1 U963 ( .A(G2090), .B(G2678), .ZN(n864) );
  XNOR2_X1 U964 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U965 ( .A(n866), .B(KEYINPUT110), .Z(n868) );
  XNOR2_X1 U966 ( .A(G2067), .B(G2072), .ZN(n867) );
  XNOR2_X1 U967 ( .A(n868), .B(n867), .ZN(n872) );
  XOR2_X1 U968 ( .A(KEYINPUT42), .B(G2100), .Z(n870) );
  XNOR2_X1 U969 ( .A(G2084), .B(G2078), .ZN(n869) );
  XNOR2_X1 U970 ( .A(n870), .B(n869), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n872), .B(n871), .ZN(G227) );
  NAND2_X1 U972 ( .A1(n903), .A2(G124), .ZN(n873) );
  XNOR2_X1 U973 ( .A(n873), .B(KEYINPUT44), .ZN(n875) );
  NAND2_X1 U974 ( .A1(G112), .A2(n904), .ZN(n874) );
  NAND2_X1 U975 ( .A1(n875), .A2(n874), .ZN(n879) );
  NAND2_X1 U976 ( .A1(G100), .A2(n898), .ZN(n877) );
  NAND2_X1 U977 ( .A1(G136), .A2(n899), .ZN(n876) );
  NAND2_X1 U978 ( .A1(n877), .A2(n876), .ZN(n878) );
  NOR2_X1 U979 ( .A1(n879), .A2(n878), .ZN(G162) );
  XOR2_X1 U980 ( .A(G162), .B(n945), .Z(n882) );
  XOR2_X1 U981 ( .A(G164), .B(n880), .Z(n881) );
  XNOR2_X1 U982 ( .A(n882), .B(n881), .ZN(n886) );
  XOR2_X1 U983 ( .A(KEYINPUT48), .B(KEYINPUT116), .Z(n884) );
  XNOR2_X1 U984 ( .A(KEYINPUT117), .B(KEYINPUT46), .ZN(n883) );
  XNOR2_X1 U985 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U986 ( .A(n886), .B(n885), .Z(n897) );
  NAND2_X1 U987 ( .A1(G103), .A2(n898), .ZN(n888) );
  NAND2_X1 U988 ( .A1(G139), .A2(n899), .ZN(n887) );
  NAND2_X1 U989 ( .A1(n888), .A2(n887), .ZN(n894) );
  NAND2_X1 U990 ( .A1(G127), .A2(n903), .ZN(n890) );
  NAND2_X1 U991 ( .A1(G115), .A2(n904), .ZN(n889) );
  NAND2_X1 U992 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U993 ( .A(KEYINPUT115), .B(n891), .ZN(n892) );
  XNOR2_X1 U994 ( .A(KEYINPUT47), .B(n892), .ZN(n893) );
  NOR2_X1 U995 ( .A1(n894), .A2(n893), .ZN(n932) );
  XOR2_X1 U996 ( .A(n895), .B(n932), .Z(n896) );
  XNOR2_X1 U997 ( .A(n897), .B(n896), .ZN(n914) );
  NAND2_X1 U998 ( .A1(G106), .A2(n898), .ZN(n901) );
  NAND2_X1 U999 ( .A1(G142), .A2(n899), .ZN(n900) );
  NAND2_X1 U1000 ( .A1(n901), .A2(n900), .ZN(n902) );
  XNOR2_X1 U1001 ( .A(n902), .B(KEYINPUT45), .ZN(n909) );
  NAND2_X1 U1002 ( .A1(G130), .A2(n903), .ZN(n906) );
  NAND2_X1 U1003 ( .A1(G118), .A2(n904), .ZN(n905) );
  NAND2_X1 U1004 ( .A1(n906), .A2(n905), .ZN(n907) );
  XOR2_X1 U1005 ( .A(KEYINPUT114), .B(n907), .Z(n908) );
  NAND2_X1 U1006 ( .A1(n909), .A2(n908), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(n910), .B(G160), .ZN(n911) );
  XOR2_X1 U1008 ( .A(n912), .B(n911), .Z(n913) );
  XNOR2_X1 U1009 ( .A(n914), .B(n913), .ZN(n915) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n915), .ZN(G395) );
  INV_X1 U1011 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U1012 ( .A(G171), .B(n981), .ZN(n916) );
  XNOR2_X1 U1013 ( .A(n916), .B(G286), .ZN(n918) );
  XNOR2_X1 U1014 ( .A(n918), .B(n917), .ZN(n919) );
  NOR2_X1 U1015 ( .A1(G37), .A2(n919), .ZN(G397) );
  NOR2_X1 U1016 ( .A1(G229), .A2(G227), .ZN(n920) );
  XOR2_X1 U1017 ( .A(KEYINPUT49), .B(n920), .Z(n923) );
  NOR2_X1 U1018 ( .A1(G401), .A2(n929), .ZN(n921) );
  XNOR2_X1 U1019 ( .A(KEYINPUT118), .B(n921), .ZN(n922) );
  NAND2_X1 U1020 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1021 ( .A(KEYINPUT119), .B(n924), .ZN(n926) );
  NOR2_X1 U1022 ( .A1(G395), .A2(G397), .ZN(n925) );
  NAND2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(G225) );
  XOR2_X1 U1024 ( .A(KEYINPUT120), .B(G225), .Z(G308) );
  INV_X1 U1026 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(G325) );
  INV_X1 U1028 ( .A(G325), .ZN(G261) );
  INV_X1 U1029 ( .A(n929), .ZN(G319) );
  INV_X1 U1030 ( .A(G69), .ZN(G235) );
  INV_X1 U1031 ( .A(KEYINPUT55), .ZN(n977) );
  XNOR2_X1 U1032 ( .A(G2084), .B(G160), .ZN(n931) );
  NAND2_X1 U1033 ( .A1(n931), .A2(n930), .ZN(n939) );
  XOR2_X1 U1034 ( .A(G2072), .B(n932), .Z(n934) );
  XOR2_X1 U1035 ( .A(G164), .B(G2078), .Z(n933) );
  NOR2_X1 U1036 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1037 ( .A(n935), .B(KEYINPUT50), .ZN(n937) );
  NAND2_X1 U1038 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1039 ( .A1(n939), .A2(n938), .ZN(n951) );
  XNOR2_X1 U1040 ( .A(G2090), .B(G162), .ZN(n940) );
  XNOR2_X1 U1041 ( .A(n940), .B(KEYINPUT121), .ZN(n941) );
  NOR2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1043 ( .A(KEYINPUT51), .B(n943), .ZN(n944) );
  NOR2_X1 U1044 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n949) );
  NOR2_X1 U1046 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1048 ( .A(KEYINPUT52), .B(n952), .ZN(n953) );
  XOR2_X1 U1049 ( .A(KEYINPUT122), .B(n953), .Z(n954) );
  NAND2_X1 U1050 ( .A1(n977), .A2(n954), .ZN(n955) );
  NAND2_X1 U1051 ( .A1(n955), .A2(G29), .ZN(n1035) );
  XNOR2_X1 U1052 ( .A(KEYINPUT54), .B(G34), .ZN(n956) );
  XNOR2_X1 U1053 ( .A(n956), .B(KEYINPUT125), .ZN(n957) );
  XNOR2_X1 U1054 ( .A(G2084), .B(n957), .ZN(n975) );
  XNOR2_X1 U1055 ( .A(G2090), .B(G35), .ZN(n973) );
  XNOR2_X1 U1056 ( .A(G32), .B(n958), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(G2067), .B(G26), .ZN(n961) );
  XNOR2_X1 U1058 ( .A(G27), .B(n959), .ZN(n960) );
  NOR2_X1 U1059 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1060 ( .A1(n963), .A2(n962), .ZN(n965) );
  XNOR2_X1 U1061 ( .A(G33), .B(G2072), .ZN(n964) );
  NOR2_X1 U1062 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1063 ( .A(KEYINPUT124), .B(n966), .ZN(n967) );
  NAND2_X1 U1064 ( .A1(n967), .A2(G28), .ZN(n970) );
  XOR2_X1 U1065 ( .A(G25), .B(G1991), .Z(n968) );
  XNOR2_X1 U1066 ( .A(KEYINPUT123), .B(n968), .ZN(n969) );
  NOR2_X1 U1067 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1068 ( .A(KEYINPUT53), .B(n971), .ZN(n972) );
  NOR2_X1 U1069 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1071 ( .A(n977), .B(n976), .ZN(n979) );
  INV_X1 U1072 ( .A(G29), .ZN(n978) );
  NAND2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1074 ( .A1(G11), .A2(n980), .ZN(n1033) );
  XNOR2_X1 U1075 ( .A(G16), .B(KEYINPUT56), .ZN(n1005) );
  XNOR2_X1 U1076 ( .A(G1348), .B(n981), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n1003) );
  XNOR2_X1 U1079 ( .A(G1966), .B(G168), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1081 ( .A(n988), .B(KEYINPUT57), .ZN(n989) );
  XNOR2_X1 U1082 ( .A(KEYINPUT126), .B(n989), .ZN(n998) );
  XNOR2_X1 U1083 ( .A(n990), .B(G1956), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(G301), .B(G1961), .ZN(n992) );
  XNOR2_X1 U1085 ( .A(G303), .B(G1971), .ZN(n991) );
  NOR2_X1 U1086 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n1001) );
  XNOR2_X1 U1090 ( .A(G1341), .B(n999), .ZN(n1000) );
  NOR2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1031) );
  INV_X1 U1094 ( .A(G16), .ZN(n1029) );
  XOR2_X1 U1095 ( .A(G1986), .B(G24), .Z(n1009) );
  XNOR2_X1 U1096 ( .A(G1971), .B(G22), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(G23), .B(G1976), .ZN(n1006) );
  NOR2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(KEYINPUT127), .B(KEYINPUT58), .ZN(n1010) );
  XNOR2_X1 U1101 ( .A(n1011), .B(n1010), .ZN(n1015) );
  XNOR2_X1 U1102 ( .A(G1966), .B(G21), .ZN(n1013) );
  XNOR2_X1 U1103 ( .A(G5), .B(G1961), .ZN(n1012) );
  NOR2_X1 U1104 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1026) );
  XNOR2_X1 U1106 ( .A(G20), .B(n1016), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(G1341), .B(G19), .ZN(n1018) );
  XNOR2_X1 U1108 ( .A(G1981), .B(G6), .ZN(n1017) );
  NOR2_X1 U1109 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1110 ( .A1(n1020), .A2(n1019), .ZN(n1023) );
  XOR2_X1 U1111 ( .A(KEYINPUT59), .B(G1348), .Z(n1021) );
  XNOR2_X1 U1112 ( .A(G4), .B(n1021), .ZN(n1022) );
  NOR2_X1 U1113 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1114 ( .A(KEYINPUT60), .B(n1024), .Z(n1025) );
  NOR2_X1 U1115 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1116 ( .A(KEYINPUT61), .B(n1027), .ZN(n1028) );
  NAND2_X1 U1117 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1118 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1119 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1120 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XOR2_X1 U1121 ( .A(KEYINPUT62), .B(n1036), .Z(G311) );
  INV_X1 U1122 ( .A(G311), .ZN(G150) );
endmodule

