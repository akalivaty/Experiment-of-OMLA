//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 1 1 0 0 0 1 1 1 0 0 1 1 1 1 1 0 1 0 0 0 1 0 0 1 0 0 0 1 0 0 1 1 1 0 1 0 1 0 1 0 0 1 1 0 0 0 0 0 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999;
  XNOR2_X1  g000(.A(G143), .B(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(KEYINPUT0), .A2(G128), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  OR2_X1    g003(.A1(KEYINPUT0), .A2(G128), .ZN(new_n190));
  AND2_X1   g004(.A1(new_n190), .A2(new_n188), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n189), .B1(new_n191), .B2(new_n187), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G125), .ZN(new_n193));
  INV_X1    g007(.A(G128), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(KEYINPUT1), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G143), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G146), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n195), .A2(new_n197), .A3(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n198), .A2(KEYINPUT1), .A3(G146), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n200), .B(new_n201), .C1(G128), .C2(new_n187), .ZN(new_n202));
  INV_X1    g016(.A(G125), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G224), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(G953), .ZN(new_n206));
  OR2_X1    g020(.A1(new_n206), .A2(KEYINPUT85), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n193), .A2(new_n204), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n206), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT7), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n210), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n193), .A2(new_n204), .A3(new_n207), .A4(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G104), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT3), .B1(new_n215), .B2(G107), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT3), .ZN(new_n217));
  INV_X1    g031(.A(G107), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n218), .A3(G104), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n215), .A2(G107), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n216), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G101), .ZN(new_n222));
  INV_X1    g036(.A(G101), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n216), .A2(new_n219), .A3(new_n223), .A4(new_n220), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n222), .A2(KEYINPUT4), .A3(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT4), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n221), .A2(new_n226), .A3(G101), .ZN(new_n227));
  NOR2_X1   g041(.A1(KEYINPUT2), .A2(G113), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT68), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n230), .B1(KEYINPUT2), .B2(G113), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(KEYINPUT2), .A2(G113), .ZN(new_n233));
  AND2_X1   g047(.A1(KEYINPUT69), .A2(G119), .ZN(new_n234));
  NOR2_X1   g048(.A1(KEYINPUT69), .A2(G119), .ZN(new_n235));
  OAI21_X1  g049(.A(G116), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G119), .ZN(new_n237));
  OR2_X1    g051(.A1(new_n237), .A2(G116), .ZN(new_n238));
  AOI22_X1  g052(.A1(new_n232), .A2(new_n233), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  AND4_X1   g053(.A1(new_n232), .A2(new_n236), .A3(new_n233), .A4(new_n238), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n225), .B(new_n227), .C1(new_n239), .C2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n236), .A2(KEYINPUT5), .A3(new_n238), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT69), .B(G119), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT5), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n243), .A2(new_n244), .A3(G116), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n242), .A2(G113), .A3(new_n245), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n232), .A2(new_n236), .A3(new_n233), .A4(new_n238), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n218), .A2(G104), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n215), .A2(G107), .ZN(new_n249));
  OAI21_X1  g063(.A(G101), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n224), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n246), .A2(new_n247), .A3(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(G110), .B(G122), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n241), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n214), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  AOI211_X1 g070(.A(KEYINPUT84), .B(new_n251), .C1(new_n247), .C2(new_n246), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT84), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n246), .A2(new_n247), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n224), .A2(new_n250), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n252), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n253), .B(KEYINPUT8), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(G902), .B1(new_n256), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n193), .A2(new_n204), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n266), .B(new_n209), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n241), .A2(new_n252), .ZN(new_n269));
  XOR2_X1   g083(.A(new_n253), .B(KEYINPUT83), .Z(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n268), .B1(new_n271), .B2(new_n254), .ZN(new_n272));
  INV_X1    g086(.A(new_n270), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n273), .B1(new_n241), .B2(new_n252), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n274), .A2(KEYINPUT6), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n267), .B1(new_n272), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(G210), .B1(G237), .B2(G902), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n265), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT87), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n277), .B(KEYINPUT86), .ZN(new_n281));
  INV_X1    g095(.A(G902), .ZN(new_n282));
  INV_X1    g096(.A(new_n263), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n251), .B1(new_n246), .B2(new_n247), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n284), .B(new_n258), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n283), .B1(new_n285), .B2(new_n252), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n282), .B1(new_n286), .B2(new_n255), .ZN(new_n287));
  INV_X1    g101(.A(new_n267), .ZN(new_n288));
  INV_X1    g102(.A(new_n254), .ZN(new_n289));
  OAI21_X1  g103(.A(KEYINPUT6), .B1(new_n289), .B2(new_n274), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n271), .A2(new_n268), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n288), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n281), .B1(new_n287), .B2(new_n292), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n265), .A2(new_n276), .A3(KEYINPUT87), .A4(new_n277), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n280), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G953), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G952), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n297), .B1(G234), .B2(G237), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  XOR2_X1   g113(.A(KEYINPUT74), .B(G902), .Z(new_n300));
  NAND2_X1  g114(.A1(G234), .A2(G237), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(G953), .A3(new_n301), .ZN(new_n302));
  XOR2_X1   g116(.A(KEYINPUT21), .B(G898), .Z(new_n303));
  OAI21_X1  g117(.A(new_n299), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(G214), .B1(G237), .B2(G902), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n295), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G469), .ZN(new_n307));
  INV_X1    g121(.A(new_n300), .ZN(new_n308));
  OR2_X1    g122(.A1(new_n187), .A2(G128), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n260), .A2(new_n201), .A3(new_n309), .A4(new_n200), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n202), .A2(new_n224), .A3(new_n250), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AND2_X1   g126(.A1(KEYINPUT65), .A2(G137), .ZN(new_n313));
  NOR2_X1   g127(.A1(KEYINPUT65), .A2(G137), .ZN(new_n314));
  OAI211_X1 g128(.A(KEYINPUT11), .B(G134), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G137), .ZN(new_n316));
  OAI21_X1  g130(.A(KEYINPUT67), .B1(new_n316), .B2(G134), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT67), .ZN(new_n318));
  INV_X1    g132(.A(G134), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(new_n319), .A3(G137), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n316), .A2(G134), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT11), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n315), .A2(new_n321), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G131), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT66), .B(G131), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n315), .A2(new_n321), .A3(new_n324), .A4(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  AND3_X1   g143(.A1(new_n312), .A2(KEYINPUT12), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(KEYINPUT12), .B1(new_n312), .B2(new_n329), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n329), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n225), .A2(new_n192), .A3(new_n227), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n311), .A2(KEYINPUT10), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT10), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n336), .B1(new_n251), .B2(new_n202), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n333), .B(new_n334), .C1(new_n335), .C2(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(G110), .B(G140), .ZN(new_n339));
  INV_X1    g153(.A(G227), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n340), .A2(G953), .ZN(new_n341));
  XOR2_X1   g155(.A(new_n339), .B(new_n341), .Z(new_n342));
  NAND2_X1  g156(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n332), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n334), .B1(new_n335), .B2(new_n337), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n329), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n342), .B1(new_n346), .B2(new_n338), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n307), .B(new_n308), .C1(new_n344), .C2(new_n347), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n338), .A2(new_n342), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n346), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n338), .B1(new_n330), .B2(new_n331), .ZN(new_n351));
  INV_X1    g165(.A(new_n342), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(G902), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n348), .B(KEYINPUT81), .C1(new_n354), .C2(new_n307), .ZN(new_n355));
  XNOR2_X1  g169(.A(KEYINPUT9), .B(G234), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n356), .B(KEYINPUT79), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n282), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G221), .ZN(new_n359));
  XOR2_X1   g173(.A(new_n359), .B(KEYINPUT80), .Z(new_n360));
  INV_X1    g174(.A(KEYINPUT81), .ZN(new_n361));
  AOI22_X1  g175(.A1(new_n346), .A2(new_n349), .B1(new_n351), .B2(new_n352), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n361), .B(G469), .C1(new_n362), .C2(G902), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n355), .A2(new_n360), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT82), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n355), .A2(KEYINPUT82), .A3(new_n360), .A4(new_n363), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n306), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G110), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT23), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n370), .B1(new_n243), .B2(G128), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n237), .A2(G128), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n372), .B1(new_n243), .B2(G128), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n369), .B(new_n371), .C1(new_n373), .C2(new_n370), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT77), .ZN(new_n375));
  XOR2_X1   g189(.A(KEYINPUT24), .B(G110), .Z(new_n376));
  OAI21_X1  g190(.A(new_n375), .B1(new_n373), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(G128), .B1(new_n234), .B2(new_n235), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n378), .B1(new_n237), .B2(G128), .ZN(new_n379));
  INV_X1    g193(.A(new_n376), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(KEYINPUT77), .A3(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n374), .A2(new_n377), .A3(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT78), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G140), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G125), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n203), .A2(G140), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n387), .A3(KEYINPUT16), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT16), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(new_n385), .A3(G125), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT76), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n389), .A2(new_n385), .A3(KEYINPUT76), .A4(G125), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n388), .A2(new_n392), .A3(G146), .A4(new_n393), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n374), .A2(new_n377), .A3(new_n381), .A4(KEYINPUT78), .ZN(new_n395));
  XNOR2_X1  g209(.A(G125), .B(G140), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n196), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n384), .A2(new_n394), .A3(new_n395), .A4(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n371), .B1(new_n373), .B2(new_n370), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G110), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(KEYINPUT75), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n373), .A2(new_n376), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n388), .A2(new_n392), .A3(new_n393), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n196), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n394), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT75), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n399), .A2(new_n406), .A3(G110), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n401), .A2(new_n402), .A3(new_n405), .A4(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n398), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(KEYINPUT22), .B(G137), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n296), .A2(G221), .A3(G234), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n410), .B(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n398), .A2(new_n408), .A3(new_n412), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(new_n308), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT25), .ZN(new_n417));
  INV_X1    g231(.A(G217), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n418), .B1(new_n308), .B2(G234), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT25), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n414), .A2(new_n420), .A3(new_n308), .A4(new_n415), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n417), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  AND2_X1   g236(.A1(new_n414), .A2(new_n415), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n419), .A2(G902), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT72), .ZN(new_n427));
  AND4_X1   g241(.A1(new_n315), .A2(new_n321), .A3(new_n324), .A4(new_n327), .ZN(new_n428));
  INV_X1    g242(.A(G131), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n317), .A2(new_n320), .B1(new_n322), .B2(new_n323), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n429), .B1(new_n430), .B2(new_n315), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n192), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n240), .A2(new_n239), .ZN(new_n433));
  NOR3_X1   g247(.A1(new_n313), .A2(new_n314), .A3(G134), .ZN(new_n434));
  INV_X1    g248(.A(new_n322), .ZN(new_n435));
  OAI21_X1  g249(.A(G131), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n328), .A2(new_n436), .A3(new_n202), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n432), .A2(new_n433), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n432), .A2(KEYINPUT30), .A3(new_n437), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT70), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n432), .A2(KEYINPUT70), .A3(KEYINPUT30), .A4(new_n437), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n197), .A2(new_n199), .B1(new_n190), .B2(new_n188), .ZN(new_n445));
  AND3_X1   g259(.A1(new_n197), .A2(new_n199), .A3(new_n188), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n447), .B1(new_n326), .B2(new_n328), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n328), .A2(new_n436), .A3(new_n202), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n444), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n433), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n438), .B1(new_n443), .B2(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(G237), .A2(G953), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(G210), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(new_n223), .ZN(new_n456));
  XNOR2_X1  g270(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n457));
  XOR2_X1   g271(.A(new_n456), .B(new_n457), .Z(new_n458));
  OAI21_X1  g272(.A(new_n427), .B1(new_n453), .B2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n458), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n450), .A2(new_n451), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n461), .B1(new_n441), .B2(new_n442), .ZN(new_n462));
  OAI211_X1 g276(.A(KEYINPUT72), .B(new_n460), .C1(new_n462), .C2(new_n438), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT29), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT28), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n451), .B1(new_n448), .B2(new_n449), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n432), .A2(new_n433), .A3(new_n437), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n467), .A2(new_n465), .ZN(new_n469));
  OAI21_X1  g283(.A(KEYINPUT71), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n433), .B1(new_n432), .B2(new_n437), .ZN(new_n471));
  OAI21_X1  g285(.A(KEYINPUT28), .B1(new_n438), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT71), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n470), .A2(new_n458), .A3(new_n474), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n459), .A2(new_n463), .A3(new_n464), .A4(new_n475), .ZN(new_n476));
  OR2_X1    g290(.A1(new_n467), .A2(KEYINPUT73), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n467), .A2(KEYINPUT73), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(new_n466), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT28), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n467), .A2(new_n465), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n480), .A2(KEYINPUT29), .A3(new_n458), .A4(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n476), .A2(new_n308), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(G472), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT32), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n443), .A2(new_n452), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(new_n458), .A3(new_n467), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT31), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n473), .B1(new_n472), .B2(new_n481), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n468), .A2(KEYINPUT71), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n460), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT31), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n453), .A2(new_n492), .A3(new_n458), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n488), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(G472), .A2(G902), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n485), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n494), .A2(new_n485), .A3(new_n495), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n484), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n327), .ZN(new_n499));
  INV_X1    g313(.A(G237), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(new_n296), .A3(G214), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n501), .A2(new_n198), .ZN(new_n502));
  AOI21_X1  g316(.A(G143), .B1(new_n454), .B2(G214), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n499), .B(KEYINPUT17), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n404), .A2(new_n394), .A3(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT90), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n501), .B(new_n198), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n499), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n502), .A2(new_n503), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n327), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT17), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n509), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n404), .A2(KEYINPUT90), .A3(new_n394), .A4(new_n504), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n507), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(G113), .B(G122), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n516), .B(new_n215), .ZN(new_n517));
  NAND2_X1  g331(.A1(KEYINPUT18), .A2(G131), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n510), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT88), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n396), .B(new_n196), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT88), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n510), .A2(new_n522), .A3(new_n518), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n508), .A2(KEYINPUT18), .A3(G131), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n520), .A2(new_n521), .A3(new_n523), .A4(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n515), .A2(new_n517), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n509), .A2(new_n511), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT89), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n396), .A2(new_n528), .A3(KEYINPUT19), .ZN(new_n529));
  AOI21_X1  g343(.A(KEYINPUT19), .B1(new_n396), .B2(new_n528), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n196), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n527), .A2(new_n394), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n525), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n517), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n526), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(G475), .A2(G902), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n538), .A2(KEYINPUT91), .A3(KEYINPUT20), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT91), .ZN(new_n540));
  INV_X1    g354(.A(new_n537), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n541), .B1(new_n526), .B2(new_n535), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT20), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n540), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n536), .A2(new_n543), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n537), .B(KEYINPUT92), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n539), .B(new_n544), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n526), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n517), .B1(new_n515), .B2(new_n525), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n282), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  XOR2_X1   g364(.A(KEYINPUT93), .B(G475), .Z(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n198), .A2(G128), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n194), .A2(G143), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT94), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n555), .B1(new_n553), .B2(new_n554), .ZN(new_n557));
  NOR3_X1   g371(.A1(new_n556), .A2(new_n557), .A3(G134), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n194), .A2(G143), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n198), .A2(G128), .ZN(new_n560));
  OAI21_X1  g374(.A(KEYINPUT94), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n319), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(KEYINPUT95), .B1(new_n558), .B2(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(G116), .B(G122), .ZN(new_n565));
  AND2_X1   g379(.A1(new_n565), .A2(new_n218), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT14), .ZN(new_n567));
  INV_X1    g381(.A(G122), .ZN(new_n568));
  NOR3_X1   g382(.A1(new_n567), .A2(new_n568), .A3(G116), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n569), .B1(new_n567), .B2(new_n565), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n566), .B1(new_n570), .B2(G107), .ZN(new_n571));
  OAI21_X1  g385(.A(G134), .B1(new_n556), .B2(new_n557), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n561), .A2(new_n319), .A3(new_n562), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT95), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n564), .A2(new_n571), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n553), .A2(new_n554), .A3(KEYINPUT13), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n577), .B(G134), .C1(KEYINPUT13), .C2(new_n553), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n565), .A2(new_n218), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n573), .B(new_n578), .C1(new_n579), .C2(new_n566), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n357), .A2(G217), .A3(new_n296), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT96), .ZN(new_n584));
  INV_X1    g398(.A(new_n582), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n576), .A2(new_n580), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n576), .A2(KEYINPUT96), .A3(new_n580), .A4(new_n585), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n587), .A2(new_n308), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(G478), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n590), .A2(KEYINPUT15), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n591), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n587), .A2(new_n308), .A3(new_n588), .A4(new_n593), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n547), .A2(new_n552), .A3(new_n592), .A4(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n368), .A2(new_n426), .A3(new_n498), .A4(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(G101), .ZN(G3));
  NAND2_X1  g412(.A1(new_n422), .A2(new_n425), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n599), .B1(new_n366), .B2(new_n367), .ZN(new_n600));
  INV_X1    g414(.A(G472), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n601), .B1(new_n494), .B2(new_n308), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n602), .B1(new_n495), .B2(new_n494), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n547), .A2(new_n552), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT33), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n587), .A2(new_n606), .A3(new_n588), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n300), .A2(new_n590), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT98), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n586), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n576), .A2(KEYINPUT98), .A3(new_n580), .A4(new_n585), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n610), .A2(new_n583), .A3(KEYINPUT33), .A4(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n607), .A2(new_n608), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(KEYINPUT99), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n589), .A2(new_n590), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT99), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n607), .A2(new_n616), .A3(new_n608), .A4(new_n612), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n614), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n605), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT100), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n605), .A2(new_n618), .A3(KEYINPUT100), .ZN(new_n622));
  INV_X1    g436(.A(new_n305), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n277), .B1(new_n265), .B2(new_n276), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n623), .B1(new_n624), .B2(KEYINPUT97), .ZN(new_n625));
  INV_X1    g439(.A(new_n277), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n626), .B1(new_n287), .B2(new_n292), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT97), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(new_n628), .A3(new_n278), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n304), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n621), .A2(new_n622), .A3(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n604), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT34), .B(G104), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  NAND2_X1  g450(.A1(new_n592), .A2(new_n594), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n536), .A2(new_n543), .A3(new_n537), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n539), .A2(new_n544), .A3(new_n638), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n639), .A2(new_n552), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n632), .A2(new_n637), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n641), .A2(new_n603), .A3(new_n600), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT35), .B(G107), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  NOR2_X1   g458(.A1(new_n413), .A2(KEYINPUT36), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n409), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n424), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n422), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n368), .A2(new_n596), .A3(new_n603), .A4(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT37), .B(G110), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G12));
  OAI21_X1  g466(.A(new_n299), .B1(new_n302), .B2(G900), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n639), .A2(new_n637), .A3(new_n552), .A4(new_n653), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n648), .A2(new_n630), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n366), .A2(new_n367), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n655), .A2(new_n498), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(KEYINPUT101), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT101), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n655), .A2(new_n498), .A3(new_n656), .A4(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G128), .ZN(G30));
  XOR2_X1   g476(.A(new_n653), .B(KEYINPUT39), .Z(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n656), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT40), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n453), .A2(new_n460), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n282), .B1(new_n479), .B2(new_n458), .ZN(new_n668));
  OAI21_X1  g482(.A(G472), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n669), .B1(new_n497), .B2(new_n496), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(KEYINPUT102), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT102), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n672), .B(new_n669), .C1(new_n497), .C2(new_n496), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n648), .ZN(new_n675));
  INV_X1    g489(.A(new_n295), .ZN(new_n676));
  OR2_X1    g490(.A1(new_n676), .A2(KEYINPUT38), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(KEYINPUT38), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n605), .A2(new_n637), .A3(new_n305), .ZN(new_n680));
  NOR4_X1   g494(.A1(new_n666), .A2(new_n675), .A3(new_n679), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(new_n198), .ZN(G45));
  AND3_X1   g496(.A1(new_n605), .A2(new_n618), .A3(new_n653), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n648), .A2(new_n630), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n498), .A2(new_n656), .A3(new_n683), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G146), .ZN(G48));
  INV_X1    g500(.A(new_n344), .ZN(new_n687));
  INV_X1    g501(.A(new_n347), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n307), .B1(new_n689), .B2(new_n308), .ZN(new_n690));
  INV_X1    g504(.A(new_n348), .ZN(new_n691));
  INV_X1    g505(.A(new_n359), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n498), .A2(new_n426), .A3(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n621), .ZN(new_n696));
  INV_X1    g510(.A(new_n622), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n695), .A2(new_n698), .A3(new_n632), .ZN(new_n699));
  XNOR2_X1  g513(.A(KEYINPUT41), .B(G113), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G15));
  NAND2_X1  g515(.A1(new_n695), .A2(new_n641), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G116), .ZN(G18));
  NOR2_X1   g517(.A1(new_n595), .A2(new_n631), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n498), .A2(new_n684), .A3(new_n693), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G119), .ZN(G21));
  NAND4_X1  g520(.A1(new_n605), .A2(new_n637), .A3(new_n629), .A4(new_n625), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n690), .A2(new_n691), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n359), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT103), .ZN(new_n711));
  INV_X1    g525(.A(new_n495), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n488), .A2(new_n493), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n480), .A2(new_n481), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n460), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n712), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n716), .A2(new_n602), .A3(new_n599), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n710), .A2(new_n711), .A3(new_n304), .A4(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n630), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n719), .A2(new_n605), .A3(new_n637), .A4(new_n693), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n494), .A2(new_n308), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(G472), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n715), .A2(new_n493), .A3(new_n488), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n495), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n722), .A2(new_n426), .A3(new_n724), .A4(new_n304), .ZN(new_n725));
  OAI21_X1  g539(.A(KEYINPUT103), .B1(new_n720), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n718), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G122), .ZN(G24));
  NOR3_X1   g542(.A1(new_n648), .A2(new_n716), .A3(new_n602), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n709), .A2(new_n630), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n729), .A2(new_n683), .A3(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G125), .ZN(G27));
  NAND3_X1  g546(.A1(new_n605), .A2(new_n618), .A3(new_n653), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n280), .A2(new_n293), .A3(new_n294), .A4(new_n305), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g549(.A(G469), .B1(new_n362), .B2(G902), .ZN(new_n736));
  AOI21_X1  g550(.A(KEYINPUT104), .B1(new_n736), .B2(new_n348), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n736), .A2(KEYINPUT104), .A3(new_n348), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n692), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n735), .A2(new_n426), .A3(new_n498), .A4(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT42), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n494), .A2(new_n495), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(KEYINPUT32), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n494), .A2(new_n485), .A3(new_n495), .ZN(new_n746));
  AOI22_X1  g560(.A1(new_n745), .A2(new_n746), .B1(G472), .B2(new_n483), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n747), .A2(new_n599), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n748), .A2(KEYINPUT42), .A3(new_n735), .A4(new_n740), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n743), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G131), .ZN(G33));
  INV_X1    g565(.A(new_n739), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n359), .B1(new_n752), .B2(new_n737), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n747), .A2(new_n599), .A3(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT105), .ZN(new_n755));
  INV_X1    g569(.A(new_n654), .ZN(new_n756));
  INV_X1    g570(.A(new_n734), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n754), .A2(new_n755), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n498), .A2(new_n756), .A3(new_n426), .A4(new_n740), .ZN(new_n759));
  OAI21_X1  g573(.A(KEYINPUT105), .B1(new_n759), .B2(new_n734), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G134), .ZN(G36));
  NAND2_X1  g576(.A1(new_n350), .A2(new_n353), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(KEYINPUT106), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n763), .A2(new_n764), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(G469), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(G469), .A2(G902), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT46), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n348), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n770), .A2(new_n771), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n359), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT107), .ZN(new_n776));
  OR3_X1    g590(.A1(new_n775), .A2(new_n776), .A3(new_n663), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n776), .B1(new_n775), .B2(new_n663), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n547), .A2(new_n552), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n618), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT43), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n780), .B(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n603), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n782), .A2(new_n783), .A3(new_n649), .ZN(new_n784));
  AOI22_X1  g598(.A1(new_n777), .A2(new_n778), .B1(KEYINPUT44), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n784), .A2(KEYINPUT44), .ZN(new_n786));
  XOR2_X1   g600(.A(new_n734), .B(KEYINPUT108), .Z(new_n787));
  NOR2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G137), .ZN(G39));
  INV_X1    g604(.A(KEYINPUT47), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n775), .A2(new_n791), .ZN(new_n792));
  OAI211_X1 g606(.A(KEYINPUT47), .B(new_n359), .C1(new_n773), .C2(new_n774), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n794), .A2(new_n735), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n747), .A2(new_n599), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G140), .ZN(G42));
  AND2_X1   g613(.A1(new_n782), .A2(new_n298), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n709), .A2(new_n305), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT114), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n801), .A2(KEYINPUT114), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n803), .B1(new_n677), .B2(new_n678), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n800), .A2(new_n717), .A3(new_n802), .A4(new_n804), .ZN(new_n805));
  XOR2_X1   g619(.A(new_n805), .B(KEYINPUT50), .Z(new_n806));
  INV_X1    g620(.A(new_n787), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n800), .A2(new_n717), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  XOR2_X1   g623(.A(new_n708), .B(KEYINPUT109), .Z(new_n810));
  NOR2_X1   g624(.A1(new_n810), .A2(new_n360), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n807), .B(new_n809), .C1(new_n794), .C2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n674), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n709), .A2(new_n734), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n813), .A2(new_n426), .A3(new_n298), .A4(new_n814), .ZN(new_n815));
  OR3_X1    g629(.A1(new_n815), .A2(new_n605), .A3(new_n618), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n800), .A2(new_n814), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n729), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n806), .A2(new_n812), .A3(new_n816), .A4(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT51), .B1(new_n812), .B2(KEYINPUT115), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n815), .A2(new_n696), .A3(new_n697), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT116), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n823), .B1(new_n824), .B2(new_n297), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n297), .A2(new_n824), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n809), .A2(new_n730), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n825), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT117), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n825), .A2(KEYINPUT117), .A3(new_n827), .A4(new_n828), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n818), .A2(new_n748), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT48), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n831), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n820), .A2(new_n821), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n822), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n595), .B1(new_n779), .B2(new_n618), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n306), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n840), .A2(new_n600), .A3(new_n841), .A4(new_n603), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n597), .A2(new_n650), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n649), .A2(new_n653), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n640), .A2(new_n592), .A3(new_n594), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n498), .A2(new_n656), .A3(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n716), .A2(new_n602), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n847), .A2(new_n740), .A3(new_n605), .A4(new_n618), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n844), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n757), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n761), .A2(new_n843), .A3(new_n850), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n718), .A2(new_n726), .B1(new_n695), .B2(new_n641), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n705), .B1(new_n694), .B2(new_n633), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n852), .A2(new_n750), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n707), .A2(new_n753), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n674), .A2(new_n648), .A3(new_n653), .A4(new_n857), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n731), .A2(new_n685), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n661), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT52), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n661), .A2(new_n858), .A3(new_n859), .A4(KEYINPUT52), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n856), .A2(new_n864), .ZN(new_n865));
  XOR2_X1   g679(.A(KEYINPUT110), .B(KEYINPUT53), .Z(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  OR3_X1    g681(.A1(new_n865), .A2(KEYINPUT111), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT111), .B1(new_n865), .B2(new_n867), .ZN(new_n869));
  INV_X1    g683(.A(new_n865), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n868), .B(new_n869), .C1(KEYINPUT53), .C2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT54), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT113), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n862), .A2(new_n863), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n854), .A2(new_n702), .A3(new_n727), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n597), .A2(new_n650), .A3(new_n842), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n876), .B1(new_n757), .B2(new_n849), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n875), .A2(new_n877), .A3(new_n750), .A4(new_n761), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n867), .B1(new_n874), .B2(new_n878), .ZN(new_n879));
  AND4_X1   g693(.A1(KEYINPUT53), .A2(new_n761), .A3(new_n843), .A4(new_n850), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n855), .A2(KEYINPUT112), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT112), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n852), .A2(new_n750), .A3(new_n882), .A4(new_n854), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n864), .A2(new_n880), .A3(new_n881), .A4(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n879), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n873), .B1(new_n885), .B2(KEYINPUT54), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n885), .A2(KEYINPUT54), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(KEYINPUT113), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n838), .A2(new_n872), .A3(new_n886), .A4(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n833), .A2(new_n834), .ZN(new_n890));
  OAI22_X1  g704(.A1(new_n889), .A2(new_n890), .B1(G952), .B2(G953), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n810), .B(KEYINPUT49), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n426), .A2(new_n360), .A3(new_n305), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n892), .A2(new_n780), .A3(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n894), .A2(new_n813), .A3(new_n679), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n891), .A2(new_n895), .ZN(G75));
  AND4_X1   g710(.A1(new_n864), .A2(new_n880), .A3(new_n881), .A4(new_n883), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n866), .B1(new_n856), .B2(new_n864), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n899), .A2(new_n308), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT56), .B1(new_n900), .B2(new_n626), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n272), .A2(new_n275), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(new_n267), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT55), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n904), .B(KEYINPUT119), .ZN(new_n906));
  XOR2_X1   g720(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n907));
  AOI211_X1 g721(.A(new_n906), .B(new_n907), .C1(new_n900), .C2(new_n281), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n296), .A2(G952), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n905), .A2(new_n908), .A3(new_n909), .ZN(G51));
  XOR2_X1   g724(.A(new_n769), .B(KEYINPUT57), .Z(new_n911));
  AND2_X1   g725(.A1(new_n885), .A2(KEYINPUT54), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n911), .B1(new_n912), .B2(new_n887), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT120), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI211_X1 g729(.A(KEYINPUT120), .B(new_n911), .C1(new_n912), .C2(new_n887), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n915), .A2(new_n689), .A3(new_n916), .ZN(new_n917));
  OR3_X1    g731(.A1(new_n899), .A2(new_n308), .A3(new_n768), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n909), .B1(new_n917), .B2(new_n918), .ZN(G54));
  NAND3_X1  g733(.A1(new_n900), .A2(KEYINPUT58), .A3(G475), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(new_n536), .Z(new_n921));
  NOR2_X1   g735(.A1(new_n921), .A2(new_n909), .ZN(G60));
  NAND3_X1  g736(.A1(new_n872), .A2(new_n886), .A3(new_n888), .ZN(new_n923));
  NAND2_X1  g737(.A1(G478), .A2(G902), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT59), .Z(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  AOI22_X1  g740(.A1(new_n923), .A2(new_n926), .B1(new_n607), .B2(new_n612), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n912), .A2(new_n887), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n607), .A2(new_n612), .A3(new_n926), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n927), .A2(new_n909), .A3(new_n930), .ZN(G63));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n932));
  NAND2_X1  g746(.A1(G217), .A2(G902), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT121), .Z(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT60), .Z(new_n935));
  OAI211_X1 g749(.A(new_n646), .B(new_n935), .C1(new_n897), .C2(new_n898), .ZN(new_n936));
  INV_X1    g750(.A(new_n909), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n423), .B1(new_n885), .B2(new_n935), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n932), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT122), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT123), .ZN(new_n943));
  INV_X1    g757(.A(new_n935), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n879), .B2(new_n884), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n943), .B1(new_n945), .B2(new_n423), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n909), .B1(new_n945), .B2(new_n646), .ZN(new_n947));
  INV_X1    g761(.A(new_n423), .ZN(new_n948));
  OAI211_X1 g762(.A(KEYINPUT123), .B(new_n948), .C1(new_n899), .C2(new_n944), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n946), .A2(new_n947), .A3(new_n949), .A4(KEYINPUT61), .ZN(new_n950));
  OAI211_X1 g764(.A(KEYINPUT122), .B(new_n932), .C1(new_n938), .C2(new_n939), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n942), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT124), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n942), .A2(KEYINPUT124), .A3(new_n950), .A4(new_n951), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(G66));
  INV_X1    g770(.A(new_n303), .ZN(new_n957));
  OAI21_X1  g771(.A(G953), .B1(new_n957), .B2(new_n205), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n875), .A2(new_n843), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n958), .B1(new_n959), .B2(G953), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n902), .B1(G898), .B2(new_n296), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(G69));
  NAND2_X1  g776(.A1(new_n443), .A2(new_n450), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n529), .A2(new_n530), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n963), .B(new_n964), .Z(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n665), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n967), .A2(new_n748), .A3(new_n757), .A4(new_n840), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n789), .A2(new_n798), .A3(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT125), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(KEYINPUT62), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n661), .A2(new_n859), .A3(new_n971), .ZN(new_n972));
  OAI22_X1  g786(.A1(new_n681), .A2(new_n972), .B1(new_n970), .B2(KEYINPUT62), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n661), .A2(new_n859), .ZN(new_n974));
  OR4_X1    g788(.A1(new_n970), .A2(new_n681), .A3(KEYINPUT62), .A4(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n969), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n966), .B1(new_n976), .B2(new_n296), .ZN(new_n977));
  AOI22_X1  g791(.A1(new_n785), .A2(new_n788), .B1(new_n795), .B2(new_n797), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n707), .B1(new_n777), .B2(new_n778), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n974), .B1(new_n979), .B2(new_n748), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n761), .A2(new_n750), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n978), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n296), .ZN(new_n983));
  INV_X1    g797(.A(G900), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(G953), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT126), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n965), .B1(new_n983), .B2(new_n986), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n977), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(G953), .B1(new_n340), .B2(new_n984), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n988), .B(new_n989), .ZN(G72));
  NAND2_X1  g804(.A1(G472), .A2(G902), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT63), .Z(new_n992));
  NAND2_X1  g806(.A1(new_n875), .A2(new_n843), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n992), .B1(new_n976), .B2(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n909), .B1(new_n994), .B2(new_n667), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n992), .B1(new_n982), .B2(new_n993), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n996), .A2(new_n460), .A3(new_n453), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n459), .A2(new_n487), .A3(new_n463), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n871), .A2(new_n992), .A3(new_n998), .ZN(new_n999));
  AND3_X1   g813(.A1(new_n995), .A2(new_n997), .A3(new_n999), .ZN(G57));
endmodule


