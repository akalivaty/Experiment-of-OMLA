//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 0 1 0 0 1 0 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 1 0 1 1 1 1 0 1 0 1 0 1 1 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n810, new_n811, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XOR2_X1   g002(.A(new_n188), .B(KEYINPUT83), .Z(new_n189));
  INV_X1    g003(.A(G469), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(G110), .B(G140), .ZN(new_n193));
  INV_X1    g007(.A(G953), .ZN(new_n194));
  AND2_X1   g008(.A1(new_n194), .A2(G227), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n193), .B(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G143), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(KEYINPUT1), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  AND3_X1   g015(.A1(new_n201), .A2(KEYINPUT65), .A3(G146), .ZN(new_n202));
  AOI21_X1  g016(.A(KEYINPUT65), .B1(new_n201), .B2(G146), .ZN(new_n203));
  OAI211_X1 g017(.A(new_n198), .B(new_n200), .C1(new_n202), .C2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n205), .B1(new_n197), .B2(G143), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n201), .A2(KEYINPUT65), .A3(G146), .ZN(new_n207));
  AOI22_X1  g021(.A1(new_n206), .A2(new_n207), .B1(G143), .B2(new_n197), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT1), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n209), .B1(G143), .B2(new_n197), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(new_n199), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n204), .B1(new_n208), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G104), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT3), .B1(new_n213), .B2(G107), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n215));
  INV_X1    g029(.A(G107), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n216), .A3(G104), .ZN(new_n217));
  INV_X1    g031(.A(G101), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n213), .A2(G107), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n214), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n213), .A2(G107), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n216), .A2(G104), .ZN(new_n222));
  OAI21_X1  g036(.A(G101), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AND2_X1   g037(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n212), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT10), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n214), .A2(new_n217), .A3(new_n219), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G101), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(KEYINPUT4), .A3(new_n220), .ZN(new_n230));
  NAND2_X1  g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(KEYINPUT64), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT64), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(KEYINPUT0), .A3(G128), .ZN(new_n235));
  AND2_X1   g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n201), .A2(G146), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT0), .ZN(new_n238));
  AOI22_X1  g052(.A1(new_n198), .A2(new_n237), .B1(new_n238), .B2(new_n199), .ZN(new_n239));
  AOI22_X1  g053(.A1(new_n232), .A2(new_n208), .B1(new_n236), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT4), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n228), .A2(new_n241), .A3(G101), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n230), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n198), .A2(new_n237), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT66), .B(G128), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n244), .B1(new_n245), .B2(new_n210), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n226), .B1(new_n204), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(new_n224), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n227), .A2(new_n243), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT11), .ZN(new_n250));
  INV_X1    g064(.A(G134), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n250), .B1(new_n251), .B2(G137), .ZN(new_n252));
  INV_X1    g066(.A(G137), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(KEYINPUT11), .A3(G134), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n251), .A2(G137), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n252), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G131), .ZN(new_n257));
  INV_X1    g071(.A(G131), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n252), .A2(new_n254), .A3(new_n258), .A4(new_n255), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(KEYINPUT84), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n249), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n261), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n225), .A2(new_n226), .B1(new_n224), .B2(new_n247), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n263), .B1(new_n264), .B2(new_n243), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n196), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n220), .A2(new_n223), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(new_n246), .A3(new_n204), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n225), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n257), .A2(new_n259), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT12), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n264), .A2(new_n260), .A3(new_n243), .ZN(new_n273));
  INV_X1    g087(.A(new_n196), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n260), .B1(new_n225), .B2(new_n268), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT12), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n272), .A2(new_n273), .A3(new_n274), .A4(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(G902), .B1(new_n266), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n192), .B1(new_n279), .B2(new_n190), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n275), .A2(new_n276), .ZN(new_n281));
  AOI211_X1 g095(.A(KEYINPUT12), .B(new_n260), .C1(new_n225), .C2(new_n268), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n273), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n196), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n249), .A2(new_n261), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n264), .A2(new_n263), .A3(new_n243), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n287), .A3(new_n274), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n285), .A2(G469), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n189), .B1(new_n280), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(G214), .B1(G237), .B2(G902), .ZN(new_n291));
  OAI21_X1  g105(.A(G210), .B1(G237), .B2(G902), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n208), .A2(new_n232), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n238), .A2(new_n199), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n244), .A2(new_n294), .A3(new_n233), .A4(new_n235), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G125), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT1), .B1(new_n201), .B2(G146), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT66), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n299), .A2(G128), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n199), .A2(KEYINPUT66), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n298), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  AOI22_X1  g116(.A1(new_n208), .A2(new_n200), .B1(new_n302), .B2(new_n244), .ZN(new_n303));
  INV_X1    g117(.A(G125), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n297), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G224), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n307), .A2(G953), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n305), .B(new_n297), .C1(new_n307), .C2(G953), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT68), .ZN(new_n312));
  INV_X1    g126(.A(G116), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT69), .B1(new_n313), .B2(G119), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT69), .ZN(new_n315));
  INV_X1    g129(.A(G119), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(new_n316), .A3(G116), .ZN(new_n317));
  AND2_X1   g131(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT70), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n319), .B1(new_n316), .B2(G116), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n313), .A2(KEYINPUT70), .A3(G119), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n312), .B1(new_n318), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT2), .ZN(new_n324));
  INV_X1    g138(.A(G113), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT67), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT67), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n327), .A2(KEYINPUT2), .A3(G113), .ZN(new_n328));
  AOI22_X1  g142(.A1(new_n326), .A2(new_n328), .B1(new_n324), .B2(new_n325), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n323), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n314), .A2(new_n317), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(new_n320), .A3(new_n321), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(new_n312), .A3(new_n329), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n331), .A2(new_n334), .A3(new_n242), .A4(new_n230), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n318), .A2(new_n322), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n329), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n332), .A2(KEYINPUT5), .A3(new_n320), .A4(new_n321), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT5), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(new_n316), .A3(G116), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n340), .A2(G113), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n337), .A2(new_n224), .A3(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(G110), .B(G122), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n335), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n335), .A2(new_n343), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n344), .A2(KEYINPUT85), .ZN(new_n347));
  AOI22_X1  g161(.A1(new_n345), .A2(KEYINPUT6), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT6), .ZN(new_n349));
  INV_X1    g163(.A(new_n347), .ZN(new_n350));
  AOI211_X1 g164(.A(new_n349), .B(new_n350), .C1(new_n335), .C2(new_n343), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n311), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT86), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OAI211_X1 g168(.A(KEYINPUT86), .B(new_n311), .C1(new_n348), .C2(new_n351), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  XOR2_X1   g170(.A(new_n344), .B(KEYINPUT8), .Z(new_n357));
  AOI22_X1  g171(.A1(new_n336), .A2(new_n329), .B1(new_n338), .B2(new_n341), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n357), .B1(new_n358), .B2(new_n267), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT87), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n340), .A2(new_n360), .A3(G113), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n360), .B1(new_n340), .B2(G113), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI22_X1  g177(.A1(new_n338), .A2(new_n363), .B1(new_n336), .B2(new_n329), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n224), .B1(new_n364), .B2(KEYINPUT88), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(new_n338), .ZN(new_n366));
  AND3_X1   g180(.A1(new_n366), .A2(new_n337), .A3(KEYINPUT88), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n359), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n240), .A2(new_n304), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n204), .A2(new_n246), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n370), .A2(G125), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT7), .ZN(new_n372));
  OAI22_X1  g186(.A1(new_n369), .A2(new_n371), .B1(new_n372), .B2(new_n308), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT89), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT89), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n306), .B(new_n375), .C1(new_n372), .C2(new_n308), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n368), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n345), .B1(new_n310), .B2(new_n372), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n191), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n292), .B1(new_n356), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n292), .ZN(new_n382));
  AOI211_X1 g196(.A(new_n382), .B(new_n379), .C1(new_n354), .C2(new_n355), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n290), .B(new_n291), .C1(new_n381), .C2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT94), .ZN(new_n385));
  INV_X1    g199(.A(G140), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G125), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n304), .A2(G140), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT80), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n387), .A2(new_n388), .A3(KEYINPUT80), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n197), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n389), .A2(G146), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G237), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(new_n194), .A3(G214), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n201), .ZN(new_n398));
  NOR2_X1   g212(.A1(G237), .A2(G953), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(G143), .A3(G214), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(KEYINPUT18), .A2(G131), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n403), .ZN(new_n405));
  AOI21_X1  g219(.A(KEYINPUT90), .B1(new_n401), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT90), .ZN(new_n407));
  AOI211_X1 g221(.A(new_n407), .B(new_n403), .C1(new_n398), .C2(new_n400), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n395), .B(new_n404), .C1(new_n406), .C2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT91), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n393), .A2(new_n394), .B1(new_n402), .B2(new_n403), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT91), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n411), .B(new_n412), .C1(new_n406), .C2(new_n408), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(G113), .B(G122), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n415), .B(G104), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n417), .A2(KEYINPUT93), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n401), .A2(G131), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n258), .B1(new_n398), .B2(new_n400), .ZN(new_n420));
  NOR3_X1   g234(.A1(new_n419), .A2(KEYINPUT17), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n387), .A2(new_n388), .A3(KEYINPUT16), .ZN(new_n423));
  OR3_X1    g237(.A1(new_n304), .A2(KEYINPUT16), .A3(G140), .ZN(new_n424));
  AOI21_X1  g238(.A(G146), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT79), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n423), .A2(new_n424), .A3(G146), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  AND4_X1   g243(.A1(KEYINPUT79), .A2(new_n423), .A3(G146), .A4(new_n424), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n429), .A2(new_n431), .B1(KEYINPUT17), .B2(new_n420), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT92), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n422), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n423), .A2(G146), .A3(new_n424), .ZN(new_n435));
  NOR3_X1   g249(.A1(new_n435), .A2(new_n425), .A3(KEYINPUT79), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT17), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n401), .A2(G131), .ZN(new_n438));
  OAI22_X1  g252(.A1(new_n436), .A2(new_n430), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n439), .A2(KEYINPUT92), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n414), .B(new_n418), .C1(new_n434), .C2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n191), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n421), .B1(new_n439), .B2(KEYINPUT92), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n432), .A2(new_n433), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n418), .B1(new_n445), .B2(new_n414), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n385), .B1(new_n442), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n414), .B1(new_n434), .B2(new_n440), .ZN(new_n448));
  INV_X1    g262(.A(new_n418), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n450), .A2(KEYINPUT94), .A3(new_n191), .A4(new_n441), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n447), .A2(G475), .A3(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT19), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n391), .A2(new_n453), .A3(new_n392), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n389), .A2(KEYINPUT19), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n454), .A2(new_n197), .A3(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n428), .B1(new_n419), .B2(new_n420), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n416), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n458), .B1(new_n410), .B2(new_n413), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(G475), .A2(G902), .ZN(new_n461));
  AOI22_X1  g275(.A1(new_n443), .A2(new_n444), .B1(new_n413), .B2(new_n410), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n460), .B(new_n461), .C1(new_n462), .C2(new_n416), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(KEYINPUT20), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n459), .B1(new_n448), .B2(new_n417), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT20), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n465), .A2(new_n466), .A3(new_n461), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n194), .A2(G952), .ZN(new_n469));
  INV_X1    g283(.A(G234), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n469), .B1(new_n470), .B2(new_n396), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  AOI211_X1 g286(.A(new_n191), .B(new_n194), .C1(G234), .C2(G237), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT21), .B(G898), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n313), .A2(G122), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n216), .B1(new_n477), .B2(KEYINPUT14), .ZN(new_n478));
  XNOR2_X1  g292(.A(G116), .B(G122), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT14), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n482), .B(KEYINPUT96), .ZN(new_n483));
  OR3_X1    g297(.A1(new_n199), .A2(KEYINPUT95), .A3(G143), .ZN(new_n484));
  OAI21_X1  g298(.A(KEYINPUT95), .B1(new_n199), .B2(G143), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n245), .A2(G143), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(G134), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n486), .A2(new_n487), .A3(new_n251), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n479), .A2(new_n216), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n483), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n479), .B(new_n216), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT13), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n486), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n484), .A2(KEYINPUT13), .A3(new_n485), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n496), .A2(new_n497), .A3(new_n487), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n490), .B(new_n494), .C1(new_n498), .C2(new_n251), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n493), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(G217), .ZN(new_n501));
  NOR3_X1   g315(.A1(new_n187), .A2(new_n501), .A3(G953), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n493), .A2(new_n499), .A3(new_n502), .ZN(new_n505));
  AOI21_X1  g319(.A(G902), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(G478), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n507), .A2(KEYINPUT15), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n506), .B(new_n508), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n452), .A2(new_n468), .A3(new_n476), .A4(new_n509), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n384), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT32), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n333), .A2(new_n312), .A3(new_n329), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n329), .B1(new_n333), .B2(new_n312), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n240), .A2(new_n270), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT30), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n251), .A2(G137), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n253), .A2(G134), .ZN(new_n519));
  OAI21_X1  g333(.A(G131), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n259), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n370), .A2(new_n521), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n516), .A2(new_n517), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n517), .B1(new_n516), .B2(new_n522), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n515), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(KEYINPUT26), .B(G101), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT72), .ZN(new_n529));
  OR2_X1    g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n399), .A2(G210), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n528), .A2(new_n529), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n531), .B1(new_n530), .B2(new_n532), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n527), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n535), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(new_n526), .A3(new_n533), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n516), .B(new_n522), .C1(new_n514), .C2(new_n513), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n525), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT31), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n525), .A2(KEYINPUT31), .A3(new_n539), .A4(new_n540), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT28), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n259), .A2(new_n520), .ZN(new_n547));
  OAI22_X1  g361(.A1(new_n260), .A2(new_n296), .B1(new_n303), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n515), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n331), .A2(new_n334), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n550), .A2(KEYINPUT28), .A3(new_n516), .A4(new_n522), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n546), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n536), .A2(new_n538), .ZN(new_n553));
  AOI22_X1  g367(.A1(new_n543), .A2(new_n544), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(G472), .A2(G902), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n512), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n552), .A2(new_n553), .ZN(new_n558));
  INV_X1    g372(.A(new_n540), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n548), .A2(KEYINPUT30), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n516), .A2(new_n517), .A3(new_n522), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n559), .B1(new_n562), .B2(new_n515), .ZN(new_n563));
  AOI21_X1  g377(.A(KEYINPUT31), .B1(new_n563), .B2(new_n539), .ZN(new_n564));
  INV_X1    g378(.A(new_n544), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n558), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n566), .A2(KEYINPUT32), .A3(new_n555), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT73), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n549), .A2(new_n568), .A3(new_n540), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n548), .A2(new_n515), .A3(KEYINPUT73), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n569), .A2(KEYINPUT28), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n546), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT29), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n572), .A2(new_n573), .A3(new_n553), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n573), .B1(new_n552), .B2(new_n553), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n539), .B1(new_n525), .B2(new_n540), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n191), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(G472), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n557), .A2(new_n567), .A3(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(G217), .B1(new_n470), .B2(G902), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(KEYINPUT74), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT77), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n582), .B1(new_n316), .B2(G128), .ZN(new_n583));
  OAI21_X1  g397(.A(KEYINPUT23), .B1(new_n199), .B2(G119), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n199), .A2(KEYINPUT77), .A3(G119), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n199), .A2(KEYINPUT66), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n299), .A2(G128), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n587), .A2(new_n588), .A3(KEYINPUT23), .A4(G119), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(KEYINPUT78), .B1(new_n590), .B2(G110), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT78), .ZN(new_n592));
  INV_X1    g406(.A(G110), .ZN(new_n593));
  AOI211_X1 g407(.A(new_n592), .B(new_n593), .C1(new_n586), .C2(new_n589), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT75), .B1(new_n199), .B2(G119), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n596), .B1(new_n245), .B2(G119), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT75), .ZN(new_n598));
  AND4_X1   g412(.A1(new_n598), .A2(new_n587), .A3(new_n588), .A4(G119), .ZN(new_n599));
  OAI21_X1  g413(.A(KEYINPUT76), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  XOR2_X1   g414(.A(KEYINPUT24), .B(G110), .Z(new_n601));
  NAND3_X1  g415(.A1(new_n587), .A2(new_n588), .A3(G119), .ZN(new_n602));
  INV_X1    g416(.A(new_n596), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n245), .A2(new_n598), .A3(G119), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT76), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n600), .A2(new_n601), .A3(new_n607), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n595), .A2(new_n431), .A3(new_n429), .A4(new_n608), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n393), .A2(new_n428), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n601), .B1(new_n600), .B2(new_n607), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n590), .A2(G110), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(KEYINPUT22), .B(G137), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n194), .A2(G221), .A3(G234), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n609), .A2(new_n613), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n616), .B1(new_n609), .B2(new_n613), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(KEYINPUT25), .B1(new_n619), .B2(new_n191), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n609), .A2(new_n613), .ZN(new_n621));
  INV_X1    g435(.A(new_n616), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n609), .A2(new_n613), .A3(new_n616), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n623), .A2(KEYINPUT25), .A3(new_n191), .A4(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n581), .B1(new_n620), .B2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT81), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n623), .A2(new_n191), .A3(new_n624), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT25), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n625), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n633), .A2(KEYINPUT81), .A3(new_n581), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n581), .A2(G902), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(KEYINPUT82), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n619), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n629), .A2(new_n634), .A3(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n579), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n511), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G101), .ZN(G3));
  INV_X1    g455(.A(KEYINPUT97), .ZN(new_n642));
  INV_X1    g456(.A(G472), .ZN(new_n643));
  OAI211_X1 g457(.A(new_n566), .B(new_n191), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n645), .B1(new_n554), .B2(G902), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n266), .A2(new_n278), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n648), .A2(new_n190), .A3(new_n191), .ZN(new_n649));
  INV_X1    g463(.A(new_n192), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n649), .A2(new_n289), .A3(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n189), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n647), .A2(new_n653), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n629), .A2(new_n634), .A3(new_n637), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n654), .A2(new_n655), .A3(KEYINPUT98), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n291), .B(new_n476), .C1(new_n381), .C2(new_n383), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT33), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n658), .B1(new_n503), .B2(KEYINPUT99), .ZN(new_n659));
  AND3_X1   g473(.A1(new_n504), .A2(new_n505), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n659), .B1(new_n504), .B2(new_n505), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n507), .A2(G902), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g478(.A(KEYINPUT100), .B1(new_n506), .B2(G478), .ZN(new_n665));
  INV_X1    g479(.A(new_n505), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n502), .B1(new_n493), .B2(new_n499), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n191), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT100), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n668), .A2(new_n669), .A3(new_n507), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n665), .A2(new_n670), .ZN(new_n671));
  AOI22_X1  g485(.A1(new_n452), .A2(new_n468), .B1(new_n664), .B2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n657), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT98), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n290), .A2(new_n646), .A3(new_n644), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n675), .B1(new_n676), .B2(new_n638), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n656), .A2(new_n674), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT34), .B(G104), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G6));
  INV_X1    g494(.A(new_n509), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n681), .A2(new_n452), .A3(new_n468), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n657), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n656), .A2(new_n677), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT35), .B(G107), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT101), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n684), .B(new_n686), .ZN(G9));
  AOI21_X1  g501(.A(KEYINPUT81), .B1(new_n633), .B2(new_n581), .ZN(new_n688));
  INV_X1    g502(.A(new_n581), .ZN(new_n689));
  AOI211_X1 g503(.A(new_n628), .B(new_n689), .C1(new_n632), .C2(new_n625), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT102), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n621), .B(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n622), .A2(KEYINPUT36), .ZN(new_n694));
  AND2_X1   g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n693), .A2(new_n694), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n636), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n647), .B1(new_n691), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n511), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT37), .B(G110), .Z(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G12));
  INV_X1    g515(.A(new_n291), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n345), .A2(KEYINPUT6), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n346), .A2(new_n347), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n351), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g521(.A(KEYINPUT86), .B1(new_n707), .B2(new_n311), .ZN(new_n708));
  INV_X1    g522(.A(new_n355), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n380), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n382), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n356), .A2(new_n292), .A3(new_n380), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n702), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n557), .A2(new_n567), .A3(new_n578), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n629), .A2(new_n634), .A3(new_n697), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n713), .A2(new_n714), .A3(new_n715), .A4(new_n290), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n452), .A2(new_n468), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n473), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n471), .B1(new_n719), .B2(G900), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(KEYINPUT103), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n718), .A2(new_n681), .A3(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n716), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(new_n199), .ZN(G30));
  NOR2_X1   g539(.A1(new_n381), .A2(new_n383), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(KEYINPUT38), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n569), .A2(new_n553), .A3(new_n570), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n541), .A2(new_n729), .A3(G472), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n643), .A2(new_n191), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  AND3_X1   g546(.A1(new_n730), .A2(KEYINPUT104), .A3(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(KEYINPUT104), .B1(new_n730), .B2(new_n732), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n557), .A3(new_n567), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n717), .A2(new_n681), .ZN(new_n738));
  NOR4_X1   g552(.A1(new_n737), .A2(new_n738), .A3(new_n715), .A4(new_n702), .ZN(new_n739));
  XOR2_X1   g553(.A(new_n721), .B(KEYINPUT39), .Z(new_n740));
  AND2_X1   g554(.A1(new_n290), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(KEYINPUT40), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n728), .A2(new_n739), .A3(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(KEYINPUT105), .B(G143), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n743), .B(new_n744), .ZN(G45));
  INV_X1    g559(.A(new_n716), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n672), .A2(new_n722), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G146), .ZN(G48));
  AND4_X1   g564(.A1(new_n274), .A2(new_n272), .A3(new_n273), .A4(new_n277), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n274), .B1(new_n286), .B2(new_n287), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n191), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(G469), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n652), .A3(new_n649), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n579), .A2(new_n638), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n674), .ZN(new_n757));
  XNOR2_X1  g571(.A(KEYINPUT41), .B(G113), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(G15));
  AOI211_X1 g573(.A(new_n702), .B(new_n475), .C1(new_n711), .C2(new_n712), .ZN(new_n760));
  INV_X1    g574(.A(new_n682), .ZN(new_n761));
  INV_X1    g575(.A(new_n755), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n639), .A2(new_n760), .A3(new_n761), .A4(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G116), .ZN(G18));
  AOI211_X1 g578(.A(new_n702), .B(new_n755), .C1(new_n711), .C2(new_n712), .ZN(new_n765));
  INV_X1    g579(.A(new_n510), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n765), .A2(new_n714), .A3(new_n766), .A4(new_n715), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G119), .ZN(G21));
  NOR2_X1   g582(.A1(new_n554), .A2(G902), .ZN(new_n769));
  XOR2_X1   g583(.A(KEYINPUT106), .B(G472), .Z(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  AOI22_X1  g585(.A1(new_n543), .A2(new_n544), .B1(new_n572), .B2(new_n553), .ZN(new_n772));
  OAI22_X1  g586(.A1(new_n769), .A2(new_n771), .B1(new_n556), .B2(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n754), .A2(new_n652), .A3(new_n649), .A4(new_n476), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n638), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n291), .B1(new_n381), .B2(new_n383), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n776), .A2(new_n738), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G122), .ZN(G24));
  NAND2_X1  g593(.A1(new_n543), .A2(new_n544), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n572), .A2(new_n553), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n556), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n566), .A2(new_n191), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n782), .B1(new_n783), .B2(new_n770), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n715), .A2(new_n672), .A3(new_n722), .A4(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n713), .A2(new_n762), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(new_n304), .ZN(G27));
  NAND3_X1  g602(.A1(new_n691), .A2(new_n714), .A3(new_n637), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT108), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n274), .B1(new_n283), .B2(new_n273), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n262), .A2(new_n265), .A3(new_n196), .ZN(new_n793));
  OAI21_X1  g607(.A(KEYINPUT107), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT107), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n288), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n794), .A2(G469), .A3(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n189), .B1(new_n797), .B2(new_n280), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n798), .A2(new_n711), .A3(new_n291), .A4(new_n712), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n664), .A2(new_n671), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n717), .A2(KEYINPUT42), .A3(new_n800), .A4(new_n722), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n655), .A2(KEYINPUT108), .A3(new_n714), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n791), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n789), .A2(new_n799), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT42), .B1(new_n806), .B2(new_n748), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(new_n258), .ZN(G33));
  NOR3_X1   g623(.A1(new_n723), .A2(new_n789), .A3(new_n799), .ZN(new_n810));
  XOR2_X1   g624(.A(KEYINPUT109), .B(G134), .Z(new_n811));
  XNOR2_X1  g625(.A(new_n810), .B(new_n811), .ZN(G36));
  INV_X1    g626(.A(KEYINPUT43), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n718), .A2(new_n813), .A3(new_n800), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n800), .A2(new_n452), .A3(new_n468), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT43), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n814), .A2(new_n816), .A3(new_n647), .A4(new_n715), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT44), .ZN(new_n818));
  OR2_X1    g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT110), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n381), .A2(new_n383), .A3(new_n702), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n822), .B1(new_n817), .B2(new_n818), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n819), .A2(new_n820), .A3(new_n823), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n794), .A2(KEYINPUT45), .A3(new_n796), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n792), .A2(new_n793), .ZN(new_n826));
  OAI21_X1  g640(.A(G469), .B1(new_n826), .B2(KEYINPUT45), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n650), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT46), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n828), .A2(new_n829), .B1(new_n190), .B2(new_n279), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n189), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n832), .A2(new_n740), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n824), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n820), .B1(new_n819), .B2(new_n823), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(new_n253), .ZN(G39));
  NOR3_X1   g651(.A1(new_n822), .A2(new_n655), .A3(new_n714), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(new_n748), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n832), .A2(KEYINPUT47), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n832), .A2(KEYINPUT47), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n839), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(new_n386), .ZN(G42));
  INV_X1    g657(.A(KEYINPUT51), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n821), .A2(new_n762), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(KEYINPUT115), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n814), .A2(new_n816), .A3(new_n472), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n846), .A2(KEYINPUT116), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT116), .B1(new_n846), .B2(new_n847), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n715), .B(new_n784), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n847), .A2(new_n655), .A3(new_n784), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n727), .A2(new_n702), .A3(new_n762), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n853), .A2(KEYINPUT50), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n853), .A2(KEYINPUT50), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n846), .A2(new_n655), .A3(new_n472), .A4(new_n737), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n717), .A2(new_n800), .ZN(new_n857));
  OAI221_X1 g671(.A(new_n850), .B1(new_n854), .B2(new_n855), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n851), .A2(new_n822), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(KEYINPUT113), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n754), .A2(new_n649), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n861), .A2(new_n652), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n840), .A2(new_n841), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n862), .B1(new_n863), .B2(KEYINPUT114), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n863), .A2(KEYINPUT114), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n860), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n844), .B1(new_n858), .B2(new_n866), .ZN(new_n867));
  OAI221_X1 g681(.A(new_n469), .B1(new_n786), .B2(new_n851), .C1(new_n856), .C2(new_n673), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n791), .A2(new_n803), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n869), .B1(new_n848), .B2(new_n849), .ZN(new_n870));
  OR2_X1    g684(.A1(new_n870), .A2(KEYINPUT48), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(KEYINPUT48), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n868), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n863), .A2(new_n862), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n874), .B(KEYINPUT117), .Z(new_n875));
  OAI21_X1  g689(.A(KEYINPUT51), .B1(new_n875), .B2(new_n860), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n867), .B(new_n873), .C1(new_n876), .C2(new_n858), .ZN(new_n877));
  INV_X1    g691(.A(new_n810), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n726), .A2(new_n715), .A3(new_n291), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n653), .A2(new_n721), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n880), .A2(new_n714), .A3(new_n509), .A4(new_n718), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n672), .A2(new_n784), .A3(new_n722), .A4(new_n798), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n879), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n878), .B(new_n884), .C1(new_n805), .C2(new_n807), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n766), .A2(new_n714), .A3(new_n715), .ZN(new_n886));
  AOI22_X1  g700(.A1(new_n765), .A2(new_n886), .B1(new_n756), .B2(new_n683), .ZN(new_n887));
  AOI22_X1  g701(.A1(new_n674), .A2(new_n756), .B1(new_n511), .B2(new_n698), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n656), .B(new_n677), .C1(new_n674), .C2(new_n683), .ZN(new_n889));
  AOI22_X1  g703(.A1(new_n639), .A2(new_n511), .B1(new_n775), .B2(new_n777), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n887), .A2(new_n888), .A3(new_n889), .A4(new_n890), .ZN(new_n891));
  OAI22_X1  g705(.A1(new_n716), .A2(new_n723), .B1(new_n785), .B2(new_n786), .ZN(new_n892));
  AOI211_X1 g706(.A(new_n189), .B(new_n721), .C1(new_n797), .C2(new_n280), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n893), .A2(new_n691), .A3(new_n736), .A4(new_n697), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n509), .B1(new_n452), .B2(new_n468), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n895), .B(new_n291), .C1(new_n381), .C2(new_n383), .ZN(new_n896));
  OAI22_X1  g710(.A1(new_n716), .A2(new_n747), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n892), .A2(new_n897), .A3(KEYINPUT52), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n885), .A2(new_n891), .A3(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT53), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n892), .A2(KEYINPUT111), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT111), .ZN(new_n903));
  OAI221_X1 g717(.A(new_n903), .B1(new_n785), .B2(new_n786), .C1(new_n716), .C2(new_n723), .ZN(new_n904));
  INV_X1    g718(.A(new_n897), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n902), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT52), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT42), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n821), .A2(new_n655), .A3(new_n714), .A4(new_n798), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n908), .B1(new_n909), .B2(new_n747), .ZN(new_n910));
  AOI211_X1 g724(.A(new_n810), .B(new_n883), .C1(new_n910), .C2(new_n804), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n889), .A2(new_n890), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n757), .A2(new_n763), .A3(new_n767), .A4(new_n699), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(KEYINPUT52), .B1(new_n892), .B2(new_n897), .ZN(new_n915));
  INV_X1    g729(.A(new_n892), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT52), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n916), .A2(new_n905), .A3(new_n917), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n911), .A2(new_n914), .A3(new_n915), .A4(new_n918), .ZN(new_n919));
  AOI22_X1  g733(.A1(new_n901), .A2(new_n907), .B1(KEYINPUT53), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(KEYINPUT54), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT112), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n911), .A2(new_n914), .A3(KEYINPUT53), .A4(new_n918), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n906), .A2(KEYINPUT52), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n899), .A2(KEYINPUT112), .A3(KEYINPUT53), .A4(new_n907), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT54), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n919), .A2(new_n900), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n925), .A2(new_n926), .A3(new_n927), .A4(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n921), .A2(new_n929), .ZN(new_n930));
  OAI22_X1  g744(.A1(new_n877), .A2(new_n930), .B1(G952), .B2(G953), .ZN(new_n931));
  AOI211_X1 g745(.A(new_n702), .B(new_n189), .C1(new_n861), .C2(KEYINPUT49), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n932), .B1(KEYINPUT49), .B2(new_n861), .ZN(new_n933));
  NOR4_X1   g747(.A1(new_n933), .A2(new_n638), .A3(new_n736), .A4(new_n815), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n727), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n931), .A2(new_n935), .ZN(G75));
  NAND3_X1  g750(.A1(new_n925), .A2(new_n926), .A3(new_n928), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n937), .A2(G210), .A3(G902), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT56), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n707), .B(KEYINPUT118), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n311), .B(KEYINPUT119), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT55), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n941), .B(new_n943), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n938), .A2(new_n939), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n944), .B1(new_n938), .B2(new_n939), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n194), .A2(G952), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(G51));
  NAND2_X1  g762(.A1(new_n937), .A2(KEYINPUT54), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n929), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n192), .B(KEYINPUT57), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n648), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n825), .A2(new_n827), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n937), .A2(G902), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n947), .B1(new_n953), .B2(new_n955), .ZN(G54));
  NAND4_X1  g770(.A1(new_n937), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n957));
  INV_X1    g771(.A(new_n465), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n957), .A2(new_n958), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n959), .A2(new_n960), .A3(new_n947), .ZN(G60));
  INV_X1    g775(.A(new_n947), .ZN(new_n962));
  INV_X1    g776(.A(new_n950), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n662), .B(KEYINPUT120), .ZN(new_n964));
  XNOR2_X1  g778(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n965));
  NAND2_X1  g779(.A1(G478), .A2(G902), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n962), .B1(new_n963), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n964), .B1(new_n930), .B2(new_n967), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n969), .A2(new_n970), .ZN(G63));
  NAND2_X1  g785(.A1(G217), .A2(G902), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT122), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT60), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n937), .A2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n619), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n937), .B(new_n974), .C1(new_n695), .C2(new_n696), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n977), .A2(new_n962), .A3(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT61), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n977), .A2(KEYINPUT61), .A3(new_n978), .A4(new_n962), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(G66));
  OAI21_X1  g797(.A(G953), .B1(new_n474), .B2(new_n307), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n984), .B1(new_n914), .B2(G953), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n941), .B1(G898), .B2(new_n194), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n985), .B(new_n986), .ZN(G69));
  AOI21_X1  g801(.A(new_n194), .B1(G227), .B2(G900), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT124), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n824), .A2(new_n833), .ZN(new_n991));
  INV_X1    g805(.A(new_n835), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n842), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n743), .A2(new_n902), .A3(new_n904), .A4(new_n749), .ZN(new_n994));
  OR2_X1    g808(.A1(new_n994), .A2(KEYINPUT62), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n639), .A2(new_n741), .A3(new_n821), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n996), .B1(new_n673), .B2(new_n682), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n997), .B1(new_n994), .B2(KEYINPUT62), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n993), .A2(new_n995), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(new_n194), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n454), .A2(new_n455), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1001), .B(KEYINPUT123), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n562), .B(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1000), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1004), .B1(G900), .B2(G953), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(new_n842), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1008), .B1(new_n834), .B2(new_n835), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n808), .A2(new_n810), .ZN(new_n1010));
  AND2_X1   g824(.A1(new_n902), .A2(new_n904), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n833), .A2(new_n777), .A3(new_n869), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n1010), .A2(new_n749), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n1009), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1007), .B1(new_n1014), .B2(new_n194), .ZN(new_n1015));
  INV_X1    g829(.A(new_n1015), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n990), .B1(new_n1005), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1003), .B1(new_n999), .B2(new_n194), .ZN(new_n1018));
  NOR3_X1   g832(.A1(new_n1018), .A2(new_n1015), .A3(KEYINPUT124), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n989), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n1005), .A2(new_n1016), .A3(new_n990), .ZN(new_n1021));
  OAI21_X1  g835(.A(KEYINPUT124), .B1(new_n1018), .B2(new_n1015), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1021), .A2(new_n988), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1020), .A2(new_n1023), .ZN(G72));
  XNOR2_X1  g838(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n732), .B(new_n1025), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1026), .B1(new_n999), .B2(new_n891), .ZN(new_n1027));
  XNOR2_X1  g841(.A(new_n563), .B(KEYINPUT126), .ZN(new_n1028));
  INV_X1    g842(.A(new_n1028), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n1027), .A2(new_n539), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g844(.A(KEYINPUT127), .ZN(new_n1031));
  AND2_X1   g845(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g846(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1033));
  NOR3_X1   g847(.A1(new_n1009), .A2(new_n1013), .A3(new_n891), .ZN(new_n1034));
  INV_X1    g848(.A(new_n1026), .ZN(new_n1035));
  OAI211_X1 g849(.A(new_n553), .B(new_n1028), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  INV_X1    g850(.A(new_n576), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n1035), .B1(new_n1037), .B2(new_n541), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n920), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g853(.A1(new_n1036), .A2(new_n1039), .A3(new_n962), .ZN(new_n1040));
  NOR3_X1   g854(.A1(new_n1032), .A2(new_n1033), .A3(new_n1040), .ZN(G57));
endmodule


