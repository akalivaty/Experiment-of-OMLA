//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 0 1 0 1 1 1 1 0 1 1 0 0 0 0 1 0 0 0 1 0 1 1 1 0 0 0 0 0 1 1 0 0 0 0 1 0 1 0 1 1 1 0 1 0 0 0 1 1 0 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:59 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n565, new_n567, new_n568, new_n570, new_n571, new_n572, new_n573,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT66), .Z(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(new_n454), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n467), .A3(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n464), .A2(KEYINPUT67), .A3(G2104), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n472), .A2(new_n467), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n475), .B1(new_n466), .B2(KEYINPUT3), .ZN(new_n476));
  NAND4_X1  g051(.A1(new_n473), .A2(G137), .A3(new_n474), .A4(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n478));
  OAI21_X1  g053(.A(KEYINPUT68), .B1(new_n466), .B2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n480), .A2(new_n474), .A3(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n478), .B1(new_n482), .B2(G101), .ZN(new_n483));
  INV_X1    g058(.A(G101), .ZN(new_n484));
  AOI211_X1 g059(.A(KEYINPUT69), .B(new_n484), .C1(new_n479), .C2(new_n481), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n471), .B(new_n477), .C1(new_n483), .C2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G160));
  NAND4_X1  g062(.A1(new_n476), .A2(new_n472), .A3(G2105), .A4(new_n467), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  AND2_X1   g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  OR2_X1    g065(.A1(G100), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G112), .C2(new_n474), .ZN(new_n492));
  XOR2_X1   g067(.A(new_n492), .B(KEYINPUT70), .Z(new_n493));
  AND3_X1   g068(.A1(new_n473), .A2(new_n474), .A3(new_n476), .ZN(new_n494));
  AOI211_X1 g069(.A(new_n490), .B(new_n493), .C1(G136), .C2(new_n494), .ZN(G162));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n476), .A2(new_n472), .A3(new_n497), .A4(new_n467), .ZN(new_n498));
  AND2_X1   g073(.A1(new_n465), .A2(new_n467), .ZN(new_n499));
  NOR3_X1   g074(.A1(new_n496), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n498), .A2(KEYINPUT4), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G126), .ZN(new_n502));
  OR2_X1    g077(.A1(KEYINPUT71), .A2(G114), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT71), .A2(G114), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n474), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g080(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n506));
  OAI22_X1  g081(.A1(new_n488), .A2(new_n502), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n501), .A2(new_n507), .ZN(G164));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT72), .B1(new_n509), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n511), .A2(new_n512), .A3(KEYINPUT5), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n512), .A2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n514), .A2(G62), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT6), .B(G651), .ZN(new_n521));
  AND2_X1   g096(.A1(KEYINPUT73), .A2(G88), .ZN(new_n522));
  NOR2_X1   g097(.A1(KEYINPUT73), .A2(G88), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n514), .A2(new_n516), .A3(new_n521), .A4(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n521), .A2(G50), .A3(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n520), .A2(new_n528), .A3(KEYINPUT74), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT74), .ZN(new_n530));
  INV_X1    g105(.A(G651), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n531), .B1(new_n517), .B2(new_n518), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n530), .B1(new_n532), .B2(new_n527), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n529), .A2(new_n533), .ZN(G166));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT75), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n515), .B1(new_n510), .B2(new_n513), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n538), .A2(new_n521), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G89), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(KEYINPUT76), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT76), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n537), .A2(new_n543), .A3(new_n540), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n521), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  AND2_X1   g121(.A1(G63), .A2(G651), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n546), .A2(G51), .B1(new_n538), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n542), .A2(new_n544), .A3(new_n548), .ZN(G286));
  INV_X1    g124(.A(G286), .ZN(G168));
  AOI22_X1  g125(.A1(new_n538), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n551), .A2(new_n531), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n538), .A2(new_n521), .ZN(new_n553));
  INV_X1    g128(.A(G90), .ZN(new_n554));
  INV_X1    g129(.A(G52), .ZN(new_n555));
  OAI22_X1  g130(.A1(new_n553), .A2(new_n554), .B1(new_n555), .B2(new_n545), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n552), .A2(new_n556), .ZN(G171));
  AOI22_X1  g132(.A1(new_n538), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n558), .A2(new_n531), .ZN(new_n559));
  INV_X1    g134(.A(G81), .ZN(new_n560));
  INV_X1    g135(.A(G43), .ZN(new_n561));
  OAI22_X1  g136(.A1(new_n553), .A2(new_n560), .B1(new_n561), .B2(new_n545), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT77), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(G188));
  NAND3_X1  g144(.A1(new_n521), .A2(G53), .A3(G543), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT9), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n539), .A2(G91), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n538), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n573));
  OAI211_X1 g148(.A(new_n571), .B(new_n572), .C1(new_n531), .C2(new_n573), .ZN(G299));
  INV_X1    g149(.A(G171), .ZN(G301));
  INV_X1    g150(.A(G166), .ZN(G303));
  OAI21_X1  g151(.A(G651), .B1(new_n538), .B2(G74), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n538), .A2(G87), .A3(new_n521), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n521), .A2(G49), .A3(G543), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G288));
  NAND3_X1  g155(.A1(new_n521), .A2(G48), .A3(G543), .ZN(new_n581));
  INV_X1    g156(.A(G86), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n553), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n538), .A2(G61), .ZN(new_n585));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(G651), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n584), .A2(new_n588), .ZN(G305));
  INV_X1    g164(.A(G85), .ZN(new_n590));
  INV_X1    g165(.A(G47), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n553), .A2(new_n590), .B1(new_n591), .B2(new_n545), .ZN(new_n592));
  AND2_X1   g167(.A1(new_n592), .A2(KEYINPUT78), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n592), .A2(KEYINPUT78), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n538), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n593), .A2(new_n594), .B1(new_n531), .B2(new_n595), .ZN(G290));
  INV_X1    g171(.A(G92), .ZN(new_n597));
  XNOR2_X1  g172(.A(KEYINPUT79), .B(KEYINPUT10), .ZN(new_n598));
  OR3_X1    g173(.A1(new_n553), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n538), .A2(G66), .ZN(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G651), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n546), .A2(G54), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n598), .B1(new_n553), .B2(new_n597), .ZN(new_n605));
  NAND4_X1  g180(.A1(new_n599), .A2(new_n603), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(new_n607), .B2(G171), .ZN(G284));
  OAI21_X1  g184(.A(new_n608), .B1(new_n607), .B2(G171), .ZN(G321));
  NAND2_X1  g185(.A1(G299), .A2(new_n607), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(G168), .B2(new_n607), .ZN(G297));
  OAI21_X1  g187(.A(new_n611), .B1(G168), .B2(new_n607), .ZN(G280));
  INV_X1    g188(.A(new_n606), .ZN(new_n614));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G860), .ZN(G148));
  OAI21_X1  g191(.A(KEYINPUT80), .B1(new_n563), .B2(G868), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n606), .A2(G559), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n618), .A2(new_n607), .ZN(new_n619));
  MUX2_X1   g194(.A(new_n617), .B(KEYINPUT80), .S(new_n619), .Z(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT81), .Z(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g197(.A1(new_n499), .A2(new_n482), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT12), .ZN(new_n624));
  XOR2_X1   g199(.A(KEYINPUT82), .B(G2100), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n624), .B(new_n626), .ZN(new_n627));
  OR2_X1    g202(.A1(G99), .A2(G2105), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n628), .B(G2104), .C1(G111), .C2(new_n474), .ZN(new_n629));
  INV_X1    g204(.A(G123), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n488), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n631), .B1(new_n494), .B2(G135), .ZN(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n633), .A2(G2096), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(G2096), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n627), .A2(new_n634), .A3(new_n635), .ZN(G156));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT85), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2430), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(KEYINPUT14), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G1341), .B(G1348), .Z(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n643), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2451), .B(G2454), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT84), .ZN(new_n649));
  XOR2_X1   g224(.A(G2443), .B(G2446), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n647), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(G14), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT86), .ZN(G401));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT87), .ZN(new_n658));
  NOR2_X1   g233(.A1(G2072), .A2(G2078), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n442), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n656), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(KEYINPUT17), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n661), .B1(new_n658), .B2(new_n662), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n656), .B(new_n657), .C1(new_n442), .C2(new_n659), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT18), .Z(new_n665));
  NAND3_X1  g240(.A1(new_n662), .A2(new_n658), .A3(new_n656), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n663), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2096), .B(G2100), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(G227));
  XNOR2_X1  g244(.A(G1971), .B(G1976), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G1956), .B(G2474), .Z(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  AND2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT20), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n673), .A2(new_n674), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n672), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT89), .ZN(new_n680));
  OR3_X1    g255(.A1(new_n672), .A2(new_n675), .A3(new_n678), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n677), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G1991), .B(G1996), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1981), .B(G1986), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(G229));
  NOR2_X1   g264(.A1(G29), .A2(G35), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(G162), .B2(G29), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT29), .Z(new_n692));
  INV_X1    g267(.A(G2090), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n692), .A2(new_n693), .ZN(new_n695));
  INV_X1    g270(.A(G16), .ZN(new_n696));
  NOR2_X1   g271(.A1(G171), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(G5), .B2(new_n696), .ZN(new_n698));
  INV_X1    g273(.A(G1961), .ZN(new_n699));
  INV_X1    g274(.A(G29), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G27), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(G164), .B2(new_n700), .ZN(new_n702));
  AOI22_X1  g277(.A1(new_n698), .A2(new_n699), .B1(new_n702), .B2(G2078), .ZN(new_n703));
  INV_X1    g278(.A(G2084), .ZN(new_n704));
  INV_X1    g279(.A(G34), .ZN(new_n705));
  AOI21_X1  g280(.A(G29), .B1(new_n705), .B2(KEYINPUT24), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(KEYINPUT24), .B2(new_n705), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(new_n486), .B2(new_n700), .ZN(new_n708));
  OAI221_X1 g283(.A(new_n703), .B1(G2078), .B2(new_n702), .C1(new_n704), .C2(new_n708), .ZN(new_n709));
  OR3_X1    g284(.A1(new_n694), .A2(new_n695), .A3(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT97), .B(KEYINPUT28), .Z(new_n711));
  NAND2_X1  g286(.A1(new_n700), .A2(G26), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n489), .A2(G128), .ZN(new_n714));
  OAI21_X1  g289(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G116), .B2(new_n474), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT96), .ZN(new_n718));
  AOI211_X1 g293(.A(new_n714), .B(new_n718), .C1(G140), .C2(new_n494), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n713), .B1(new_n719), .B2(new_n700), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(G2067), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n696), .A2(G20), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT23), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n571), .A2(new_n572), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n573), .A2(new_n531), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n723), .B1(new_n726), .B2(new_n696), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G1956), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n696), .A2(G19), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(new_n563), .B2(new_n696), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G1341), .ZN(new_n731));
  NOR3_X1   g306(.A1(new_n721), .A2(new_n728), .A3(new_n731), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT25), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n499), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n735), .A2(new_n474), .ZN(new_n736));
  AOI211_X1 g311(.A(new_n734), .B(new_n736), .C1(G139), .C2(new_n494), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G29), .ZN(new_n738));
  NOR2_X1   g313(.A1(G29), .A2(G33), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT98), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n738), .A2(G2072), .A3(new_n740), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT31), .B(G11), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT30), .B(G28), .Z(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(new_n743), .B2(G29), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n632), .B2(G29), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n708), .A2(new_n704), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n698), .B2(new_n699), .ZN(new_n748));
  AOI21_X1  g323(.A(G2072), .B1(new_n738), .B2(new_n740), .ZN(new_n749));
  NOR3_X1   g324(.A1(new_n746), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n696), .A2(G4), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n614), .B2(new_n696), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(G1348), .Z(new_n753));
  NAND3_X1  g328(.A1(new_n732), .A2(new_n750), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n494), .A2(G141), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT99), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n482), .A2(G105), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT100), .B(KEYINPUT26), .ZN(new_n758));
  NAND3_X1  g333(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  AOI211_X1 g335(.A(new_n757), .B(new_n760), .C1(G129), .C2(new_n489), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n756), .A2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n763), .A2(G29), .ZN(new_n764));
  NOR2_X1   g339(.A1(G29), .A2(G32), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(KEYINPUT101), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(KEYINPUT101), .B2(new_n764), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT27), .B(G1996), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n696), .A2(G21), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G168), .B2(new_n696), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT103), .B(G1966), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT102), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n771), .B(new_n773), .ZN(new_n774));
  NOR4_X1   g349(.A1(new_n710), .A2(new_n754), .A3(new_n769), .A4(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n696), .A2(G23), .ZN(new_n777));
  NAND2_X1  g352(.A1(G288), .A2(KEYINPUT93), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT93), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n577), .A2(new_n578), .A3(new_n779), .A4(new_n579), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n777), .B1(new_n782), .B2(new_n696), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT94), .Z(new_n784));
  XOR2_X1   g359(.A(KEYINPUT33), .B(G1976), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT95), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n696), .A2(G6), .ZN(new_n789));
  INV_X1    g364(.A(G305), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(new_n696), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT91), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT32), .B(G1981), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT92), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n792), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n784), .A2(new_n787), .ZN(new_n796));
  NOR2_X1   g371(.A1(G16), .A2(G22), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G166), .B2(G16), .ZN(new_n798));
  INV_X1    g373(.A(G1971), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n788), .A2(new_n795), .A3(new_n796), .A4(new_n800), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(KEYINPUT34), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(KEYINPUT34), .ZN(new_n803));
  OR2_X1    g378(.A1(G16), .A2(G24), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G290), .B2(new_n696), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(G1986), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n806), .A2(G1986), .ZN(new_n808));
  NOR2_X1   g383(.A1(G25), .A2(G29), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n494), .A2(G131), .ZN(new_n810));
  INV_X1    g385(.A(G119), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n474), .A2(G107), .ZN(new_n812));
  OAI21_X1  g387(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n813));
  OAI22_X1  g388(.A1(new_n488), .A2(new_n811), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n809), .B1(new_n815), .B2(G29), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT35), .B(G1991), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT90), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n816), .B(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n808), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n802), .A2(new_n803), .A3(new_n807), .A4(new_n820), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(KEYINPUT36), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(KEYINPUT36), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n776), .B1(new_n822), .B2(new_n823), .ZN(G311));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n823), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(new_n775), .ZN(G150));
  AOI22_X1  g401(.A1(new_n538), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n827), .A2(new_n531), .ZN(new_n828));
  INV_X1    g403(.A(G93), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT105), .B(G55), .Z(new_n830));
  OAI22_X1  g405(.A1(new_n553), .A2(new_n829), .B1(new_n545), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(G860), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(KEYINPUT107), .B(KEYINPUT37), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n606), .A2(new_n615), .ZN(new_n837));
  XOR2_X1   g412(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n832), .A2(new_n563), .ZN(new_n840));
  OAI22_X1  g415(.A1(new_n828), .A2(new_n831), .B1(new_n559), .B2(new_n562), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n839), .B(new_n842), .Z(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(KEYINPUT39), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT106), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n833), .B1(new_n844), .B2(KEYINPUT39), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n836), .B1(new_n846), .B2(new_n847), .ZN(G145));
  XNOR2_X1  g423(.A(new_n762), .B(new_n737), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n489), .A2(G130), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n474), .A2(G118), .ZN(new_n851));
  OAI21_X1  g426(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(G142), .B2(new_n494), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n624), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n849), .B(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n719), .B(G164), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n815), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n856), .A2(new_n858), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(G160), .B(new_n632), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(G162), .Z(new_n863));
  AOI21_X1  g438(.A(G37), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(new_n863), .B2(new_n861), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g441(.A(new_n607), .B1(new_n828), .B2(new_n831), .ZN(new_n867));
  XNOR2_X1  g442(.A(G290), .B(G305), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(G303), .A2(KEYINPUT111), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(G303), .A2(KEYINPUT111), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n781), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n872), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n874), .A2(new_n870), .A3(new_n782), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n869), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n782), .B1(new_n874), .B2(new_n870), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n871), .A2(new_n781), .A3(new_n872), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n877), .A2(new_n878), .A3(new_n868), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT42), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n842), .B(new_n618), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n614), .A2(G299), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(KEYINPUT108), .B1(new_n614), .B2(G299), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT108), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n726), .A2(new_n886), .A3(new_n606), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n884), .B1(new_n888), .B2(KEYINPUT109), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT109), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n885), .A2(new_n890), .A3(new_n887), .ZN(new_n891));
  AOI21_X1  g466(.A(KEYINPUT41), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n726), .A2(new_n886), .A3(new_n606), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n886), .B1(new_n726), .B2(new_n606), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n895), .A2(KEYINPUT110), .A3(KEYINPUT41), .A4(new_n883), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n885), .A2(KEYINPUT41), .A3(new_n883), .A4(new_n887), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT110), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n882), .B1(new_n892), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n895), .A2(new_n883), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n901), .B1(new_n903), .B2(new_n882), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n881), .B(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n867), .B1(new_n905), .B2(new_n607), .ZN(G295));
  OAI21_X1  g481(.A(new_n867), .B1(new_n905), .B2(new_n607), .ZN(G331));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n908));
  AND2_X1   g483(.A1(new_n876), .A2(new_n879), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n840), .A2(G301), .A3(new_n841), .ZN(new_n910));
  AOI21_X1  g485(.A(G301), .B1(new_n840), .B2(new_n841), .ZN(new_n911));
  OAI21_X1  g486(.A(G286), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n842), .A2(G171), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n840), .A2(G301), .A3(new_n841), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n913), .A2(G168), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n897), .B(KEYINPUT110), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT109), .B1(new_n893), .B2(new_n894), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n918), .A2(new_n891), .A3(new_n883), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT41), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n916), .B1(new_n917), .B2(new_n921), .ZN(new_n922));
  NOR3_X1   g497(.A1(new_n910), .A2(new_n911), .A3(G286), .ZN(new_n923));
  AOI21_X1  g498(.A(G168), .B1(new_n913), .B2(new_n914), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n902), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n909), .B1(new_n922), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(G37), .ZN(new_n928));
  INV_X1    g503(.A(new_n916), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n929), .B1(new_n892), .B2(new_n900), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n930), .A2(new_n880), .A3(new_n925), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n927), .A2(new_n928), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n919), .A2(KEYINPUT41), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n885), .A2(new_n920), .A3(new_n883), .A4(new_n887), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n912), .A2(new_n915), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n925), .A2(KEYINPUT112), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT112), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n916), .A2(new_n940), .A3(new_n902), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n938), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n909), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n943), .A2(new_n931), .A3(KEYINPUT43), .A4(new_n928), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n908), .B1(new_n934), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n932), .A2(KEYINPUT43), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n943), .A2(new_n931), .A3(new_n933), .A4(new_n928), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT44), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT113), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n930), .A2(new_n925), .ZN(new_n950));
  AOI21_X1  g525(.A(G37), .B1(new_n950), .B2(new_n909), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT43), .B1(new_n951), .B2(new_n931), .ZN(new_n952));
  INV_X1    g527(.A(new_n944), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT44), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n933), .B1(new_n951), .B2(new_n931), .ZN(new_n955));
  INV_X1    g530(.A(new_n947), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n908), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT113), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n954), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n949), .A2(new_n959), .ZN(G397));
  INV_X1    g535(.A(G1384), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n961), .B1(new_n501), .B2(new_n507), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G40), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n486), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  XOR2_X1   g544(.A(new_n762), .B(G1996), .Z(new_n970));
  XNOR2_X1  g545(.A(new_n719), .B(G2067), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  XOR2_X1   g547(.A(new_n815), .B(new_n817), .Z(new_n973));
  XNOR2_X1  g548(.A(new_n973), .B(KEYINPUT114), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(G290), .B(G1986), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n969), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n963), .A2(G1384), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n978), .B1(new_n501), .B2(new_n507), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT117), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT117), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n981), .B(new_n978), .C1(new_n501), .C2(new_n507), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n964), .A2(new_n967), .ZN(new_n985));
  OAI211_X1 g560(.A(KEYINPUT118), .B(new_n772), .C1(new_n984), .C2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n962), .A2(KEYINPUT50), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT50), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n988), .B(new_n961), .C1(new_n501), .C2(new_n507), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n987), .A2(new_n967), .A3(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n990), .A2(G2084), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n986), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n772), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n482), .A2(G101), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(KEYINPUT69), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n482), .A2(new_n478), .A3(G101), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n998), .A2(G40), .A3(new_n477), .A4(new_n471), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n999), .B1(new_n963), .B2(new_n962), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n994), .B1(new_n1000), .B2(new_n983), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1001), .A2(KEYINPUT118), .ZN(new_n1002));
  OAI21_X1  g577(.A(G8), .B1(new_n993), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT51), .ZN(new_n1004));
  NAND2_X1  g579(.A1(G286), .A2(G8), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT122), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT122), .ZN(new_n1007));
  NAND3_X1  g582(.A1(G286), .A2(new_n1007), .A3(G8), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1003), .A2(new_n1004), .A3(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1009), .B1(new_n993), .B2(new_n1002), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT51), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n991), .B1(new_n1001), .B2(KEYINPUT118), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n772), .B1(new_n984), .B2(new_n985), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT118), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1014), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1009), .B1(new_n1018), .B2(G8), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1011), .B1(new_n1013), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT123), .ZN(new_n1021));
  INV_X1    g596(.A(G2078), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n964), .A2(new_n967), .A3(new_n1022), .A4(new_n979), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT53), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1024), .A2(G2078), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n983), .A2(new_n964), .A3(new_n967), .A4(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n990), .A2(new_n699), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1025), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(G171), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n964), .A2(new_n967), .A3(new_n979), .A4(new_n1026), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1025), .A2(new_n1028), .A3(G301), .A4(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT54), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n529), .A2(G8), .A3(new_n533), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n529), .A2(new_n533), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n987), .A2(new_n967), .A3(new_n989), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n964), .A2(new_n967), .A3(new_n979), .ZN(new_n1040));
  AOI22_X1  g615(.A1(new_n1039), .A2(new_n693), .B1(new_n1040), .B2(new_n799), .ZN(new_n1041));
  INV_X1    g616(.A(G8), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1038), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1044));
  AOI21_X1  g619(.A(G1971), .B1(new_n1000), .B2(new_n979), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n990), .A2(G2090), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1044), .B(G8), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G1981), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n584), .A2(new_n588), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n531), .B1(new_n585), .B2(new_n586), .ZN(new_n1050));
  OAI21_X1  g625(.A(G1981), .B1(new_n583), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT115), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1049), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(G305), .A2(KEYINPUT115), .A3(G1981), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT49), .ZN(new_n1056));
  OAI21_X1  g631(.A(G8), .B1(new_n999), .B2(new_n962), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT49), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1053), .A2(new_n1059), .A3(new_n1054), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1056), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n778), .A2(G1976), .A3(new_n780), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(KEYINPUT52), .B1(new_n1063), .B2(new_n1057), .ZN(new_n1064));
  OR2_X1    g639(.A1(new_n999), .A2(new_n962), .ZN(new_n1065));
  INV_X1    g640(.A(G1976), .ZN(new_n1066));
  AOI21_X1  g641(.A(KEYINPUT52), .B1(G288), .B2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1065), .A2(new_n1062), .A3(new_n1067), .A4(G8), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n1064), .A2(new_n1068), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1043), .A2(new_n1047), .A3(new_n1061), .A4(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1025), .A2(new_n1028), .A3(new_n1031), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(G171), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1025), .A2(new_n1027), .A3(new_n1028), .A4(G301), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1072), .A2(KEYINPUT54), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT124), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT124), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1072), .A2(new_n1076), .A3(KEYINPUT54), .A4(new_n1073), .ZN(new_n1077));
  AOI211_X1 g652(.A(new_n1033), .B(new_n1070), .C1(new_n1075), .C2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT123), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1079), .B(new_n1011), .C1(new_n1013), .C2(new_n1019), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1021), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT125), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1021), .A2(new_n1078), .A3(KEYINPUT125), .A4(new_n1080), .ZN(new_n1084));
  INV_X1    g659(.A(G1956), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n990), .A2(KEYINPUT119), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT119), .B1(new_n990), .B2(new_n1085), .ZN(new_n1087));
  XOR2_X1   g662(.A(KEYINPUT56), .B(G2072), .Z(new_n1088));
  OAI22_X1  g663(.A1(new_n1086), .A2(new_n1087), .B1(new_n1040), .B2(new_n1088), .ZN(new_n1089));
  XNOR2_X1  g664(.A(G299), .B(KEYINPUT57), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  OR2_X1    g666(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1092));
  OAI22_X1  g667(.A1(new_n1039), .A2(G1348), .B1(new_n1065), .B2(G2067), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1093), .A2(new_n614), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1092), .A2(KEYINPUT61), .A3(new_n1091), .ZN(new_n1096));
  OR2_X1    g671(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1097));
  XOR2_X1   g672(.A(KEYINPUT58), .B(G1341), .Z(new_n1098));
  NAND2_X1  g673(.A1(new_n1065), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT120), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1065), .A2(KEYINPUT120), .A3(new_n1098), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1101), .B(new_n1102), .C1(G1996), .C2(new_n1040), .ZN(new_n1103));
  AOI211_X1 g678(.A(new_n562), .B(new_n559), .C1(KEYINPUT121), .C2(KEYINPUT59), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1097), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NOR3_X1   g680(.A1(new_n1093), .A2(KEYINPUT60), .A3(new_n606), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1093), .A2(new_n614), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT60), .B1(new_n1094), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1103), .A2(new_n1097), .A3(new_n1104), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1096), .A2(new_n1107), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT61), .B1(new_n1092), .B2(new_n1091), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1091), .B(new_n1095), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n1083), .A2(new_n1084), .A3(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(G288), .A2(G1976), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1061), .A2(new_n1115), .B1(new_n1048), .B2(new_n790), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT116), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1058), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1061), .A2(new_n1069), .ZN(new_n1120));
  OAI22_X1  g695(.A1(new_n1118), .A2(new_n1119), .B1(new_n1047), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT63), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1018), .A2(G8), .A3(G168), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1122), .B1(new_n1123), .B2(new_n1070), .ZN(new_n1124));
  OR3_X1    g699(.A1(new_n1123), .A2(new_n1070), .A3(new_n1122), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1121), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1021), .A2(KEYINPUT62), .A3(new_n1080), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1070), .A2(new_n1030), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT62), .B1(new_n1021), .B2(new_n1080), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1126), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n977), .B1(new_n1114), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n975), .A2(new_n969), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n968), .A2(G290), .A3(G1986), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1134), .B(KEYINPUT126), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1133), .B1(KEYINPUT48), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1136), .B1(KEYINPUT48), .B2(new_n1135), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n968), .B1(new_n971), .B2(new_n763), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT46), .B1(new_n968), .B2(G1996), .ZN(new_n1139));
  OR3_X1    g714(.A1(new_n968), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1138), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n1141), .B(KEYINPUT47), .ZN(new_n1142));
  NOR3_X1   g717(.A1(new_n810), .A2(new_n814), .A3(new_n817), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n972), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(G2067), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n719), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n968), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n1137), .A2(new_n1142), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1132), .A2(new_n1148), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g724(.A1(G401), .A2(new_n462), .A3(G227), .ZN(new_n1151));
  NAND2_X1  g725(.A1(new_n1151), .A2(new_n688), .ZN(new_n1152));
  INV_X1    g726(.A(KEYINPUT127), .ZN(new_n1153));
  XNOR2_X1  g727(.A(new_n1152), .B(new_n1153), .ZN(new_n1154));
  NAND2_X1  g728(.A1(new_n946), .A2(new_n947), .ZN(new_n1155));
  NAND3_X1  g729(.A1(new_n1154), .A2(new_n865), .A3(new_n1155), .ZN(G225));
  INV_X1    g730(.A(G225), .ZN(G308));
endmodule


