//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 1 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 1 0 0 1 1 1 0 1 0 0 1 1 0 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1192, new_n1193, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  NAND2_X1  g0009(.A1(new_n202), .A2(new_n203), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G50), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT64), .ZN(new_n212));
  NAND3_X1  g0012(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT0), .ZN(new_n217));
  OAI22_X1  g0017(.A1(new_n212), .A2(new_n213), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT65), .Z(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G68), .A2(G238), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  AND2_X1   g0024(.A1(G50), .A2(G226), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n214), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT1), .ZN(new_n227));
  AOI211_X1 g0027(.A(new_n218), .B(new_n227), .C1(new_n217), .C2(new_n216), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G264), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(G270), .Z(new_n235));
  XOR2_X1   g0035(.A(new_n232), .B(new_n235), .Z(G358));
  XNOR2_X1  g0036(.A(G50), .B(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G58), .ZN(new_n238));
  INV_X1    g0038(.A(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G97), .B(G107), .ZN(new_n241));
  INV_X1    g0041(.A(G87), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  INV_X1    g0043(.A(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n240), .B(new_n245), .Z(G351));
  OAI21_X1  g0046(.A(KEYINPUT78), .B1(new_n202), .B2(new_n203), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT78), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n248), .A2(G58), .A3(G68), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n247), .A2(new_n249), .A3(new_n210), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  AOI22_X1  g0051(.A1(new_n250), .A2(G20), .B1(G159), .B2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT77), .ZN(new_n253));
  AND2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NOR3_X1   g0055(.A1(new_n254), .A2(new_n255), .A3(G20), .ZN(new_n256));
  XOR2_X1   g0056(.A(KEYINPUT76), .B(KEYINPUT7), .Z(new_n257));
  AOI21_X1  g0057(.A(new_n203), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT3), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G20), .ZN(new_n262));
  NAND2_X1  g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT7), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n253), .B1(new_n258), .B2(new_n265), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT76), .B(KEYINPUT7), .ZN(new_n267));
  OAI21_X1  g0067(.A(G68), .B1(new_n264), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT7), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n254), .A2(new_n255), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n269), .B1(new_n270), .B2(new_n262), .ZN(new_n271));
  NOR3_X1   g0071(.A1(new_n268), .A2(new_n271), .A3(KEYINPUT77), .ZN(new_n272));
  OAI211_X1 g0072(.A(KEYINPUT16), .B(new_n252), .C1(new_n266), .C2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(KEYINPUT67), .B1(new_n214), .B2(new_n260), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G1), .A2(G13), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT67), .ZN(new_n276));
  NAND4_X1  g0076(.A1(new_n276), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n274), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n261), .A2(new_n269), .A3(new_n262), .A4(new_n263), .ZN(new_n280));
  OAI211_X1 g0080(.A(G68), .B(new_n280), .C1(new_n256), .C2(new_n257), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n279), .B1(new_n252), .B2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(KEYINPUT80), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT80), .ZN(new_n284));
  AOI211_X1 g0084(.A(new_n284), .B(new_n279), .C1(new_n252), .C2(new_n281), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n273), .B(new_n278), .C1(new_n283), .C2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT68), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n278), .A2(new_n287), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n274), .A2(KEYINPUT68), .A3(new_n275), .A4(new_n277), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G1), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(G13), .A3(G20), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n292), .A2(G20), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n296), .B(KEYINPUT70), .ZN(new_n297));
  XNOR2_X1  g0097(.A(KEYINPUT8), .B(G58), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n295), .A2(new_n299), .B1(new_n294), .B2(new_n298), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n286), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G274), .ZN(new_n302));
  XNOR2_X1  g0102(.A(KEYINPUT66), .B(G45), .ZN(new_n303));
  INV_X1    g0103(.A(G41), .ZN(new_n304));
  AOI211_X1 g0104(.A(G1), .B(new_n302), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n261), .A2(new_n263), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n306), .A2(G226), .A3(G1698), .ZN(new_n307));
  NAND2_X1  g0107(.A1(G33), .A2(G87), .ZN(new_n308));
  INV_X1    g0108(.A(G1698), .ZN(new_n309));
  OAI211_X1 g0109(.A(G223), .B(new_n309), .C1(new_n254), .C2(new_n255), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n307), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n275), .B1(G33), .B2(G41), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n305), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G45), .ZN(new_n314));
  AOI21_X1  g0114(.A(G1), .B1(new_n304), .B2(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G232), .ZN(new_n317));
  AND3_X1   g0117(.A1(new_n313), .A2(G179), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G169), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n319), .B1(new_n313), .B2(new_n317), .ZN(new_n320));
  OR2_X1    g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n301), .A2(KEYINPUT18), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT81), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n318), .A2(new_n320), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n325), .B1(new_n286), .B2(new_n300), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n326), .A2(KEYINPUT81), .A3(KEYINPUT18), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n301), .A2(new_n321), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT18), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n324), .A2(new_n327), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n313), .A2(new_n317), .ZN(new_n332));
  INV_X1    g0132(.A(G200), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n334), .B1(G190), .B2(new_n332), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n335), .A2(new_n286), .A3(new_n300), .ZN(new_n336));
  XNOR2_X1  g0136(.A(new_n336), .B(KEYINPUT17), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n331), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(G1698), .B1(new_n261), .B2(new_n263), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n339), .A2(G222), .B1(new_n270), .B2(G77), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n309), .B1(new_n261), .B2(new_n263), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(G223), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n305), .B1(new_n343), .B2(new_n312), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n316), .A2(G226), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G190), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n348), .B1(G200), .B2(new_n346), .ZN(new_n349));
  NOR4_X1   g0149(.A1(new_n291), .A2(new_n201), .A3(new_n297), .A4(new_n294), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n204), .A2(G20), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT69), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n260), .A2(G20), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n298), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(KEYINPUT69), .B1(new_n204), .B2(G20), .ZN(new_n357));
  INV_X1    g0157(.A(new_n251), .ZN(new_n358));
  INV_X1    g0158(.A(G150), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR4_X1   g0160(.A1(new_n353), .A2(new_n356), .A3(new_n357), .A4(new_n360), .ZN(new_n361));
  OAI22_X1  g0161(.A1(new_n361), .A2(new_n290), .B1(G50), .B2(new_n293), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n350), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT9), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NOR3_X1   g0165(.A1(new_n350), .A2(new_n362), .A3(KEYINPUT9), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n349), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT10), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n346), .A2(G200), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n369), .B(KEYINPUT72), .C1(new_n347), .C2(new_n346), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n367), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  OAI221_X1 g0171(.A(new_n349), .B1(KEYINPUT72), .B2(KEYINPUT10), .C1(new_n365), .C2(new_n366), .ZN(new_n372));
  INV_X1    g0172(.A(new_n363), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n346), .A2(new_n319), .ZN(new_n374));
  INV_X1    g0174(.A(G179), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n344), .A2(new_n375), .A3(new_n345), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n373), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n371), .A2(new_n372), .A3(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n305), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n316), .A2(G244), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n341), .A2(G238), .B1(new_n270), .B2(G107), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n306), .A2(G232), .A3(new_n309), .ZN(new_n382));
  AND2_X1   g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI211_X1 g0183(.A(G1), .B(G13), .C1(new_n260), .C2(new_n304), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n379), .B(new_n380), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  OR2_X1    g0185(.A1(new_n385), .A2(G179), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n293), .A2(KEYINPUT71), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT71), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n388), .A2(new_n292), .A3(G13), .A4(G20), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NOR3_X1   g0190(.A1(new_n297), .A2(new_n390), .A3(new_n278), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(G77), .ZN(new_n392));
  OAI22_X1  g0192(.A1(new_n298), .A2(new_n358), .B1(new_n262), .B2(new_n239), .ZN(new_n393));
  XNOR2_X1  g0193(.A(KEYINPUT15), .B(G87), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n394), .A2(new_n355), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n278), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  AND2_X1   g0196(.A1(new_n387), .A2(new_n389), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n392), .B(new_n396), .C1(G77), .C2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n385), .A2(new_n319), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n386), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NOR3_X1   g0201(.A1(new_n338), .A2(new_n378), .A3(new_n401), .ZN(new_n402));
  OAI211_X1 g0202(.A(G226), .B(new_n309), .C1(new_n254), .C2(new_n255), .ZN(new_n403));
  OAI211_X1 g0203(.A(G232), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G97), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n406), .A2(new_n312), .B1(new_n316), .B2(G238), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n379), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT13), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT73), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT13), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n407), .A2(new_n411), .A3(new_n379), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n409), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n408), .A2(KEYINPUT73), .A3(KEYINPUT13), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(G179), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n409), .A2(new_n412), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT14), .B1(new_n417), .B2(new_n319), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n409), .A2(new_n412), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT14), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(new_n420), .A3(G169), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n416), .A2(new_n418), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT75), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n354), .A2(G77), .B1(new_n251), .B2(G50), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n262), .B2(G68), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n291), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g0227(.A(new_n427), .B(KEYINPUT11), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n391), .A2(G68), .ZN(new_n429));
  INV_X1    g0229(.A(G13), .ZN(new_n430));
  NOR3_X1   g0230(.A1(new_n430), .A2(KEYINPUT12), .A3(G1), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n431), .A2(G20), .A3(new_n203), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n397), .A2(G68), .ZN(new_n433));
  XOR2_X1   g0233(.A(KEYINPUT74), .B(KEYINPUT12), .Z(new_n434));
  OAI21_X1  g0234(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n428), .A2(new_n429), .A3(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n416), .A2(KEYINPUT75), .A3(new_n421), .A4(new_n418), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n424), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n417), .A2(new_n333), .ZN(new_n439));
  AOI211_X1 g0239(.A(new_n439), .B(new_n436), .C1(G190), .C2(new_n415), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n398), .B1(new_n385), .B2(G200), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(new_n347), .B2(new_n385), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n402), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n341), .A2(G244), .B1(G33), .B2(G116), .ZN(new_n447));
  AOI21_X1  g0247(.A(KEYINPUT83), .B1(new_n339), .B2(G238), .ZN(new_n448));
  OAI211_X1 g0248(.A(G238), .B(new_n309), .C1(new_n254), .C2(new_n255), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT83), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n447), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT84), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n449), .A2(new_n450), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n306), .A2(KEYINPUT83), .A3(G238), .A4(new_n309), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n457), .A2(KEYINPUT84), .A3(new_n447), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n454), .A2(new_n312), .A3(new_n458), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n384), .B(G250), .C1(G1), .C2(new_n314), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n314), .A2(G1), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G274), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n459), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n319), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n459), .A2(new_n375), .A3(new_n464), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT19), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n468), .B1(new_n355), .B2(new_n206), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n306), .A2(new_n262), .A3(G68), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n262), .B1(new_n405), .B2(new_n468), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n471), .B1(G87), .B2(new_n208), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n469), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n473), .A2(new_n278), .B1(new_n390), .B2(new_n394), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n260), .A2(G1), .ZN(new_n475));
  AOI211_X1 g0275(.A(new_n294), .B(new_n475), .C1(new_n288), .C2(new_n289), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n474), .B1(new_n477), .B2(new_n394), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n466), .A2(new_n467), .A3(new_n478), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n457), .A2(KEYINPUT84), .A3(new_n447), .ZN(new_n480));
  AOI21_X1  g0280(.A(KEYINPUT84), .B1(new_n457), .B2(new_n447), .ZN(new_n481));
  NOR3_X1   g0281(.A1(new_n480), .A2(new_n481), .A3(new_n384), .ZN(new_n482));
  OAI21_X1  g0282(.A(G200), .B1(new_n482), .B2(new_n463), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n476), .A2(G87), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n484), .A2(new_n474), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n459), .A2(G190), .A3(new_n464), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n483), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n479), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n341), .A2(G257), .ZN(new_n489));
  XNOR2_X1  g0289(.A(KEYINPUT89), .B(G294), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G33), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n306), .A2(G250), .A3(new_n309), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n489), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n312), .ZN(new_n494));
  XNOR2_X1  g0294(.A(KEYINPUT5), .B(G41), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n495), .A2(G274), .A3(new_n461), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n312), .B1(new_n461), .B2(new_n495), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G264), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n494), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n333), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n494), .A2(new_n347), .A3(new_n496), .A4(new_n498), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g0302(.A(KEYINPUT22), .B(G87), .C1(new_n254), .C2(new_n255), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G33), .A2(G116), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT22), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n262), .B(G87), .C1(new_n254), .C2(new_n255), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n505), .A2(new_n262), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT24), .ZN(new_n509));
  OAI21_X1  g0309(.A(KEYINPUT88), .B1(new_n262), .B2(G107), .ZN(new_n510));
  XNOR2_X1  g0310(.A(new_n510), .B(KEYINPUT23), .ZN(new_n511));
  AND3_X1   g0311(.A1(new_n508), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n509), .B1(new_n508), .B2(new_n511), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n278), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n476), .A2(G107), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n293), .A2(G107), .ZN(new_n516));
  XNOR2_X1  g0316(.A(new_n516), .B(KEYINPUT25), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n502), .A2(new_n514), .A3(new_n515), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n294), .A2(new_n206), .ZN(new_n519));
  XNOR2_X1  g0319(.A(KEYINPUT82), .B(KEYINPUT6), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n241), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NOR3_X1   g0322(.A1(new_n520), .A2(new_n206), .A3(G107), .ZN(new_n523));
  OAI21_X1  g0323(.A(G20), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n251), .A2(G77), .ZN(new_n525));
  OAI211_X1 g0325(.A(G107), .B(new_n280), .C1(new_n256), .C2(new_n257), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n278), .A2(new_n527), .B1(new_n476), .B2(G97), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n306), .A2(G244), .A3(new_n309), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT4), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(G33), .A2(G283), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n341), .A2(G250), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n339), .A2(KEYINPUT4), .A3(G244), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n531), .A2(new_n532), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n312), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n497), .A2(G257), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n496), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n536), .A2(new_n347), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(G200), .B1(new_n536), .B2(new_n539), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n519), .B(new_n528), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n527), .A2(new_n278), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n476), .A2(G97), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n543), .A2(new_n519), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n536), .A2(new_n539), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n319), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n538), .B1(new_n312), .B2(new_n535), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n375), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n545), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n518), .A2(new_n542), .A3(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n488), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n514), .A2(new_n515), .A3(new_n517), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n499), .A2(new_n319), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n494), .A2(new_n498), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n555), .A2(new_n375), .A3(new_n496), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n553), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n339), .A2(G257), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT85), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n270), .A2(G303), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n339), .A2(KEYINPUT85), .A3(G257), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n341), .A2(G264), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n560), .A2(new_n561), .A3(new_n562), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n312), .ZN(new_n565));
  INV_X1    g0365(.A(new_n496), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n566), .B1(new_n497), .B2(G270), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n319), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT86), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(new_n397), .B2(G116), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n390), .A2(KEYINPUT86), .A3(new_n244), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n390), .A2(new_n278), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n475), .A2(new_n244), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n570), .A2(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(G20), .B1(G33), .B2(G283), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n260), .A2(G97), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n575), .A2(new_n576), .B1(G20), .B2(new_n244), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n278), .A2(KEYINPUT20), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT20), .B1(new_n278), .B2(new_n577), .ZN(new_n579));
  OR2_X1    g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT87), .B1(new_n574), .B2(new_n580), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n274), .A2(new_n275), .A3(new_n277), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n397), .A2(new_n582), .A3(new_n573), .ZN(new_n583));
  AOI21_X1  g0383(.A(KEYINPUT86), .B1(new_n390), .B2(new_n244), .ZN(new_n584));
  AOI211_X1 g0384(.A(new_n569), .B(G116), .C1(new_n387), .C2(new_n389), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n578), .A2(new_n579), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT87), .ZN(new_n588));
  NOR3_X1   g0388(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n568), .B1(new_n581), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT21), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n568), .B(KEYINPUT21), .C1(new_n581), .C2(new_n589), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n565), .A2(new_n567), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n594), .A2(new_n375), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n581), .B2(new_n589), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n557), .A2(new_n592), .A3(new_n593), .A4(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n581), .A2(new_n589), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n565), .A2(new_n567), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(G190), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n594), .A2(G200), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n552), .A2(new_n598), .A3(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n446), .A2(new_n604), .ZN(G372));
  INV_X1    g0405(.A(new_n446), .ZN(new_n606));
  INV_X1    g0406(.A(new_n479), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n607), .B1(new_n552), .B2(new_n597), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n545), .A2(new_n547), .A3(new_n549), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n479), .A2(new_n487), .A3(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT26), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT90), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n479), .A2(new_n487), .A3(KEYINPUT26), .A4(new_n609), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n610), .A2(KEYINPUT90), .A3(new_n611), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n608), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n606), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g0418(.A(new_n618), .B(KEYINPUT91), .ZN(new_n619));
  INV_X1    g0419(.A(new_n377), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT17), .ZN(new_n621));
  XNOR2_X1  g0421(.A(new_n336), .B(new_n621), .ZN(new_n622));
  AOI211_X1 g0422(.A(new_n440), .B(new_n622), .C1(new_n438), .C2(new_n400), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n330), .A2(new_n322), .ZN(new_n624));
  OR2_X1    g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n371), .A2(new_n372), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n620), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n619), .A2(new_n627), .ZN(G369));
  INV_X1    g0428(.A(new_n603), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n592), .A2(new_n593), .A3(new_n596), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n430), .A2(G20), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n292), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(G213), .A3(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(G343), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n599), .A2(new_n638), .ZN(new_n639));
  OR2_X1    g0439(.A1(new_n630), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n630), .A2(new_n639), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n629), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(G330), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n553), .A2(new_n637), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n518), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n646), .A2(new_n557), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n557), .A2(new_n637), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n644), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n630), .A2(new_n638), .ZN(new_n651));
  OAI22_X1  g0451(.A1(new_n647), .A2(new_n651), .B1(new_n557), .B2(new_n637), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n650), .A2(new_n653), .ZN(G399));
  INV_X1    g0454(.A(new_n215), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n655), .A2(G41), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n208), .A2(G87), .A3(G116), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(G1), .A3(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n659), .B1(new_n212), .B2(new_n657), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n660), .B(KEYINPUT28), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT93), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n479), .A2(new_n487), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n518), .A2(new_n550), .A3(new_n542), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(new_n597), .A3(new_n664), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n665), .A2(new_n616), .A3(new_n479), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n637), .B1(new_n666), .B2(new_n615), .ZN(new_n667));
  XNOR2_X1  g0467(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n662), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n612), .A2(new_n614), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n608), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n671), .A2(KEYINPUT29), .A3(new_n638), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n617), .A2(new_n638), .ZN(new_n673));
  INV_X1    g0473(.A(new_n668), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(KEYINPUT93), .A3(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n669), .A2(new_n672), .A3(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n459), .A2(new_n548), .A3(new_n464), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n678), .A2(KEYINPUT30), .A3(new_n555), .A4(new_n595), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT30), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n600), .A2(G179), .A3(new_n555), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n680), .B1(new_n681), .B2(new_n677), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n600), .A2(G179), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n683), .A2(new_n546), .A3(new_n499), .A4(new_n465), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n679), .A2(new_n682), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n637), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT31), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n685), .A2(KEYINPUT31), .A3(new_n637), .ZN(new_n689));
  OAI211_X1 g0489(.A(new_n688), .B(new_n689), .C1(new_n604), .C2(new_n637), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G330), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n676), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n661), .B1(new_n693), .B2(G1), .ZN(G364));
  NAND3_X1  g0494(.A1(G355), .A2(new_n306), .A3(new_n215), .ZN(new_n695));
  INV_X1    g0495(.A(new_n303), .ZN(new_n696));
  OAI22_X1  g0496(.A1(new_n240), .A2(new_n314), .B1(new_n212), .B2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n655), .A2(new_n306), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  OAI221_X1 g0499(.A(new_n695), .B1(G116), .B2(new_n215), .C1(new_n697), .C2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(G13), .A2(G33), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(G20), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n275), .B1(G20), .B2(new_n319), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n700), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n704), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n347), .A2(G179), .A3(G200), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(new_n262), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(new_n206), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n262), .A2(new_n375), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(G200), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(G190), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n710), .B1(G68), .B2(new_n713), .ZN(new_n714));
  XOR2_X1   g0514(.A(new_n714), .B(KEYINPUT96), .Z(new_n715));
  NOR2_X1   g0515(.A1(new_n333), .A2(G179), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n716), .A2(G20), .A3(G190), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(G87), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n712), .A2(new_n347), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n262), .A2(G190), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(new_n375), .A3(new_n333), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G159), .ZN(new_n725));
  OAI22_X1  g0525(.A1(new_n721), .A2(new_n201), .B1(new_n725), .B2(KEYINPUT32), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n726), .B1(KEYINPUT32), .B2(new_n725), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n722), .A2(G179), .A3(new_n333), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n716), .A2(G20), .A3(new_n347), .ZN(new_n729));
  OAI221_X1 g0529(.A(new_n306), .B1(new_n728), .B2(new_n239), .C1(new_n207), .C2(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n711), .A2(G190), .A3(new_n333), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT95), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n711), .A2(KEYINPUT95), .A3(G190), .A4(new_n333), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n730), .B1(new_n736), .B2(G58), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n715), .A2(new_n719), .A3(new_n727), .A4(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n490), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n709), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n713), .ZN(new_n741));
  INV_X1    g0541(.A(G317), .ZN(new_n742));
  AND2_X1   g0542(.A1(new_n742), .A2(KEYINPUT33), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(KEYINPUT33), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n741), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  AOI211_X1 g0545(.A(new_n740), .B(new_n745), .C1(G326), .C2(new_n720), .ZN(new_n746));
  INV_X1    g0546(.A(new_n728), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G311), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n717), .B(KEYINPUT97), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G303), .ZN(new_n751));
  INV_X1    g0551(.A(G283), .ZN(new_n752));
  INV_X1    g0552(.A(G329), .ZN(new_n753));
  OAI221_X1 g0553(.A(new_n270), .B1(new_n729), .B2(new_n752), .C1(new_n753), .C2(new_n723), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n754), .B1(new_n736), .B2(G322), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n746), .A2(new_n748), .A3(new_n751), .A4(new_n755), .ZN(new_n756));
  AND2_X1   g0556(.A1(new_n738), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n703), .ZN(new_n758));
  OAI221_X1 g0558(.A(new_n706), .B1(new_n707), .B2(new_n757), .C1(new_n642), .C2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n631), .A2(G45), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n657), .A2(G1), .A3(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  OR3_X1    g0563(.A1(new_n642), .A2(KEYINPUT94), .A3(G330), .ZN(new_n764));
  OAI21_X1  g0564(.A(KEYINPUT94), .B1(new_n642), .B2(G330), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n644), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n763), .B1(new_n766), .B2(new_n762), .ZN(new_n767));
  XOR2_X1   g0567(.A(new_n767), .B(KEYINPUT98), .Z(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(G396));
  NAND2_X1  g0569(.A1(new_n398), .A2(new_n637), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n401), .B1(new_n445), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n400), .A2(new_n637), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n665), .A2(new_n616), .A3(new_n479), .ZN(new_n774));
  AND3_X1   g0574(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n638), .B(new_n773), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n773), .B1(new_n617), .B2(new_n638), .ZN(new_n778));
  OR3_X1    g0578(.A1(new_n777), .A2(new_n778), .A3(new_n691), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(new_n761), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(KEYINPUT101), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n691), .B1(new_n777), .B2(new_n778), .ZN(new_n782));
  INV_X1    g0582(.A(KEYINPUT101), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n779), .A2(new_n783), .A3(new_n761), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n781), .A2(new_n782), .A3(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n741), .A2(new_n752), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n710), .B(new_n786), .C1(G303), .C2(new_n720), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n724), .A2(G311), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n750), .A2(G107), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n270), .B1(new_n728), .B2(new_n244), .C1(new_n242), .C2(new_n729), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(new_n736), .B2(G294), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n787), .A2(new_n788), .A3(new_n789), .A4(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT99), .ZN(new_n793));
  AOI22_X1  g0593(.A1(G137), .A2(new_n720), .B1(new_n713), .B2(G150), .ZN(new_n794));
  INV_X1    g0594(.A(G159), .ZN(new_n795));
  INV_X1    g0595(.A(G143), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n794), .B1(new_n795), .B2(new_n728), .C1(new_n796), .C2(new_n735), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT34), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n709), .A2(new_n202), .B1(new_n729), .B2(new_n203), .ZN(new_n801));
  INV_X1    g0601(.A(G132), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n306), .B1(new_n802), .B2(new_n723), .C1(new_n749), .C2(new_n201), .ZN(new_n803));
  NOR4_X1   g0603(.A1(new_n799), .A2(new_n800), .A3(new_n801), .A4(new_n803), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n793), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n761), .B1(new_n805), .B2(new_n704), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n704), .A2(new_n701), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n806), .B1(G77), .B2(new_n808), .C1(new_n702), .C2(new_n773), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT100), .Z(new_n810));
  NAND2_X1  g0610(.A1(new_n785), .A2(new_n810), .ZN(G384));
  INV_X1    g0611(.A(new_n635), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n301), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n813), .B(new_n336), .C1(KEYINPUT103), .C2(new_n326), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n301), .A2(KEYINPUT103), .A3(new_n321), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT37), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(KEYINPUT105), .B1(new_n814), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n813), .A2(new_n336), .ZN(new_n819));
  OAI21_X1  g0619(.A(KEYINPUT37), .B1(new_n819), .B2(new_n326), .ZN(new_n820));
  INV_X1    g0620(.A(new_n336), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n635), .B1(new_n286), .B2(new_n300), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(KEYINPUT37), .B1(new_n326), .B2(KEYINPUT103), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT103), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n328), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT105), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n823), .A2(new_n824), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n818), .A2(new_n820), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n822), .B1(new_n624), .B2(new_n622), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT38), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n252), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n258), .A2(new_n253), .A3(new_n265), .ZN(new_n835));
  OAI21_X1  g0635(.A(KEYINPUT77), .B1(new_n268), .B2(new_n271), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n273), .B1(new_n837), .B2(new_n279), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n838), .A2(new_n290), .ZN(new_n839));
  INV_X1    g0639(.A(new_n300), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n812), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n338), .A2(new_n842), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n839), .A2(new_n840), .B1(new_n321), .B2(new_n812), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n816), .B1(new_n844), .B2(new_n336), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n817), .B2(new_n814), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n843), .A2(KEYINPUT38), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n833), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n436), .A2(new_n637), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n442), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n438), .A2(new_n441), .A3(new_n850), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n690), .A2(new_n773), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n849), .A2(KEYINPUT40), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  XOR2_X1   g0656(.A(KEYINPUT106), .B(KEYINPUT40), .Z(new_n857));
  AOI21_X1  g0657(.A(KEYINPUT38), .B1(new_n843), .B2(new_n847), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n841), .B1(new_n331), .B2(new_n337), .ZN(new_n859));
  AOI21_X1  g0659(.A(KEYINPUT103), .B1(new_n301), .B2(new_n321), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n819), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n845), .B1(new_n861), .B2(new_n824), .ZN(new_n862));
  NOR3_X1   g0662(.A1(new_n859), .A2(new_n862), .A3(new_n832), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n858), .A2(new_n863), .ZN(new_n864));
  AND3_X1   g0664(.A1(new_n438), .A2(new_n441), .A3(new_n850), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n850), .B1(new_n438), .B2(new_n441), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n690), .B(new_n773), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n857), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n856), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n606), .A2(new_n690), .ZN(new_n870));
  XOR2_X1   g0670(.A(new_n869), .B(new_n870), .Z(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(G330), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n669), .A2(new_n606), .A3(new_n672), .A4(new_n675), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n627), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n872), .B(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n772), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n776), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n832), .B1(new_n859), .B2(new_n862), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n848), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n877), .A2(new_n879), .A3(new_n854), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n624), .A2(new_n635), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n424), .A2(new_n437), .A3(new_n436), .A4(new_n638), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT104), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT39), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n833), .A2(new_n886), .A3(new_n848), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT39), .B1(new_n858), .B2(new_n863), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n885), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n882), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n875), .B(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(new_n292), .B2(new_n631), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n522), .A2(new_n523), .ZN(new_n893));
  XOR2_X1   g0693(.A(new_n893), .B(KEYINPUT102), .Z(new_n894));
  INV_X1    g0694(.A(KEYINPUT35), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n213), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n896), .B(G116), .C1(new_n895), .C2(new_n894), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n897), .B(KEYINPUT36), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n247), .A2(new_n249), .A3(G77), .ZN(new_n899));
  OAI22_X1  g0699(.A1(new_n212), .A2(new_n899), .B1(G50), .B2(new_n203), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n900), .A2(G1), .A3(new_n430), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n892), .A2(new_n898), .A3(new_n901), .ZN(G367));
  OAI221_X1 g0702(.A(new_n705), .B1(new_n215), .B2(new_n394), .C1(new_n235), .C2(new_n699), .ZN(new_n903));
  OAI22_X1  g0703(.A1(new_n741), .A2(new_n795), .B1(new_n203), .B2(new_n709), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(G143), .B2(new_n720), .ZN(new_n905));
  INV_X1    g0705(.A(G137), .ZN(new_n906));
  OAI22_X1  g0706(.A1(new_n723), .A2(new_n906), .B1(new_n728), .B2(new_n201), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n736), .B2(G150), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n718), .A2(G58), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n306), .B1(new_n729), .B2(new_n239), .ZN(new_n910));
  XOR2_X1   g0710(.A(new_n910), .B(KEYINPUT110), .Z(new_n911));
  NAND4_X1  g0711(.A1(new_n905), .A2(new_n908), .A3(new_n909), .A4(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT46), .B1(new_n718), .B2(G116), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n741), .A2(new_n739), .B1(new_n207), .B2(new_n709), .ZN(new_n914));
  AOI211_X1 g0714(.A(new_n913), .B(new_n914), .C1(G311), .C2(new_n720), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n750), .A2(KEYINPUT46), .A3(G116), .ZN(new_n916));
  OAI221_X1 g0716(.A(new_n270), .B1(new_n728), .B2(new_n752), .C1(new_n206), .C2(new_n729), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n917), .B1(new_n736), .B2(G303), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n915), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n723), .A2(new_n742), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n912), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n921), .B(KEYINPUT47), .Z(new_n922));
  OAI211_X1 g0722(.A(new_n762), .B(new_n903), .C1(new_n922), .C2(new_n707), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT111), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n485), .A2(new_n638), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n663), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n479), .B2(new_n925), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n927), .A2(new_n758), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n924), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n651), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n609), .A2(new_n637), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n545), .A2(new_n637), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n542), .A2(new_n550), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n649), .A2(new_n930), .A3(new_n934), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n935), .B(KEYINPUT42), .Z(new_n936));
  OAI21_X1  g0736(.A(new_n550), .B1(new_n933), .B2(new_n557), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n638), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n936), .A2(new_n938), .B1(KEYINPUT43), .B2(new_n927), .ZN(new_n939));
  INV_X1    g0739(.A(new_n934), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n650), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n939), .B(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n927), .A2(KEYINPUT43), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n942), .B(new_n943), .Z(new_n944));
  XOR2_X1   g0744(.A(KEYINPUT107), .B(KEYINPUT41), .Z(new_n945));
  XOR2_X1   g0745(.A(new_n656), .B(new_n945), .Z(new_n946));
  NAND2_X1  g0746(.A1(new_n652), .A2(new_n940), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT44), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n947), .B(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n653), .A2(KEYINPUT45), .A3(new_n934), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT45), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n652), .B2(new_n940), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n949), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n650), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n949), .A2(new_n953), .A3(new_n650), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n649), .B(new_n930), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(new_n644), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n676), .A2(new_n960), .A3(new_n691), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(KEYINPUT108), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT108), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n676), .A2(new_n960), .A3(new_n963), .A4(new_n691), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n958), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n946), .B1(new_n965), .B2(new_n692), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n760), .A2(G1), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT109), .Z(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n929), .B1(new_n944), .B2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(G387));
  INV_X1    g0772(.A(new_n960), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n692), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n974), .A2(new_n656), .A3(new_n961), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n960), .A2(new_n968), .ZN(new_n976));
  AOI22_X1  g0776(.A1(G311), .A2(new_n713), .B1(new_n720), .B2(G322), .ZN(new_n977));
  INV_X1    g0777(.A(G303), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n977), .B1(new_n978), .B2(new_n728), .C1(new_n742), .C2(new_n735), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT48), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n980), .B1(new_n752), .B2(new_n709), .C1(new_n739), .C2(new_n717), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT49), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n724), .A2(G326), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n981), .A2(new_n982), .ZN(new_n985));
  INV_X1    g0785(.A(new_n729), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n306), .B1(new_n986), .B2(G116), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n983), .A2(new_n984), .A3(new_n985), .A4(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n723), .A2(new_n359), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n795), .A2(new_n721), .B1(new_n741), .B2(new_n298), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n709), .A2(new_n394), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n717), .A2(new_n239), .B1(new_n728), .B2(new_n203), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(new_n736), .B2(G50), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n270), .B1(new_n986), .B2(G97), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n992), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n988), .B1(new_n989), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n658), .B1(new_n203), .B2(new_n239), .ZN(new_n998));
  NOR3_X1   g0798(.A1(new_n298), .A2(KEYINPUT50), .A3(G50), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(KEYINPUT50), .B1(new_n298), .B2(G50), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n1000), .A2(new_n314), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n699), .B1(new_n232), .B2(new_n696), .ZN(new_n1003));
  NOR3_X1   g0803(.A1(new_n658), .A2(new_n655), .A3(new_n270), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1002), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(G107), .B2(new_n215), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n997), .A2(new_n704), .B1(new_n705), .B2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1007), .B(new_n762), .C1(new_n649), .C2(new_n758), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT112), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n975), .A2(new_n976), .A3(new_n1009), .ZN(G393));
  AND2_X1   g0810(.A1(new_n958), .A2(new_n961), .ZN(new_n1011));
  NOR3_X1   g0811(.A1(new_n965), .A2(new_n657), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT113), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n958), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n956), .A2(KEYINPUT113), .A3(new_n957), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1014), .A2(new_n968), .A3(new_n1015), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n736), .A2(G159), .B1(G150), .B2(new_n720), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1017), .A2(KEYINPUT51), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n203), .A2(new_n717), .B1(new_n723), .B2(new_n796), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n298), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1019), .B1(new_n1020), .B2(new_n747), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n239), .B2(new_n709), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1018), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1017), .A2(KEYINPUT51), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n713), .A2(G50), .B1(new_n986), .B2(G87), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1023), .A2(new_n306), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(G294), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n728), .A2(new_n1027), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n736), .A2(G311), .B1(G317), .B2(new_n720), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1029), .A2(KEYINPUT52), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(KEYINPUT52), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n741), .A2(new_n978), .B1(new_n207), .B2(new_n729), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n270), .B1(new_n709), .B2(new_n244), .ZN(new_n1033));
  INV_X1    g0833(.A(G322), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n752), .A2(new_n717), .B1(new_n723), .B2(new_n1034), .ZN(new_n1035));
  NOR3_X1   g0835(.A1(new_n1032), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1030), .A2(new_n1031), .A3(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1026), .B1(new_n1028), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n761), .B1(new_n1038), .B2(new_n704), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n245), .A2(new_n698), .B1(G97), .B2(new_n655), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n705), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1039), .B(new_n1041), .C1(new_n758), .C2(new_n934), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1016), .A2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1012), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(G390));
  AOI22_X1  g0845(.A1(new_n776), .A2(new_n876), .B1(new_n853), .B2(new_n852), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n887), .B(new_n888), .C1(new_n1046), .C2(new_n884), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n637), .B(new_n771), .C1(new_n608), .C2(new_n670), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n854), .B1(new_n1048), .B2(new_n772), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1049), .A2(new_n849), .A3(new_n885), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n854), .A2(G330), .A3(new_n690), .A4(new_n773), .ZN(new_n1051));
  AND3_X1   g0851(.A1(new_n1047), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1051), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n690), .A2(G330), .A3(new_n773), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n865), .A2(new_n866), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1048), .A2(new_n772), .ZN(new_n1057));
  AND3_X1   g0857(.A1(new_n1051), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n1051), .A2(new_n1056), .B1(new_n876), .B2(new_n776), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n606), .A2(G330), .A3(new_n690), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n873), .A2(new_n627), .A3(new_n1061), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n1052), .A2(new_n1053), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n887), .A2(new_n888), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n884), .B1(new_n877), .B2(new_n854), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1050), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1051), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1047), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1069));
  AND3_X1   g0869(.A1(new_n873), .A2(new_n627), .A3(new_n1061), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1051), .A2(new_n1056), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n877), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1051), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .A4(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1063), .A2(new_n1075), .A3(new_n656), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1064), .A2(new_n702), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n808), .A2(new_n1020), .ZN(new_n1078));
  XOR2_X1   g0878(.A(KEYINPUT54), .B(G143), .Z(new_n1079));
  AOI22_X1  g0879(.A1(new_n713), .A2(G137), .B1(new_n747), .B2(new_n1079), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT114), .Z(new_n1081));
  INV_X1    g0881(.A(new_n709), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1081), .B1(G159), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(G128), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n735), .A2(new_n802), .B1(new_n1084), .B2(new_n721), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT116), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n717), .A2(new_n359), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT53), .ZN(new_n1088));
  INV_X1    g0888(.A(G125), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n306), .B1(new_n729), .B2(new_n201), .C1(new_n1089), .C2(new_n723), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT115), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1083), .A2(new_n1086), .A3(new_n1088), .A4(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT117), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n741), .A2(new_n207), .B1(new_n721), .B2(new_n752), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(G77), .B2(new_n1082), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(G116), .A2(new_n736), .B1(new_n750), .B2(G87), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n306), .B1(new_n747), .B2(G97), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n723), .A2(new_n1027), .B1(new_n729), .B2(new_n203), .ZN(new_n1098));
  XOR2_X1   g0898(.A(new_n1098), .B(KEYINPUT118), .Z(new_n1099));
  NAND4_X1  g0899(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .A4(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n707), .B1(new_n1093), .B2(new_n1100), .ZN(new_n1101));
  NOR4_X1   g0901(.A1(new_n1077), .A2(new_n761), .A3(new_n1078), .A4(new_n1101), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1102), .B1(new_n1103), .B2(new_n968), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n1076), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(G378));
  INV_X1    g0906(.A(KEYINPUT57), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1062), .B1(new_n1103), .B2(new_n1074), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n856), .A2(new_n868), .A3(G330), .ZN(new_n1109));
  AOI21_X1  g0909(.A(KEYINPUT38), .B1(new_n829), .B2(new_n830), .ZN(new_n1110));
  NOR3_X1   g0910(.A1(new_n1110), .A2(new_n863), .A3(KEYINPUT39), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n886), .B1(new_n848), .B2(new_n878), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n884), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1046), .A2(new_n879), .B1(new_n624), .B2(new_n635), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n378), .B(KEYINPUT119), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n363), .A2(new_n635), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1116), .B(new_n1117), .ZN(new_n1118));
  XOR2_X1   g0918(.A(new_n1115), .B(new_n1118), .Z(new_n1119));
  AND3_X1   g0919(.A1(new_n1113), .A2(new_n1114), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1119), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1109), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1115), .B(new_n1118), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n882), .B2(new_n889), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n856), .A2(new_n868), .A3(G330), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1113), .A2(new_n1114), .A3(new_n1119), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1122), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1107), .B1(new_n1108), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1075), .A2(new_n1070), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1130), .A2(KEYINPUT57), .A3(new_n1127), .A4(new_n1122), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1129), .A2(new_n656), .A3(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1122), .A2(new_n968), .A3(new_n1127), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n721), .A2(new_n1089), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n741), .A2(new_n802), .B1(new_n359), .B2(new_n709), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n1134), .B(new_n1135), .C1(new_n718), .C2(new_n1079), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n1136), .B1(new_n1084), .B2(new_n735), .C1(new_n906), .C2(new_n728), .ZN(new_n1137));
  XOR2_X1   g0937(.A(new_n1137), .B(KEYINPUT59), .Z(new_n1138));
  AOI21_X1  g0938(.A(G41), .B1(new_n724), .B2(G124), .ZN(new_n1139));
  AOI21_X1  g0939(.A(G33), .B1(new_n986), .B2(G159), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n201), .B1(new_n254), .B2(G41), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n304), .B(new_n270), .C1(new_n717), .C2(new_n239), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n741), .A2(new_n206), .B1(new_n721), .B2(new_n244), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1143), .B(new_n1144), .C1(G68), .C2(new_n1082), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n723), .A2(new_n752), .B1(new_n729), .B2(new_n202), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(new_n736), .B2(G107), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1145), .B(new_n1147), .C1(new_n394), .C2(new_n728), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1148), .B(KEYINPUT58), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1141), .A2(new_n1142), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n761), .B1(new_n1150), .B2(new_n704), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n1151), .B1(G50), .B2(new_n808), .C1(new_n1123), .C2(new_n702), .ZN(new_n1152));
  AND2_X1   g0952(.A1(new_n1133), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1132), .A2(new_n1153), .ZN(G375));
  NAND2_X1  g0954(.A1(new_n1070), .A2(new_n1074), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1155), .A2(new_n1156), .A3(new_n946), .ZN(new_n1157));
  XOR2_X1   g0957(.A(new_n1157), .B(KEYINPUT120), .Z(new_n1158));
  NOR2_X1   g0958(.A1(new_n741), .A2(new_n244), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n991), .B(new_n1159), .C1(G294), .C2(new_n720), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n270), .B1(new_n728), .B2(new_n207), .C1(new_n239), .C2(new_n729), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n750), .B2(G97), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n724), .A2(G303), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n736), .A2(G283), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1160), .A2(new_n1162), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(G137), .A2(new_n736), .B1(new_n750), .B2(G159), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n721), .A2(new_n802), .B1(new_n723), .B2(new_n1084), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(new_n713), .B2(new_n1079), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n709), .A2(new_n201), .B1(new_n728), .B2(new_n359), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT121), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n306), .B1(new_n729), .B2(new_n202), .ZN(new_n1171));
  XOR2_X1   g0971(.A(new_n1171), .B(KEYINPUT122), .Z(new_n1172));
  NAND4_X1  g0972(.A1(new_n1166), .A2(new_n1168), .A3(new_n1170), .A4(new_n1172), .ZN(new_n1173));
  AND2_X1   g0973(.A1(new_n1165), .A2(new_n1173), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n762), .B1(G68), .B2(new_n808), .C1(new_n1174), .C2(new_n707), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT123), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n1055), .B2(new_n701), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n1074), .B2(new_n968), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1158), .A2(new_n1178), .ZN(G381));
  NOR2_X1   g0979(.A1(G381), .A2(G390), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n768), .A2(new_n975), .A3(new_n976), .A4(new_n1009), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1181), .A2(G384), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT124), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1076), .A2(new_n1133), .A3(new_n1104), .A4(new_n1152), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1125), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n1130), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n657), .B1(new_n1188), .B2(new_n1107), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1184), .B1(new_n1189), .B2(new_n1131), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1180), .A2(new_n971), .A3(new_n1183), .A4(new_n1190), .ZN(G407));
  INV_X1    g0991(.A(G213), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n1190), .B2(new_n636), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(G407), .A2(new_n1193), .ZN(G409));
  NAND2_X1  g0994(.A1(G393), .A2(G396), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n1181), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1044), .A2(new_n1196), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1195), .B(new_n1181), .C1(new_n1012), .C2(new_n1043), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(G387), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n971), .A2(new_n1198), .A3(new_n1197), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT60), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n1070), .B2(new_n1074), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1060), .A2(new_n1062), .A3(KEYINPUT60), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1204), .A2(new_n656), .A3(new_n1155), .A4(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1206), .A2(G384), .A3(new_n1178), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(KEYINPUT126), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1206), .A2(new_n1178), .ZN(new_n1209));
  INV_X1    g1009(.A(G384), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT126), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1206), .A2(new_n1212), .A3(G384), .A4(new_n1178), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1208), .A2(new_n1211), .A3(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1192), .A2(G343), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(G2897), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1214), .A2(new_n1217), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1208), .A2(new_n1211), .A3(new_n1213), .A4(new_n1216), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1215), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1187), .A2(KEYINPUT125), .A3(new_n1130), .A4(new_n946), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1105), .A2(new_n1153), .A3(new_n1221), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1108), .A2(new_n1128), .ZN(new_n1223));
  AOI21_X1  g1023(.A(KEYINPUT125), .B1(new_n1223), .B2(new_n946), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1220), .B1(new_n1222), .B2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1105), .B1(new_n1132), .B2(new_n1153), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1218), .B(new_n1219), .C1(new_n1225), .C2(new_n1226), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(new_n1225), .A2(new_n1226), .A3(new_n1214), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT62), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1227), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n946), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(new_n1108), .A2(new_n1128), .A3(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1184), .B1(KEYINPUT125), .B2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT125), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n1188), .B2(new_n1231), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1215), .B1(new_n1233), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(G375), .A2(G378), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1214), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1236), .A2(new_n1237), .A3(new_n1229), .A4(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT61), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1202), .B1(new_n1230), .B2(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1200), .A2(new_n1240), .A3(new_n1201), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n1228), .B2(KEYINPUT63), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT63), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1235), .A2(new_n1105), .A3(new_n1153), .A4(new_n1221), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1153), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(new_n1189), .B2(new_n1131), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1220), .B(new_n1247), .C1(new_n1249), .C2(new_n1105), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1245), .B1(new_n1246), .B2(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1244), .B1(new_n1251), .B2(new_n1228), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1242), .A2(new_n1252), .ZN(G405));
  NOR2_X1   g1053(.A1(new_n1214), .A2(KEYINPUT127), .ZN(new_n1254));
  OR3_X1    g1054(.A1(new_n1254), .A2(new_n1190), .A3(new_n1226), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1202), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1254), .B1(new_n1190), .B2(new_n1226), .ZN(new_n1257));
  AND3_X1   g1057(.A1(new_n1255), .A2(new_n1256), .A3(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1256), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1258), .A2(new_n1259), .ZN(G402));
endmodule


