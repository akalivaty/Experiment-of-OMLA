//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 0 0 1 1 1 1 1 0 0 1 0 0 0 1 0 1 1 0 0 0 0 0 1 1 1 0 0 1 0 0 1 0 1 0 0 1 0 1 1 1 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT74), .ZN(new_n189));
  INV_X1    g003(.A(G104), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT74), .A2(G104), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(G107), .A3(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G107), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n194), .B1(new_n190), .B2(KEYINPUT3), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n191), .A2(new_n194), .A3(new_n192), .ZN(new_n197));
  AND3_X1   g011(.A1(new_n197), .A2(KEYINPUT75), .A3(KEYINPUT3), .ZN(new_n198));
  AOI21_X1  g012(.A(KEYINPUT75), .B1(new_n197), .B2(KEYINPUT3), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n196), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G101), .ZN(new_n201));
  INV_X1    g015(.A(G101), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n202), .B(new_n196), .C1(new_n198), .C2(new_n199), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n201), .A2(KEYINPUT4), .A3(new_n203), .ZN(new_n204));
  XOR2_X1   g018(.A(KEYINPUT2), .B(G113), .Z(new_n205));
  XNOR2_X1  g019(.A(G116), .B(G119), .ZN(new_n206));
  XNOR2_X1  g020(.A(new_n205), .B(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT4), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n200), .A2(new_n208), .A3(G101), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n204), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT76), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n211), .B1(new_n194), .B2(G104), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n190), .A2(KEYINPUT76), .A3(G107), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n197), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT77), .ZN(new_n215));
  AND3_X1   g029(.A1(new_n214), .A2(new_n215), .A3(G101), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n215), .B1(new_n214), .B2(G101), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n205), .A2(new_n206), .ZN(new_n219));
  INV_X1    g033(.A(G116), .ZN(new_n220));
  NOR3_X1   g034(.A1(new_n220), .A2(KEYINPUT5), .A3(G119), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n221), .B1(new_n206), .B2(KEYINPUT5), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n219), .B1(G113), .B2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n218), .A2(new_n203), .A3(new_n223), .ZN(new_n224));
  XOR2_X1   g038(.A(G110), .B(G122), .Z(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n210), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G146), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G143), .ZN(new_n229));
  INV_X1    g043(.A(G143), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G146), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT0), .ZN(new_n233));
  INV_X1    g047(.A(G128), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NOR2_X1   g049(.A1(KEYINPUT0), .A2(G128), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n232), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  XNOR2_X1  g051(.A(G143), .B(G146), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n238), .B1(new_n233), .B2(new_n234), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G125), .ZN(new_n241));
  NOR3_X1   g055(.A1(new_n232), .A2(KEYINPUT1), .A3(new_n234), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT64), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT64), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n245), .B(KEYINPUT1), .C1(new_n230), .C2(G146), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n244), .A2(G128), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n242), .B1(new_n247), .B2(new_n232), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n241), .B1(new_n248), .B2(G125), .ZN(new_n249));
  INV_X1    g063(.A(G953), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G224), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT7), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n249), .B(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n218), .A2(new_n203), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n254), .B(new_n223), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n225), .B(KEYINPUT8), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n227), .B(new_n253), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G902), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n210), .A2(new_n224), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(new_n225), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n261), .A2(KEYINPUT6), .A3(new_n227), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n249), .B(new_n251), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT6), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n260), .A2(new_n264), .A3(new_n225), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n262), .A2(new_n263), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT80), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n262), .A2(KEYINPUT80), .A3(new_n263), .A4(new_n265), .ZN(new_n269));
  AOI211_X1 g083(.A(new_n188), .B(new_n259), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT81), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n268), .A2(new_n269), .ZN(new_n272));
  INV_X1    g086(.A(new_n259), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n188), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT81), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n272), .A2(new_n187), .A3(new_n273), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G475), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT18), .ZN(new_n280));
  INV_X1    g094(.A(G131), .ZN(new_n281));
  INV_X1    g095(.A(G237), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT66), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT66), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G237), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(KEYINPUT67), .B(G953), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n287), .A3(G214), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n230), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n286), .A2(new_n287), .A3(G143), .A4(G214), .ZN(new_n290));
  AOI211_X1 g104(.A(new_n280), .B(new_n281), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(KEYINPUT18), .A2(G131), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n289), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G125), .ZN(new_n294));
  INV_X1    g108(.A(G140), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(G125), .A2(G140), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n296), .A2(KEYINPUT83), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(KEYINPUT83), .B1(new_n296), .B2(new_n297), .ZN(new_n299));
  OAI21_X1  g113(.A(G146), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n296), .A2(new_n297), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n228), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n293), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(KEYINPUT84), .B1(new_n291), .B2(new_n304), .ZN(new_n305));
  OR2_X1    g119(.A1(KEYINPUT67), .A2(G953), .ZN(new_n306));
  NAND2_X1  g120(.A1(KEYINPUT67), .A2(G953), .ZN(new_n307));
  AOI22_X1  g121(.A1(new_n283), .A2(new_n285), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(G143), .B1(new_n308), .B2(G214), .ZN(new_n309));
  INV_X1    g123(.A(new_n290), .ZN(new_n310));
  OAI211_X1 g124(.A(KEYINPUT18), .B(G131), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT84), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n311), .A2(new_n312), .A3(new_n293), .A4(new_n303), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n305), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(G131), .B1(new_n309), .B2(new_n310), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT17), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n289), .A2(new_n281), .A3(new_n290), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NOR3_X1   g132(.A1(new_n294), .A2(KEYINPUT16), .A3(G140), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n319), .B1(new_n301), .B2(KEYINPUT16), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n320), .A2(G146), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n320), .A2(G146), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n318), .B(new_n323), .C1(new_n316), .C2(new_n315), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n314), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(G113), .B(G122), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n326), .B(new_n190), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n314), .A2(new_n327), .A3(new_n324), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n279), .B1(new_n331), .B2(new_n258), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT19), .B1(new_n296), .B2(new_n297), .ZN(new_n333));
  OR2_X1    g147(.A1(new_n298), .A2(new_n299), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n333), .B1(new_n334), .B2(KEYINPUT19), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n321), .B1(new_n335), .B2(new_n228), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n315), .A2(new_n317), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n314), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(KEYINPUT85), .A3(new_n328), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT85), .ZN(new_n341));
  AOI22_X1  g155(.A1(new_n305), .A2(new_n313), .B1(new_n337), .B2(new_n336), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n341), .B1(new_n342), .B2(new_n327), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n340), .A2(new_n343), .A3(new_n330), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(new_n279), .A3(new_n258), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT82), .B(KEYINPUT20), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT20), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n344), .A2(new_n348), .A3(new_n279), .A4(new_n258), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n332), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT90), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n230), .A2(G128), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT13), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n230), .A2(G128), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n356), .B(KEYINPUT86), .C1(new_n354), .C2(new_n355), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n357), .B(G134), .C1(KEYINPUT86), .C2(new_n356), .ZN(new_n358));
  OR2_X1    g172(.A1(new_n358), .A2(KEYINPUT87), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n234), .A2(G143), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n355), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n361), .B(KEYINPUT88), .ZN(new_n362));
  INV_X1    g176(.A(G134), .ZN(new_n363));
  AND2_X1   g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(G116), .B(G122), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n194), .ZN(new_n366));
  INV_X1    g180(.A(new_n365), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G107), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n364), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n358), .A2(KEYINPUT87), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n359), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  XOR2_X1   g185(.A(KEYINPUT9), .B(G234), .Z(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G217), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n373), .A2(new_n374), .A3(G953), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n220), .A2(KEYINPUT14), .A3(G122), .ZN(new_n376));
  OAI211_X1 g190(.A(G107), .B(new_n376), .C1(new_n367), .C2(KEYINPUT14), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n366), .B(KEYINPUT89), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n362), .A2(new_n363), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n377), .B(new_n378), .C1(new_n364), .C2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n371), .A2(new_n375), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n375), .B1(new_n371), .B2(new_n380), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n352), .B(new_n258), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G478), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n385), .A2(KEYINPUT15), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n384), .B(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n351), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G952), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n389), .A2(G953), .ZN(new_n390));
  INV_X1    g204(.A(G234), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n390), .B1(new_n391), .B2(new_n282), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n287), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n394), .B(G902), .C1(new_n391), .C2(new_n282), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n395), .B(KEYINPUT91), .ZN(new_n396));
  XNOR2_X1  g210(.A(KEYINPUT21), .B(G898), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n393), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(G214), .B1(G237), .B2(G902), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  AND4_X1   g215(.A1(new_n271), .A2(new_n278), .A3(new_n388), .A4(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G137), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n287), .A2(G221), .A3(G234), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT72), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n404), .B(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT22), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n404), .B(KEYINPUT72), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n409), .A2(KEYINPUT22), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n403), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(KEYINPUT22), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n406), .A2(new_n407), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n412), .A2(new_n413), .A3(G137), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n234), .A2(G119), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT23), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OR2_X1    g232(.A1(new_n234), .A2(G119), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n234), .A2(KEYINPUT23), .A3(G119), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G110), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n422), .B(KEYINPUT69), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n419), .A2(new_n416), .ZN(new_n424));
  XNOR2_X1  g238(.A(KEYINPUT24), .B(G110), .ZN(new_n425));
  OAI22_X1  g239(.A1(new_n321), .A2(new_n322), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT70), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(KEYINPUT70), .B1(new_n423), .B2(new_n426), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n321), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n424), .A2(new_n425), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n433), .B1(new_n421), .B2(G110), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n432), .A2(new_n302), .A3(new_n434), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(KEYINPUT71), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n415), .A2(new_n431), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n415), .B1(new_n431), .B2(new_n436), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n258), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(KEYINPUT25), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n374), .B1(G234), .B2(new_n258), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n431), .A2(new_n436), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n411), .A2(new_n414), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n437), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT25), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(new_n447), .A3(new_n258), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n441), .A2(new_n442), .A3(new_n448), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n442), .A2(G902), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n450), .B(KEYINPUT73), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n446), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT32), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n205), .A2(new_n206), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n219), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT11), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n457), .B1(new_n363), .B2(G137), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n363), .A2(G137), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n403), .A2(KEYINPUT11), .A3(G134), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G131), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n458), .A2(new_n460), .A3(new_n281), .A4(new_n459), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n240), .ZN(new_n465));
  INV_X1    g279(.A(new_n459), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n363), .A2(G137), .ZN(new_n467));
  OAI21_X1  g281(.A(G131), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n463), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n456), .B(new_n465), .C1(new_n248), .C2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT65), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n246), .A2(G128), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n245), .B1(new_n229), .B2(KEYINPUT1), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n232), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT1), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n238), .A2(new_n476), .A3(G128), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n469), .ZN(new_n479));
  AOI22_X1  g293(.A1(new_n478), .A2(new_n479), .B1(new_n464), .B2(new_n240), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n480), .A2(KEYINPUT65), .A3(new_n456), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n472), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n465), .B1(new_n248), .B2(new_n469), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n483), .A2(KEYINPUT30), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT30), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n480), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n207), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n488), .B(G101), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n308), .A2(G210), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n489), .B(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(KEYINPUT68), .B(KEYINPUT31), .ZN(new_n492));
  AND4_X1   g306(.A1(new_n482), .A2(new_n487), .A3(new_n491), .A4(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT28), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n470), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n480), .A2(new_n456), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n497), .B1(new_n472), .B2(new_n481), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n496), .B1(new_n498), .B2(new_n495), .ZN(new_n499));
  INV_X1    g313(.A(new_n491), .ZN(new_n500));
  AOI21_X1  g314(.A(KEYINPUT31), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n487), .A2(new_n482), .A3(new_n491), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n494), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(G472), .A2(G902), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n454), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n503), .A2(new_n454), .A3(new_n504), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n499), .A2(new_n500), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT29), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT29), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n487), .A2(new_n482), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n511), .B1(new_n512), .B2(new_n491), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n510), .B(new_n258), .C1(new_n509), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(G472), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n453), .B1(new_n508), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(G221), .B1(new_n373), .B2(G902), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(G469), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n519), .A2(new_n258), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n214), .A2(G101), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT77), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n214), .A2(new_n215), .A3(G101), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n203), .A2(new_n478), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT10), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT10), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n477), .A2(KEYINPUT78), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n243), .A2(G128), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n232), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT78), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n238), .A2(new_n530), .A3(new_n476), .A4(G128), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n527), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n218), .A2(new_n526), .A3(new_n203), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n525), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n204), .A2(new_n240), .A3(new_n209), .ZN(new_n535));
  INV_X1    g349(.A(new_n464), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT79), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n534), .A2(new_n535), .A3(KEYINPUT79), .A4(new_n536), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n478), .B1(new_n218), .B2(new_n203), .ZN(new_n542));
  AND4_X1   g356(.A1(new_n203), .A2(new_n522), .A3(new_n523), .A4(new_n532), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n464), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT12), .ZN(new_n545));
  OR2_X1    g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n544), .A2(new_n545), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n541), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n287), .A2(G227), .ZN(new_n550));
  XNOR2_X1  g364(.A(G110), .B(G140), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n550), .B(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n553), .B1(new_n539), .B2(new_n540), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n534), .A2(new_n535), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n464), .ZN(new_n556));
  AOI22_X1  g370(.A1(new_n549), .A2(new_n553), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n520), .B1(new_n557), .B2(G469), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n541), .A2(new_n552), .A3(new_n548), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n552), .B1(new_n541), .B2(new_n556), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n519), .B(new_n258), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n518), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n402), .A2(new_n516), .A3(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(G101), .ZN(G3));
  INV_X1    g378(.A(KEYINPUT31), .ZN(new_n565));
  INV_X1    g379(.A(new_n496), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n483), .A2(new_n207), .ZN(new_n567));
  AOI21_X1  g381(.A(KEYINPUT65), .B1(new_n480), .B2(new_n456), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n469), .B1(new_n475), .B2(new_n477), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n463), .A2(new_n462), .B1(new_n237), .B2(new_n239), .ZN(new_n570));
  NOR4_X1   g384(.A1(new_n569), .A2(new_n570), .A3(new_n471), .A4(new_n207), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n567), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n566), .B1(new_n572), .B2(KEYINPUT28), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n565), .B1(new_n573), .B2(new_n491), .ZN(new_n574));
  INV_X1    g388(.A(new_n502), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n493), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(G472), .B1(new_n576), .B2(G902), .ZN(new_n577));
  OR2_X1    g391(.A1(new_n577), .A2(KEYINPUT92), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n503), .A2(new_n504), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(KEYINPUT92), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n453), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n582), .A2(new_n583), .A3(new_n562), .ZN(new_n584));
  INV_X1    g398(.A(new_n398), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n385), .B(new_n258), .C1(new_n382), .C2(new_n383), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n385), .A2(new_n258), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(KEYINPUT33), .B1(new_n375), .B2(KEYINPUT93), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n383), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n590), .B1(new_n591), .B2(new_n381), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n382), .A2(new_n383), .A3(new_n589), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n586), .B(new_n588), .C1(new_n594), .C2(new_n385), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n350), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n187), .B1(new_n272), .B2(new_n273), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n597), .A2(new_n270), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n598), .A2(new_n400), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n584), .A2(new_n585), .A3(new_n596), .A4(new_n599), .ZN(new_n600));
  XOR2_X1   g414(.A(KEYINPUT34), .B(G104), .Z(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(G6));
  INV_X1    g416(.A(new_n346), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n344), .A2(new_n279), .A3(new_n258), .A4(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n332), .B1(new_n347), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n387), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AND4_X1   g422(.A1(new_n585), .A2(new_n584), .A3(new_n599), .A4(new_n608), .ZN(new_n609));
  XOR2_X1   g423(.A(KEYINPUT35), .B(G107), .Z(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(KEYINPUT94), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n609), .B(new_n611), .ZN(G9));
  AND2_X1   g426(.A1(new_n444), .A2(KEYINPUT36), .ZN(new_n613));
  OR2_X1    g427(.A1(new_n446), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n443), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n614), .A2(new_n451), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n449), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n402), .A2(new_n562), .A3(new_n582), .A4(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(new_n618), .B(KEYINPUT37), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G110), .ZN(G12));
  INV_X1    g434(.A(G900), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n393), .B1(new_n396), .B2(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT95), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n605), .A2(new_n387), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(KEYINPUT96), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT96), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n605), .A2(new_n627), .A3(new_n387), .A4(new_n624), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n399), .B(new_n617), .C1(new_n597), .C2(new_n270), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n504), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n576), .A2(KEYINPUT32), .A3(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n515), .B1(new_n634), .B2(new_n505), .ZN(new_n635));
  INV_X1    g449(.A(new_n520), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n554), .A2(new_n556), .ZN(new_n637));
  AOI22_X1  g451(.A1(new_n539), .A2(new_n540), .B1(new_n546), .B2(new_n547), .ZN(new_n638));
  OAI211_X1 g452(.A(new_n637), .B(G469), .C1(new_n552), .C2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n561), .A2(new_n636), .A3(new_n639), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n635), .A2(new_n517), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n630), .A2(new_n632), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G128), .ZN(G30));
  INV_X1    g457(.A(KEYINPUT38), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT97), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n278), .A2(new_n645), .A3(new_n271), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n645), .B1(new_n278), .B2(new_n271), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n644), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n648), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n650), .A2(KEYINPUT38), .A3(new_n646), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n512), .A2(new_n500), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(G902), .B1(new_n498), .B2(new_n500), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI22_X1  g471(.A1(new_n506), .A2(new_n507), .B1(G472), .B2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(new_n617), .ZN(new_n659));
  XOR2_X1   g473(.A(new_n623), .B(KEYINPUT39), .Z(new_n660));
  NAND2_X1  g474(.A1(new_n562), .A2(new_n660), .ZN(new_n661));
  OR2_X1    g475(.A1(new_n661), .A2(KEYINPUT40), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n351), .A2(new_n399), .A3(new_n387), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n663), .B1(new_n661), .B2(KEYINPUT40), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n653), .A2(new_n659), .A3(new_n662), .A4(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G143), .ZN(G45));
  NOR3_X1   g480(.A1(new_n350), .A2(new_n595), .A3(new_n623), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n632), .A2(KEYINPUT98), .A3(new_n641), .A4(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT98), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n667), .A2(new_n562), .A3(new_n635), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n669), .B1(new_n670), .B2(new_n631), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G146), .ZN(G48));
  NAND2_X1  g487(.A1(new_n583), .A2(new_n635), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n559), .A2(new_n560), .ZN(new_n675));
  OAI21_X1  g489(.A(G469), .B1(new_n675), .B2(G902), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n676), .A2(new_n517), .A3(new_n561), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n678), .A2(new_n599), .A3(new_n585), .A4(new_n596), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT41), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G113), .ZN(G15));
  NAND4_X1  g495(.A1(new_n678), .A2(new_n599), .A3(new_n585), .A4(new_n608), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G116), .ZN(G18));
  NOR2_X1   g497(.A1(new_n631), .A2(new_n677), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n684), .A2(new_n635), .A3(new_n585), .A4(new_n388), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G119), .ZN(G21));
  NOR2_X1   g500(.A1(new_n663), .A2(new_n598), .ZN(new_n687));
  OR3_X1    g501(.A1(new_n501), .A2(KEYINPUT99), .A3(new_n502), .ZN(new_n688));
  OAI21_X1  g502(.A(KEYINPUT99), .B1(new_n501), .B2(new_n502), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n688), .A2(new_n494), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n577), .B1(new_n690), .B2(new_n633), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n691), .A2(new_n453), .ZN(new_n692));
  INV_X1    g506(.A(new_n677), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n687), .A2(new_n692), .A3(new_n585), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G122), .ZN(G24));
  INV_X1    g509(.A(new_n667), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n696), .A2(new_n691), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n684), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G125), .ZN(G27));
  AND3_X1   g513(.A1(new_n558), .A2(KEYINPUT100), .A3(new_n561), .ZN(new_n700));
  AOI21_X1  g514(.A(KEYINPUT100), .B1(new_n558), .B2(new_n561), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n517), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(KEYINPUT101), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT100), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n640), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n558), .A2(KEYINPUT100), .A3(new_n561), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n518), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT101), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n703), .A2(new_n709), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n597), .A2(new_n270), .A3(KEYINPUT81), .ZN(new_n711));
  INV_X1    g525(.A(new_n271), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n516), .B(new_n399), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n710), .A2(new_n667), .A3(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT42), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n710), .A2(KEYINPUT42), .A3(new_n714), .A4(new_n667), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G131), .ZN(G33));
  NAND3_X1  g534(.A1(new_n710), .A2(new_n630), .A3(new_n714), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G134), .ZN(G36));
  INV_X1    g536(.A(KEYINPUT46), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n637), .B1(new_n552), .B2(new_n638), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT45), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n557), .A2(KEYINPUT45), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n726), .A2(new_n727), .A3(G469), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n723), .B1(new_n729), .B2(new_n520), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n728), .A2(KEYINPUT46), .A3(new_n636), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n730), .A2(new_n561), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n517), .ZN(new_n733));
  INV_X1    g547(.A(new_n660), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n400), .B1(new_n278), .B2(new_n271), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n738));
  OAI21_X1  g552(.A(G478), .B1(new_n592), .B2(new_n593), .ZN(new_n739));
  AND3_X1   g553(.A1(new_n739), .A2(new_n586), .A3(new_n588), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n350), .A2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT43), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n350), .A2(new_n740), .A3(KEYINPUT43), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(new_n581), .A3(new_n617), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n737), .B1(new_n738), .B2(new_n746), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n735), .B(new_n747), .C1(new_n738), .C2(new_n746), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(KEYINPUT102), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G137), .ZN(G39));
  NOR2_X1   g564(.A1(new_n696), .A2(new_n635), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n736), .A2(new_n751), .A3(new_n453), .ZN(new_n752));
  XOR2_X1   g566(.A(new_n752), .B(KEYINPUT103), .Z(new_n753));
  INV_X1    g567(.A(KEYINPUT47), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n733), .B(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G140), .ZN(G42));
  AOI21_X1  g571(.A(new_n392), .B1(new_n743), .B2(new_n744), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n736), .A2(new_n758), .A3(new_n617), .A4(new_n693), .ZN(new_n759));
  OR3_X1    g573(.A1(new_n759), .A2(KEYINPUT110), .A3(new_n691), .ZN(new_n760));
  OAI21_X1  g574(.A(KEYINPUT110), .B1(new_n759), .B2(new_n691), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n736), .A2(new_n693), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n658), .A2(new_n393), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n762), .A2(new_n453), .A3(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n351), .A2(new_n740), .ZN(new_n765));
  AOI22_X1  g579(.A1(new_n760), .A2(new_n761), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n758), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n692), .A2(new_n693), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n767), .A2(new_n768), .A3(new_n399), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n652), .A2(KEYINPUT50), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT50), .B1(new_n652), .B2(new_n769), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n766), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n737), .A2(new_n767), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n676), .A2(new_n561), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT104), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT109), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n776), .A2(new_n777), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n778), .A2(new_n779), .A3(new_n517), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n692), .B(new_n774), .C1(new_n755), .C2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n773), .A2(KEYINPUT51), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n764), .A2(new_n596), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n774), .A2(new_n678), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(KEYINPUT48), .ZN(new_n785));
  AND4_X1   g599(.A1(new_n390), .A2(new_n782), .A3(new_n783), .A4(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT111), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n772), .A2(new_n787), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n766), .B(KEYINPUT111), .C1(new_n771), .C2(new_n770), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(new_n781), .A3(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT112), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT51), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n791), .B1(new_n790), .B2(new_n792), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n786), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n736), .A2(new_n617), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n705), .A2(new_n706), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n708), .B1(new_n797), .B2(new_n517), .ZN(new_n798));
  AOI211_X1 g612(.A(KEYINPUT101), .B(new_n518), .C1(new_n705), .C2(new_n706), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n697), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n606), .A2(new_n387), .A3(new_n623), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n641), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n796), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  AOI211_X1 g617(.A(new_n629), .B(new_n713), .C1(new_n703), .C2(new_n709), .ZN(new_n804));
  OAI21_X1  g618(.A(KEYINPUT106), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT106), .ZN(new_n806));
  INV_X1    g620(.A(new_n802), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n807), .B1(new_n710), .B2(new_n697), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n806), .B(new_n721), .C1(new_n808), .C2(new_n796), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n805), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n707), .A2(new_n687), .A3(new_n624), .A4(new_n659), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n672), .A2(new_n642), .A3(new_n698), .A4(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT52), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n641), .A2(new_n628), .A3(new_n626), .ZN(new_n815));
  AOI22_X1  g629(.A1(new_n815), .A2(new_n632), .B1(new_n684), .B2(new_n697), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n816), .A2(KEYINPUT52), .A3(new_n672), .A4(new_n811), .ZN(new_n817));
  AOI22_X1  g631(.A1(new_n814), .A2(new_n817), .B1(new_n717), .B2(new_n718), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n351), .A2(new_n607), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n278), .A2(new_n819), .A3(new_n271), .A4(new_n401), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT105), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n822), .A2(new_n584), .A3(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n711), .A2(new_n712), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n584), .A2(new_n825), .A3(new_n401), .A4(new_n596), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n824), .A2(new_n826), .A3(new_n563), .A4(new_n618), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n685), .A2(new_n679), .A3(new_n682), .A4(new_n694), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n810), .A2(new_n818), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n810), .A2(new_n818), .A3(KEYINPUT53), .A4(new_n829), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n832), .A2(KEYINPUT107), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT107), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n830), .A2(new_n835), .A3(new_n831), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n834), .A2(KEYINPUT54), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT108), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n828), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(KEYINPUT53), .B1(new_n828), .B2(new_n839), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n827), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n842), .A2(new_n810), .A3(new_n818), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n832), .A2(new_n838), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n837), .A2(new_n844), .ZN(new_n845));
  NOR4_X1   g659(.A1(new_n767), .A2(new_n768), .A3(new_n598), .A4(new_n400), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n795), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n389), .A2(new_n250), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(KEYINPUT113), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n776), .B(KEYINPUT49), .ZN(new_n850));
  NOR4_X1   g664(.A1(new_n653), .A2(new_n453), .A3(new_n850), .A4(new_n518), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n851), .A2(new_n399), .A3(new_n658), .ZN(new_n852));
  OAI22_X1  g666(.A1(new_n847), .A2(new_n849), .B1(new_n741), .B2(new_n852), .ZN(G75));
  AOI21_X1  g667(.A(new_n258), .B1(new_n832), .B2(new_n843), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT56), .B1(new_n854), .B2(G210), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n262), .A2(new_n265), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(new_n263), .ZN(new_n857));
  XOR2_X1   g671(.A(new_n857), .B(KEYINPUT55), .Z(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  OR3_X1    g673(.A1(new_n855), .A2(KEYINPUT114), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n287), .A2(G952), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n861), .B1(new_n855), .B2(KEYINPUT114), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n859), .B1(new_n855), .B2(KEYINPUT114), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n860), .A2(new_n862), .A3(new_n863), .ZN(G51));
  INV_X1    g678(.A(KEYINPUT115), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n854), .A2(new_n729), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n520), .B(KEYINPUT57), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n832), .A2(new_n838), .A3(new_n843), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n838), .B1(new_n832), .B2(new_n843), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(new_n675), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n866), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n865), .B1(new_n872), .B2(new_n861), .ZN(new_n873));
  INV_X1    g687(.A(new_n861), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n832), .A2(new_n843), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT54), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n844), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n675), .B1(new_n877), .B2(new_n867), .ZN(new_n878));
  OAI211_X1 g692(.A(KEYINPUT115), .B(new_n874), .C1(new_n878), .C2(new_n866), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n873), .A2(new_n879), .ZN(G54));
  NAND3_X1  g694(.A1(new_n854), .A2(KEYINPUT58), .A3(G475), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT117), .ZN(new_n882));
  INV_X1    g696(.A(new_n344), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n882), .B1(new_n881), .B2(new_n883), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n874), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n854), .A2(KEYINPUT58), .A3(G475), .A4(new_n344), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT116), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n886), .A2(new_n888), .ZN(G60));
  XNOR2_X1  g703(.A(new_n587), .B(KEYINPUT59), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n877), .A2(new_n594), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n890), .B1(new_n837), .B2(new_n844), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n892), .B(new_n874), .C1(new_n893), .C2(new_n594), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(G63));
  NAND2_X1  g709(.A1(G217), .A2(G902), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT60), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n897), .B1(new_n832), .B2(new_n843), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n898), .A2(new_n446), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n899), .A2(new_n861), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n614), .A2(new_n615), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n898), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n900), .A2(KEYINPUT61), .A3(new_n903), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n898), .A2(KEYINPUT119), .A3(new_n902), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT119), .B1(new_n898), .B2(new_n902), .ZN(new_n906));
  NOR4_X1   g720(.A1(new_n905), .A2(new_n906), .A3(new_n899), .A4(new_n861), .ZN(new_n907));
  XNOR2_X1  g721(.A(KEYINPUT118), .B(KEYINPUT61), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n904), .B1(new_n907), .B2(new_n908), .ZN(G66));
  INV_X1    g723(.A(G224), .ZN(new_n910));
  OAI21_X1  g724(.A(G953), .B1(new_n397), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n911), .B1(new_n829), .B2(new_n394), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n856), .B1(G898), .B2(new_n287), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT120), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n912), .B(new_n914), .ZN(G69));
  AND2_X1   g729(.A1(new_n756), .A2(new_n748), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n735), .A2(new_n516), .A3(new_n687), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT123), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n816), .A2(new_n672), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n719), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n916), .A2(new_n918), .A3(new_n721), .A4(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(new_n287), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n484), .A2(new_n486), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(new_n335), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n287), .A2(G900), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT122), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n922), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n287), .B1(G227), .B2(G900), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n665), .A2(new_n919), .ZN(new_n929));
  XOR2_X1   g743(.A(KEYINPUT121), .B(KEYINPUT62), .Z(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT62), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n665), .B(new_n919), .C1(KEYINPUT121), .C2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n819), .A2(new_n596), .ZN(new_n934));
  OR3_X1    g748(.A1(new_n713), .A2(new_n661), .A3(new_n934), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n931), .A2(new_n916), .A3(new_n933), .A4(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n287), .ZN(new_n937));
  OAI221_X1 g751(.A(new_n927), .B1(KEYINPUT124), .B2(new_n928), .C1(new_n924), .C2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n928), .A2(KEYINPUT124), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(G72));
  NAND2_X1  g754(.A1(G472), .A2(G902), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT63), .Z(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT125), .Z(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n829), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n944), .B1(new_n936), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(KEYINPUT126), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT126), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n948), .B(new_n944), .C1(new_n936), .C2(new_n945), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n947), .A2(new_n654), .A3(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n944), .B1(new_n921), .B2(new_n945), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT127), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n512), .A2(new_n500), .ZN(new_n954));
  OAI211_X1 g768(.A(KEYINPUT127), .B(new_n944), .C1(new_n921), .C2(new_n945), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n950), .A2(new_n956), .A3(new_n874), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n834), .A2(new_n836), .A3(new_n942), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n958), .A2(new_n654), .A3(new_n954), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n957), .A2(new_n959), .ZN(G57));
endmodule


