//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 0 0 0 0 0 1 0 0 0 1 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 1 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n438, new_n445, new_n446, new_n447, new_n452,
    new_n456, new_n457, new_n458, new_n459, new_n460, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n564,
    new_n566, new_n567, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n614, new_n617, new_n619,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1175, new_n1176, new_n1177, new_n1178;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  OR2_X1    g011(.A1(new_n436), .A2(KEYINPUT65), .ZN(new_n437));
  NAND2_X1  g012(.A1(new_n436), .A2(KEYINPUT65), .ZN(new_n438));
  NAND2_X1  g013(.A1(new_n437), .A2(new_n438), .ZN(G220));
  XNOR2_X1  g014(.A(KEYINPUT66), .B(G96), .ZN(G221));
  INV_X1    g015(.A(G69), .ZN(G235));
  INV_X1    g016(.A(G120), .ZN(G236));
  INV_X1    g017(.A(G57), .ZN(G237));
  INV_X1    g018(.A(G108), .ZN(G238));
  INV_X1    g019(.A(G2072), .ZN(new_n445));
  INV_X1    g020(.A(G2078), .ZN(new_n446));
  NOR2_X1   g021(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g022(.A1(new_n447), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g023(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g024(.A(G452), .Z(G391));
  AND2_X1   g025(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g026(.A1(G7), .A2(G661), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g028(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g029(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR3_X1   g030(.A1(G221), .A2(G218), .A3(G219), .ZN(new_n456));
  NAND3_X1  g031(.A1(new_n437), .A2(new_n456), .A3(new_n438), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT2), .ZN(new_n458));
  NOR4_X1   g033(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n458), .A2(new_n460), .ZN(G325));
  INV_X1    g036(.A(G325), .ZN(G261));
  NAND2_X1  g037(.A1(new_n458), .A2(G2106), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(KEYINPUT67), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n464), .B1(G567), .B2(new_n460), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(KEYINPUT67), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(G319));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  AND2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(G137), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT68), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n471), .B1(new_n474), .B2(new_n479), .ZN(new_n480));
  XNOR2_X1  g055(.A(KEYINPUT68), .B(G2105), .ZN(new_n481));
  OAI21_X1  g056(.A(G125), .B1(new_n472), .B2(new_n473), .ZN(new_n482));
  NAND2_X1  g057(.A1(G113), .A2(G2104), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n480), .A2(new_n484), .ZN(G160));
  OAI221_X1 g060(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n481), .C2(G112), .ZN(new_n486));
  INV_X1    g061(.A(G124), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT3), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(new_n469), .ZN(new_n489));
  NAND2_X1  g064(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(new_n479), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n486), .B1(new_n487), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n472), .A2(new_n473), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT69), .B1(new_n494), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n491), .A2(new_n496), .A3(new_n475), .ZN(new_n497));
  AND2_X1   g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n493), .B1(G136), .B2(new_n498), .ZN(G162));
  NOR2_X1   g074(.A1(new_n475), .A2(G114), .ZN(new_n500));
  OAI21_X1  g075(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT70), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OR2_X1    g077(.A1(G102), .A2(G2105), .ZN(new_n503));
  INV_X1    g078(.A(G114), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G2105), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n503), .A2(new_n505), .A3(new_n506), .A4(G2104), .ZN(new_n507));
  AND2_X1   g082(.A1(G126), .A2(G2105), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n502), .A2(new_n507), .B1(new_n491), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g084(.A(G138), .B1(new_n472), .B2(new_n473), .ZN(new_n510));
  NOR3_X1   g085(.A1(new_n510), .A2(new_n479), .A3(KEYINPUT4), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT4), .ZN(new_n512));
  INV_X1    g087(.A(G138), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n513), .B1(new_n489), .B2(new_n490), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n512), .B1(new_n514), .B2(new_n481), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n509), .B1(new_n511), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(G164));
  OR2_X1    g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT5), .B(G543), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G543), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n523), .B1(new_n518), .B2(new_n519), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n522), .A2(G88), .B1(G50), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT71), .ZN(new_n526));
  INV_X1    g101(.A(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n521), .A2(G62), .ZN(new_n528));
  NAND2_X1  g103(.A1(G75), .A2(G543), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n525), .B1(new_n526), .B2(new_n530), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n530), .A2(new_n526), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(G166));
  XOR2_X1   g108(.A(KEYINPUT72), .B(KEYINPUT7), .Z(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n534), .B(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n524), .A2(G51), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n520), .A2(new_n521), .ZN(new_n540));
  INV_X1    g115(.A(G89), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n538), .A2(new_n542), .ZN(G286));
  INV_X1    g118(.A(G286), .ZN(G168));
  NAND2_X1  g119(.A1(new_n524), .A2(G52), .ZN(new_n545));
  INV_X1    g120(.A(G90), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n540), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(new_n527), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n547), .A2(new_n549), .ZN(G171));
  AND3_X1   g125(.A1(new_n520), .A2(new_n521), .A3(G81), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT73), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n524), .A2(G43), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n554), .ZN(new_n556));
  OAI21_X1  g131(.A(KEYINPUT73), .B1(new_n556), .B2(new_n551), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n559), .A2(new_n527), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n564));
  XOR2_X1   g139(.A(new_n564), .B(KEYINPUT74), .Z(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  NAND3_X1  g143(.A1(new_n522), .A2(KEYINPUT75), .A3(G91), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n570));
  INV_X1    g145(.A(G91), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n540), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(new_n521), .ZN(new_n574));
  XNOR2_X1  g149(.A(KEYINPUT76), .B(G65), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n569), .A2(new_n572), .B1(G651), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n524), .A2(G53), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT9), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n577), .A2(new_n579), .ZN(G299));
  INV_X1    g155(.A(G171), .ZN(G301));
  INV_X1    g156(.A(G166), .ZN(G303));
  NAND2_X1  g157(.A1(new_n524), .A2(G49), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n520), .A2(new_n521), .A3(G87), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(G288));
  NAND2_X1  g161(.A1(new_n524), .A2(G48), .ZN(new_n587));
  INV_X1    g162(.A(G86), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n540), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n521), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n590), .A2(new_n527), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G305));
  NAND2_X1  g168(.A1(new_n524), .A2(G47), .ZN(new_n594));
  INV_X1    g169(.A(G85), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n540), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n597), .A2(new_n527), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  AND3_X1   g176(.A1(new_n520), .A2(new_n521), .A3(G92), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT10), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  XOR2_X1   g179(.A(KEYINPUT77), .B(G66), .Z(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n574), .B2(new_n605), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n606), .A2(G651), .B1(G54), .B2(new_n524), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n601), .B1(new_n609), .B2(G868), .ZN(G284));
  OAI21_X1  g185(.A(new_n601), .B1(new_n609), .B2(G868), .ZN(G321));
  NAND2_X1  g186(.A1(G286), .A2(G868), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT78), .Z(new_n613));
  INV_X1    g188(.A(G299), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(G868), .B2(new_n614), .ZN(G297));
  OAI21_X1  g190(.A(new_n613), .B1(G868), .B2(new_n614), .ZN(G280));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n609), .B1(new_n617), .B2(G860), .ZN(G148));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n561), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n608), .A2(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(new_n619), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n491), .A2(new_n470), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT12), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2100), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n494), .A2(new_n481), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G123), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT79), .Z(new_n630));
  NAND2_X1  g205(.A1(new_n498), .A2(G135), .ZN(new_n631));
  OAI221_X1 g206(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n481), .C2(G111), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n633), .A2(G2096), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(G2096), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n627), .A2(new_n634), .A3(new_n635), .ZN(G156));
  INV_X1    g211(.A(G14), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2427), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(KEYINPUT14), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n637), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  INV_X1    g226(.A(KEYINPUT80), .ZN(new_n652));
  AND2_X1   g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n650), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(G401));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  XNOR2_X1  g232(.A(G2072), .B(G2078), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT18), .Z(new_n661));
  AOI21_X1  g236(.A(new_n659), .B1(new_n658), .B2(KEYINPUT81), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n662), .B1(KEYINPUT81), .B2(new_n658), .ZN(new_n663));
  INV_X1    g238(.A(new_n657), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n658), .B(KEYINPUT17), .Z(new_n665));
  INV_X1    g240(.A(new_n659), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n663), .B(new_n664), .C1(new_n665), .C2(new_n666), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n665), .A2(new_n666), .A3(new_n657), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n661), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G2096), .B(G2100), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(G227));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1956), .B(G2474), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1961), .B(G1966), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n675), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n673), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n680), .A2(KEYINPUT83), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n679), .B(new_n681), .Z(new_n682));
  NAND2_X1  g257(.A1(new_n680), .A2(new_n676), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n684));
  XOR2_X1   g259(.A(new_n683), .B(new_n684), .Z(new_n685));
  NOR2_X1   g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  AND2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  XOR2_X1   g264(.A(G1991), .B(G1996), .Z(new_n690));
  OR3_X1    g265(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n690), .B1(new_n688), .B2(new_n689), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n693), .B(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(G229));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT30), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n698), .B1(new_n699), .B2(G28), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT97), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n699), .A2(G28), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(new_n701), .B2(new_n702), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT31), .B(G11), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n707), .A2(G21), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G286), .B2(G16), .ZN(new_n709));
  INV_X1    g284(.A(G1966), .ZN(new_n710));
  OAI22_X1  g285(.A1(new_n709), .A2(new_n710), .B1(new_n633), .B2(new_n698), .ZN(new_n711));
  AOI211_X1 g286(.A(new_n706), .B(new_n711), .C1(new_n710), .C2(new_n709), .ZN(new_n712));
  NOR2_X1   g287(.A1(G4), .A2(G16), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT91), .Z(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(new_n608), .B2(new_n707), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT92), .B(G1348), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n698), .A2(G26), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT28), .Z(new_n719));
  NAND2_X1  g294(.A1(new_n498), .A2(G140), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n628), .A2(G128), .ZN(new_n721));
  OAI221_X1 g296(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n481), .C2(G116), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n719), .B1(new_n724), .B2(G29), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G2067), .ZN(new_n726));
  NOR2_X1   g301(.A1(G16), .A2(G19), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n562), .B2(G16), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G1341), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n712), .A2(new_n717), .A3(new_n726), .A4(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n698), .A2(G35), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G162), .B2(new_n698), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT29), .Z(new_n733));
  INV_X1    g308(.A(G2090), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT100), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n698), .A2(G27), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G164), .B2(new_n698), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(new_n446), .ZN(new_n738));
  OAI22_X1  g313(.A1(new_n733), .A2(new_n734), .B1(new_n735), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n730), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n733), .A2(new_n734), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n738), .A2(new_n735), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n707), .A2(G20), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT23), .Z(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G299), .B2(G16), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G1956), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n740), .A2(new_n741), .A3(new_n742), .A4(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(G5), .A2(G16), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT98), .Z(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G301), .B2(new_n707), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT99), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G1961), .ZN(new_n752));
  NAND2_X1  g327(.A1(G160), .A2(G29), .ZN(new_n753));
  AND2_X1   g328(.A1(KEYINPUT24), .A2(G34), .ZN(new_n754));
  NOR2_X1   g329(.A1(KEYINPUT24), .A2(G34), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n698), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT94), .Z(new_n757));
  NAND2_X1  g332(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT95), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(G2084), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n698), .A2(G33), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n491), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n762), .A2(new_n481), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT93), .Z(new_n764));
  NAND2_X1  g339(.A1(new_n498), .A2(G139), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n481), .A2(G103), .A3(G2104), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT25), .Z(new_n767));
  NAND3_X1  g342(.A1(new_n764), .A2(new_n765), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n761), .B1(new_n768), .B2(G29), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(new_n445), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n760), .A2(new_n770), .ZN(new_n771));
  OAI22_X1  g346(.A1(new_n769), .A2(new_n445), .B1(new_n728), .B2(G1341), .ZN(new_n772));
  NOR3_X1   g347(.A1(new_n752), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n698), .A2(G32), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n470), .A2(G105), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT96), .ZN(new_n776));
  NAND3_X1  g351(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT26), .Z(new_n778));
  NAND2_X1  g353(.A1(new_n628), .A2(G129), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n776), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n498), .B2(G141), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n774), .B1(new_n781), .B2(new_n698), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT27), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1996), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n773), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n747), .A2(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT36), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n707), .A2(G22), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G166), .B2(new_n707), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT90), .Z(new_n791));
  OR2_X1    g366(.A1(new_n791), .A2(G1971), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(G1971), .ZN(new_n793));
  MUX2_X1   g368(.A(G23), .B(G288), .S(G16), .Z(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT33), .B(G1976), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT89), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n794), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n707), .A2(G6), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(new_n592), .B2(new_n707), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT87), .B(KEYINPUT88), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT32), .B(G1981), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n801), .A2(new_n803), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n797), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n792), .A2(new_n793), .A3(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n807), .A2(KEYINPUT34), .ZN(new_n808));
  NOR2_X1   g383(.A1(G16), .A2(G24), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n599), .B(KEYINPUT85), .Z(new_n810));
  AOI21_X1  g385(.A(new_n809), .B1(new_n810), .B2(G16), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(G1986), .Z(new_n812));
  INV_X1    g387(.A(KEYINPUT86), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n812), .A2(new_n813), .ZN(new_n815));
  NOR2_X1   g390(.A1(G25), .A2(G29), .ZN(new_n816));
  OAI221_X1 g391(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n481), .C2(G107), .ZN(new_n817));
  INV_X1    g392(.A(G119), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(new_n492), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(G131), .B2(new_n498), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n816), .B1(new_n820), .B2(G29), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT84), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT35), .B(G1991), .Z(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n815), .A2(new_n824), .ZN(new_n825));
  NOR3_X1   g400(.A1(new_n808), .A2(new_n814), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n807), .A2(KEYINPUT34), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n788), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n826), .A2(new_n788), .A3(new_n827), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n787), .B1(new_n829), .B2(new_n830), .ZN(G311));
  INV_X1    g406(.A(new_n830), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n786), .B1(new_n832), .B2(new_n828), .ZN(G150));
  NAND2_X1  g408(.A1(new_n609), .A2(G559), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT102), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT38), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n524), .A2(G55), .ZN(new_n837));
  INV_X1    g412(.A(G93), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n837), .B1(new_n838), .B2(new_n540), .ZN(new_n839));
  AOI22_X1  g414(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n840), .A2(new_n527), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT101), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n839), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OR3_X1    g418(.A1(new_n840), .A2(new_n842), .A3(new_n527), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n561), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n558), .A2(new_n843), .A3(new_n560), .A4(new_n844), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n836), .B(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT39), .ZN(new_n850));
  AOI21_X1  g425(.A(G860), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(new_n850), .B2(new_n849), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n845), .A2(G860), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT37), .Z(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n854), .ZN(G145));
  XNOR2_X1  g430(.A(G162), .B(G160), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT103), .Z(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n633), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n724), .B(new_n516), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n768), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n860), .A2(new_n781), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n781), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n498), .A2(G142), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n628), .A2(G130), .ZN(new_n865));
  OAI221_X1 g440(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n481), .C2(G118), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n625), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(new_n820), .Z(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(KEYINPUT105), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n858), .B1(new_n863), .B2(new_n870), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n863), .A2(new_n870), .ZN(new_n872));
  AOI21_X1  g447(.A(G37), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT104), .ZN(new_n874));
  INV_X1    g449(.A(new_n869), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n863), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n861), .B(new_n862), .C1(KEYINPUT104), .C2(new_n869), .ZN(new_n877));
  OAI211_X1 g452(.A(new_n876), .B(new_n877), .C1(new_n874), .C2(new_n875), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(new_n858), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n873), .A2(new_n879), .A3(KEYINPUT40), .ZN(new_n880));
  AOI21_X1  g455(.A(KEYINPUT40), .B1(new_n873), .B2(new_n879), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(G395));
  OR2_X1    g457(.A1(new_n592), .A2(KEYINPUT107), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n592), .A2(KEYINPUT107), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n885), .A2(G166), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n599), .B(G288), .Z(new_n888));
  NAND2_X1  g463(.A1(new_n885), .A2(G166), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n888), .B1(new_n887), .B2(new_n889), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT42), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(KEYINPUT108), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n893), .A2(KEYINPUT108), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n895), .B(new_n896), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n848), .B(KEYINPUT106), .Z(new_n898));
  AND2_X1   g473(.A1(new_n898), .A2(new_n621), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(new_n621), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n614), .A2(new_n609), .ZN(new_n901));
  NAND2_X1  g476(.A1(G299), .A2(new_n608), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  OR3_X1    g479(.A1(new_n899), .A2(new_n900), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT41), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n901), .A2(new_n906), .A3(new_n902), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n903), .A2(KEYINPUT41), .ZN(new_n908));
  OAI211_X1 g483(.A(new_n907), .B(new_n908), .C1(new_n899), .C2(new_n900), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n897), .A2(new_n905), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n897), .B1(new_n905), .B2(new_n909), .ZN(new_n911));
  OAI21_X1  g486(.A(G868), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n845), .A2(new_n619), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(G295));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n913), .ZN(G331));
  OR2_X1    g490(.A1(new_n890), .A2(new_n891), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n846), .A2(G301), .A3(new_n847), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(G301), .B1(new_n846), .B2(new_n847), .ZN(new_n919));
  OAI21_X1  g494(.A(G286), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n919), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n921), .A2(G168), .A3(new_n917), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n908), .A2(new_n907), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n920), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n903), .B1(new_n920), .B2(new_n922), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n916), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(G37), .ZN(new_n927));
  AOI21_X1  g502(.A(G168), .B1(new_n921), .B2(new_n917), .ZN(new_n928));
  NOR3_X1   g503(.A1(new_n918), .A2(new_n919), .A3(G286), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n904), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n920), .A2(new_n922), .A3(new_n923), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(new_n892), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n926), .A2(new_n927), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n908), .A2(KEYINPUT109), .A3(new_n907), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n903), .A2(new_n936), .A3(KEYINPUT41), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n935), .A2(new_n920), .A3(new_n922), .A4(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n930), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n916), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n940), .A2(new_n941), .A3(new_n927), .A4(new_n932), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n934), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n943), .A2(KEYINPUT44), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n932), .A2(new_n927), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n892), .B1(new_n930), .B2(new_n938), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT111), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT111), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n940), .A2(new_n948), .A3(new_n927), .A4(new_n932), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n947), .A2(KEYINPUT43), .A3(new_n949), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n926), .A2(new_n932), .A3(new_n941), .A4(new_n927), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT110), .ZN(new_n952));
  OR2_X1    g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n952), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n950), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n944), .B1(new_n955), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g531(.A(G1384), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n516), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(G160), .A2(G40), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G2067), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n724), .B(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n963), .B1(new_n965), .B2(new_n781), .ZN(new_n966));
  OR3_X1    g541(.A1(new_n963), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT46), .B1(new_n963), .B2(G1996), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n969), .B(KEYINPUT47), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n781), .B(G1996), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n971), .A2(new_n823), .A3(new_n820), .A4(new_n965), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n720), .A2(new_n723), .A3(new_n964), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n963), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n974), .B(KEYINPUT126), .ZN(new_n975));
  XOR2_X1   g550(.A(new_n820), .B(new_n823), .Z(new_n976));
  AND3_X1   g551(.A1(new_n976), .A2(new_n965), .A3(new_n971), .ZN(new_n977));
  OR3_X1    g552(.A1(new_n963), .A2(G1986), .A3(G290), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT48), .ZN(new_n979));
  OAI22_X1  g554(.A1(new_n977), .A2(new_n963), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n980), .B1(new_n979), .B2(new_n978), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n970), .A2(new_n975), .A3(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT49), .ZN(new_n983));
  OAI21_X1  g558(.A(G1981), .B1(new_n589), .B2(new_n591), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n589), .A2(new_n591), .A3(G1981), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n983), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G1981), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n592), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n989), .A2(KEYINPUT49), .A3(new_n984), .ZN(new_n990));
  INV_X1    g565(.A(G8), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT4), .B1(new_n510), .B2(new_n479), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n491), .A2(new_n481), .A3(new_n512), .A4(G138), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(G1384), .B1(new_n994), .B2(new_n509), .ZN(new_n995));
  INV_X1    g570(.A(G40), .ZN(new_n996));
  NOR3_X1   g571(.A1(new_n480), .A2(new_n484), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n991), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n987), .A2(new_n990), .A3(new_n998), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n583), .A2(new_n584), .A3(new_n585), .A4(G1976), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n1000), .B(KEYINPUT114), .ZN(new_n1001));
  INV_X1    g576(.A(G1976), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT52), .B1(G288), .B2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n998), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n999), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1006), .B1(new_n998), .B2(new_n1001), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n997), .B1(new_n995), .B2(KEYINPUT45), .ZN(new_n1009));
  AOI211_X1 g584(.A(G1384), .B(new_n959), .C1(new_n994), .C2(new_n509), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n710), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n958), .A2(KEYINPUT50), .ZN(new_n1012));
  INV_X1    g587(.A(G2084), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT50), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n995), .A2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1012), .A2(new_n1013), .A3(new_n997), .A4(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n991), .B1(new_n1011), .B2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1008), .A2(G168), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1971), .ZN(new_n1019));
  INV_X1    g594(.A(new_n959), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n997), .B1(new_n995), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT45), .ZN(new_n1022));
  AOI211_X1 g597(.A(new_n1022), .B(G1384), .C1(new_n994), .C2(new_n509), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1019), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1012), .A2(new_n734), .A3(new_n997), .A4(new_n1015), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n991), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(G8), .B1(new_n531), .B2(new_n532), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n1027), .B(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT63), .B1(new_n1018), .B2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(G288), .A2(G1976), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n986), .B1(new_n999), .B2(new_n1032), .ZN(new_n1033));
  OR2_X1    g608(.A1(new_n1033), .A2(KEYINPUT115), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(KEYINPUT115), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1034), .A2(new_n998), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1031), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1008), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n997), .B1(new_n995), .B2(new_n1014), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n958), .A2(new_n1041), .A3(KEYINPUT50), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT116), .B1(new_n995), .B2(new_n1014), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1040), .B(new_n734), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n991), .B1(new_n1044), .B2(new_n1024), .ZN(new_n1045));
  OR2_X1    g620(.A1(new_n1045), .A2(new_n1029), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1017), .ZN(new_n1047));
  NOR3_X1   g622(.A1(new_n1047), .A2(KEYINPUT63), .A3(G286), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT113), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1026), .A2(new_n1029), .A3(KEYINPUT113), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1038), .B1(new_n1049), .B2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1037), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n1057));
  XNOR2_X1  g632(.A(G299), .B(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1059));
  XNOR2_X1  g634(.A(KEYINPUT56), .B(G2072), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1015), .A2(new_n1041), .ZN(new_n1062));
  AOI211_X1 g637(.A(KEYINPUT50), .B(G1384), .C1(new_n994), .C2(new_n509), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT116), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1039), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1058), .B(new_n1061), .C1(new_n1065), .C2(G1956), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n995), .A2(new_n1067), .A3(new_n997), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1067), .B1(new_n995), .B2(new_n997), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n964), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G1348), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(new_n1039), .B2(new_n1063), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n608), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1066), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1058), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1076));
  AOI21_X1  g651(.A(G1956), .B1(new_n1076), .B2(new_n1040), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1023), .ZN(new_n1078));
  AND4_X1   g653(.A1(new_n997), .A2(new_n1078), .A3(new_n960), .A4(new_n1060), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1075), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1074), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1040), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1083));
  INV_X1    g658(.A(G1956), .ZN(new_n1084));
  AOI22_X1  g659(.A1(new_n1083), .A2(new_n1084), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1082), .B1(new_n1085), .B2(new_n1058), .ZN(new_n1086));
  AOI22_X1  g661(.A1(new_n1086), .A2(KEYINPUT61), .B1(new_n1066), .B2(new_n1080), .ZN(new_n1087));
  AND4_X1   g662(.A1(KEYINPUT119), .A2(new_n1080), .A3(KEYINPUT61), .A4(new_n1066), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1070), .A2(new_n608), .A3(new_n1072), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT60), .B1(new_n1090), .B2(new_n1073), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n608), .A2(KEYINPUT60), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1070), .A2(new_n1072), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(G1996), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1059), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(KEYINPUT118), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT118), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1059), .A2(new_n1098), .A3(new_n1095), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT58), .B(G1341), .Z(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1097), .A2(new_n1099), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(new_n562), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT59), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT59), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1103), .A2(new_n1106), .A3(new_n562), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1094), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1081), .B1(new_n1089), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(G286), .A2(G8), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT120), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n961), .B1(new_n958), .B2(new_n1022), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1010), .ZN(new_n1113));
  AOI21_X1  g688(.A(G1966), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NOR3_X1   g689(.A1(new_n1039), .A2(G2084), .A3(new_n1063), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1111), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1011), .A2(new_n1016), .A3(KEYINPUT120), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1110), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1116), .A2(G168), .A3(new_n1117), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT51), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1120), .A2(new_n991), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1110), .ZN(new_n1123));
  NOR3_X1   g698(.A1(new_n1017), .A2(KEYINPUT51), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1118), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT123), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1026), .A2(KEYINPUT113), .A3(new_n1029), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT113), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1008), .B1(new_n1029), .B2(new_n1045), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1128), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1054), .A2(KEYINPUT123), .A3(new_n1046), .A4(new_n1008), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1059), .A2(new_n446), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT53), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1039), .A2(new_n1063), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1137), .B1(G1961), .B2(new_n1138), .ZN(new_n1139));
  XOR2_X1   g714(.A(G171), .B(KEYINPUT54), .Z(new_n1140));
  NOR2_X1   g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g716(.A(KEYINPUT121), .B(G2078), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1059), .A2(KEYINPUT53), .A3(new_n1142), .ZN(new_n1143));
  XOR2_X1   g718(.A(new_n1143), .B(KEYINPUT122), .Z(new_n1144));
  NAND4_X1  g719(.A1(new_n1112), .A2(KEYINPUT53), .A3(new_n1113), .A4(new_n446), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1137), .B(new_n1145), .C1(G1961), .C2(new_n1138), .ZN(new_n1146));
  AOI22_X1  g721(.A1(new_n1141), .A2(new_n1144), .B1(new_n1146), .B2(new_n1140), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1127), .A2(new_n1133), .A3(new_n1134), .A4(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1056), .B1(new_n1109), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT62), .ZN(new_n1150));
  OAI21_X1  g725(.A(KEYINPUT125), .B1(new_n1126), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT125), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1124), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1152), .B(KEYINPUT62), .C1(new_n1153), .C2(new_n1118), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1118), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1121), .ZN(new_n1157));
  AND3_X1   g732(.A1(new_n1011), .A2(new_n1016), .A3(KEYINPUT120), .ZN(new_n1158));
  AOI21_X1  g733(.A(KEYINPUT120), .B1(new_n1011), .B2(new_n1016), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1157), .B1(new_n1160), .B2(G168), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n1150), .B(new_n1156), .C1(new_n1161), .C2(new_n1124), .ZN(new_n1162));
  AND2_X1   g737(.A1(new_n1146), .A2(G171), .ZN(new_n1163));
  AND4_X1   g738(.A1(new_n1162), .A2(new_n1133), .A3(new_n1134), .A4(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1155), .B1(new_n1164), .B2(KEYINPUT124), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT124), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1133), .A2(new_n1134), .A3(new_n1163), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1162), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1166), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1149), .B1(new_n1165), .B2(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n599), .B(G1986), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n963), .B1(new_n977), .B2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n982), .B1(new_n1170), .B2(new_n1172), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g748(.A1(new_n467), .A2(G227), .ZN(new_n1175));
  XNOR2_X1  g749(.A(new_n1175), .B(KEYINPUT127), .ZN(new_n1176));
  AND3_X1   g750(.A1(new_n696), .A2(new_n655), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g751(.A1(new_n873), .A2(new_n879), .ZN(new_n1178));
  AND3_X1   g752(.A1(new_n1177), .A2(new_n1178), .A3(new_n943), .ZN(G308));
  NAND3_X1  g753(.A1(new_n1177), .A2(new_n1178), .A3(new_n943), .ZN(G225));
endmodule


