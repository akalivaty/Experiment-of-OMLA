//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 0 1 1 0 1 0 0 1 0 1 1 0 0 1 0 1 1 1 0 1 0 0 1 1 0 1 1 1 0 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028;
  INV_X1    g000(.A(KEYINPUT23), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G128), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(G128), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT23), .A3(G119), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n190), .A3(new_n192), .ZN(new_n193));
  OR2_X1    g007(.A1(new_n193), .A2(KEYINPUT75), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(KEYINPUT75), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(new_n195), .A3(G110), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT76), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n194), .A2(new_n195), .A3(KEYINPUT76), .A4(G110), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n191), .A2(G119), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(new_n190), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT24), .B(G110), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT77), .ZN(new_n205));
  INV_X1    g019(.A(G140), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G125), .ZN(new_n207));
  INV_X1    g021(.A(G125), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G140), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT16), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n205), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n207), .A2(new_n209), .A3(KEYINPUT77), .A4(KEYINPUT16), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n211), .A2(new_n206), .A3(G125), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n212), .A2(G146), .A3(new_n213), .A4(new_n214), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n204), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n200), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n202), .A2(new_n203), .ZN(new_n221));
  INV_X1    g035(.A(G110), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n189), .A2(new_n192), .A3(new_n222), .A4(new_n190), .ZN(new_n223));
  INV_X1    g037(.A(new_n210), .ZN(new_n224));
  AND2_X1   g038(.A1(KEYINPUT64), .A2(G146), .ZN(new_n225));
  NOR2_X1   g039(.A1(KEYINPUT64), .A2(G146), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n221), .A2(new_n223), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n218), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n220), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G953), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(G221), .A3(G234), .ZN(new_n232));
  XNOR2_X1  g046(.A(new_n232), .B(KEYINPUT22), .ZN(new_n233));
  XNOR2_X1  g047(.A(new_n233), .B(G137), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n230), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G902), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n220), .A2(new_n229), .A3(new_n234), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT25), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT25), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n236), .A2(new_n241), .A3(new_n237), .A4(new_n238), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT73), .B(G217), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n244), .B1(G234), .B2(new_n237), .ZN(new_n245));
  XOR2_X1   g059(.A(new_n245), .B(KEYINPUT74), .Z(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n240), .A2(new_n242), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n236), .A2(new_n238), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n245), .A2(G902), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(KEYINPUT78), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  OR3_X1    g066(.A1(new_n249), .A2(KEYINPUT78), .A3(new_n251), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n248), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  OR2_X1    g068(.A1(KEYINPUT2), .A2(G113), .ZN(new_n255));
  NAND2_X1  g069(.A1(KEYINPUT2), .A2(G113), .ZN(new_n256));
  NAND2_X1  g070(.A1(G116), .A2(G119), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  NOR2_X1   g072(.A1(G116), .A2(G119), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n255), .B(new_n256), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G116), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n188), .ZN(new_n262));
  INV_X1    g076(.A(new_n256), .ZN(new_n263));
  NOR2_X1   g077(.A1(KEYINPUT2), .A2(G113), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n262), .B(new_n257), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n260), .A2(new_n265), .A3(KEYINPUT67), .ZN(new_n266));
  AOI21_X1  g080(.A(KEYINPUT67), .B1(new_n260), .B2(new_n265), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT11), .ZN(new_n270));
  INV_X1    g084(.A(G134), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n270), .B1(new_n271), .B2(G137), .ZN(new_n272));
  INV_X1    g086(.A(G137), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n273), .A2(KEYINPUT11), .A3(G134), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n271), .A2(G137), .ZN(new_n276));
  INV_X1    g090(.A(G131), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT65), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT65), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G131), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n276), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n275), .A2(new_n281), .A3(KEYINPUT66), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT66), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n272), .A2(new_n274), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n276), .A2(new_n278), .A3(new_n280), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n276), .ZN(new_n288));
  OAI21_X1  g102(.A(G131), .B1(new_n284), .B2(new_n288), .ZN(new_n289));
  AND3_X1   g103(.A1(new_n287), .A2(KEYINPUT68), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT68), .B1(new_n287), .B2(new_n289), .ZN(new_n291));
  INV_X1    g105(.A(G143), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n292), .A2(G146), .ZN(new_n293));
  OR2_X1    g107(.A1(KEYINPUT64), .A2(G146), .ZN(new_n294));
  NAND2_X1  g108(.A1(KEYINPUT64), .A2(G146), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n293), .B1(new_n296), .B2(new_n292), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT0), .B(G128), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n294), .A2(G143), .A3(new_n295), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n216), .A2(G143), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(KEYINPUT0), .A2(G128), .ZN(new_n303));
  OAI22_X1  g117(.A1(new_n297), .A2(new_n298), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n290), .A2(new_n291), .A3(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n191), .A2(KEYINPUT1), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n299), .A2(new_n301), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n191), .B1(new_n299), .B2(KEYINPUT1), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n307), .B1(new_n308), .B2(new_n297), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n273), .A2(G134), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n277), .B1(new_n310), .B2(new_n276), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n311), .B1(new_n282), .B2(new_n286), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT69), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n309), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  AOI211_X1 g128(.A(KEYINPUT69), .B(new_n311), .C1(new_n282), .C2(new_n286), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(KEYINPUT30), .B1(new_n305), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n311), .ZN(new_n318));
  AOI21_X1  g132(.A(KEYINPUT66), .B1(new_n275), .B2(new_n281), .ZN(new_n319));
  NOR3_X1   g133(.A1(new_n284), .A2(new_n285), .A3(new_n283), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n309), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n304), .B1(new_n287), .B2(new_n289), .ZN(new_n324));
  NOR3_X1   g138(.A1(new_n323), .A2(new_n324), .A3(KEYINPUT30), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n269), .B1(new_n317), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n289), .B1(new_n319), .B2(new_n320), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT68), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n304), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n287), .A2(KEYINPUT68), .A3(new_n289), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n321), .A2(KEYINPUT69), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n312), .A2(new_n313), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(new_n309), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n333), .A2(new_n336), .A3(new_n269), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT26), .B(G101), .ZN(new_n338));
  NOR2_X1   g152(.A1(G237), .A2(G953), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G210), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n338), .B(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n342));
  XOR2_X1   g156(.A(new_n341), .B(new_n342), .Z(new_n343));
  NAND2_X1  g157(.A1(new_n337), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(KEYINPUT31), .B1(new_n327), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT28), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n337), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n268), .B1(new_n323), .B2(new_n324), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n333), .A2(new_n336), .A3(KEYINPUT28), .A4(new_n269), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n343), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n337), .A2(new_n343), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT31), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n333), .A2(new_n336), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n325), .B1(new_n355), .B2(KEYINPUT30), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n353), .B(new_n354), .C1(new_n269), .C2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n345), .A2(new_n352), .A3(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(G472), .A2(G902), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n358), .A2(KEYINPUT32), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(KEYINPUT32), .B1(new_n358), .B2(new_n359), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n337), .B1(new_n356), .B2(new_n269), .ZN(new_n363));
  AOI21_X1  g177(.A(KEYINPUT29), .B1(new_n363), .B2(new_n351), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n347), .A2(new_n349), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT71), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n365), .A2(new_n366), .A3(new_n343), .A4(new_n348), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT71), .B1(new_n350), .B2(new_n351), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n364), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT72), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n370), .B1(new_n337), .B2(new_n346), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n355), .A2(new_n268), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n347), .A2(new_n349), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n371), .B1(new_n373), .B2(new_n370), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n343), .A2(KEYINPUT29), .ZN(new_n375));
  AOI21_X1  g189(.A(G902), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n369), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G472), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n254), .B1(new_n362), .B2(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(G110), .B(G140), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n231), .A2(G227), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n380), .B(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n330), .A2(new_n332), .ZN(new_n383));
  INV_X1    g197(.A(G104), .ZN(new_n384));
  NOR3_X1   g198(.A1(new_n384), .A2(KEYINPUT3), .A3(G107), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  OR2_X1    g200(.A1(KEYINPUT80), .A2(G104), .ZN(new_n387));
  NAND2_X1  g201(.A1(KEYINPUT80), .A2(G104), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(G107), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(G107), .B1(new_n387), .B2(new_n388), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT3), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n386), .B(new_n389), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G101), .ZN(new_n393));
  INV_X1    g207(.A(G101), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n389), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G107), .ZN(new_n397));
  AND2_X1   g211(.A1(KEYINPUT80), .A2(G104), .ZN(new_n398));
  NOR2_X1   g212(.A1(KEYINPUT80), .A2(G104), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n397), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n385), .B1(new_n400), .B2(KEYINPUT3), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n393), .A2(KEYINPUT4), .A3(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n394), .A2(KEYINPUT4), .ZN(new_n404));
  AOI21_X1  g218(.A(KEYINPUT81), .B1(new_n392), .B2(new_n404), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n392), .A2(KEYINPUT81), .A3(new_n404), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n403), .B(new_n331), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n397), .A2(G104), .ZN(new_n408));
  OAI21_X1  g222(.A(G101), .B1(new_n390), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT82), .ZN(new_n410));
  INV_X1    g224(.A(new_n408), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n394), .B1(new_n400), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT82), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AOI22_X1  g228(.A1(new_n410), .A2(new_n414), .B1(new_n401), .B2(new_n396), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT10), .ZN(new_n416));
  NOR3_X1   g230(.A1(new_n225), .A2(new_n226), .A3(new_n292), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT1), .ZN(new_n418));
  OAI21_X1  g232(.A(G128), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n293), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n420), .B1(new_n227), .B2(G143), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n416), .B1(new_n422), .B2(new_n307), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n415), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n300), .B1(new_n227), .B2(G143), .ZN(new_n425));
  OAI21_X1  g239(.A(G128), .B1(new_n293), .B2(new_n418), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n307), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n412), .A2(new_n413), .ZN(new_n429));
  AOI211_X1 g243(.A(KEYINPUT82), .B(new_n394), .C1(new_n400), .C2(new_n411), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n428), .B(new_n402), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n416), .ZN(new_n432));
  AND4_X1   g246(.A1(new_n383), .A2(new_n407), .A3(new_n424), .A4(new_n432), .ZN(new_n433));
  AOI22_X1  g247(.A1(new_n416), .A2(new_n431), .B1(new_n415), .B2(new_n423), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n383), .B1(new_n434), .B2(new_n407), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n382), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT85), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n290), .A2(new_n291), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n431), .B1(new_n415), .B2(new_n309), .ZN(new_n440));
  AOI21_X1  g254(.A(KEYINPUT12), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n402), .B1(new_n429), .B2(new_n430), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n302), .A2(new_n426), .ZN(new_n443));
  AOI22_X1  g257(.A1(new_n443), .A2(new_n307), .B1(new_n396), .B2(new_n401), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n410), .A2(new_n414), .ZN(new_n445));
  AOI22_X1  g259(.A1(new_n442), .A2(new_n322), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n328), .A2(KEYINPUT12), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(KEYINPUT84), .B1(new_n441), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT12), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n450), .B1(new_n446), .B2(new_n383), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT84), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n440), .A2(KEYINPUT12), .A3(new_n328), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n434), .A2(new_n383), .A3(new_n407), .ZN(new_n455));
  INV_X1    g269(.A(new_n382), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n449), .A2(new_n454), .A3(new_n455), .A4(new_n456), .ZN(new_n457));
  OAI211_X1 g271(.A(KEYINPUT85), .B(new_n382), .C1(new_n433), .C2(new_n435), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n438), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(G469), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n460), .A3(new_n237), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n455), .B1(new_n441), .B2(new_n448), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n382), .B(KEYINPUT79), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n434), .A2(new_n407), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n439), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n455), .A3(new_n456), .ZN(new_n467));
  AOI21_X1  g281(.A(G902), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(KEYINPUT83), .B1(new_n468), .B2(new_n460), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT83), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n433), .A2(new_n435), .ZN(new_n471));
  AOI22_X1  g285(.A1(new_n471), .A2(new_n456), .B1(new_n462), .B2(new_n463), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n470), .B(G469), .C1(new_n472), .C2(G902), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n461), .A2(new_n469), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(G214), .B1(G237), .B2(G902), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(G110), .B(G122), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(KEYINPUT8), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n262), .A2(new_n257), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT5), .ZN(new_n480));
  INV_X1    g294(.A(G113), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n261), .A2(KEYINPUT5), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n481), .B1(new_n482), .B2(new_n188), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n263), .A2(new_n264), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n480), .A2(new_n483), .B1(new_n484), .B2(new_n479), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n485), .B1(new_n445), .B2(new_n402), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n402), .B(new_n485), .C1(new_n429), .C2(new_n430), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n478), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT87), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT87), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n491), .B(new_n478), .C1(new_n486), .C2(new_n488), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n406), .A2(new_n405), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n386), .B1(new_n390), .B2(new_n391), .ZN(new_n495));
  OAI21_X1  g309(.A(KEYINPUT4), .B1(new_n495), .B2(new_n395), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n394), .B1(new_n401), .B2(new_n389), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n268), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n477), .B(new_n487), .C1(new_n494), .C2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n422), .A2(new_n208), .A3(new_n307), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n304), .A2(G125), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT88), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT7), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n500), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n231), .A2(G224), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT7), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n506), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n500), .A2(new_n501), .A3(new_n508), .A4(new_n503), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n499), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(G902), .B1(new_n493), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n487), .B1(new_n494), .B2(new_n498), .ZN(new_n512));
  INV_X1    g326(.A(new_n477), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(KEYINPUT6), .A3(new_n499), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n500), .A2(new_n501), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n505), .B(KEYINPUT86), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n516), .B(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT6), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n512), .A2(new_n519), .A3(new_n513), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n515), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n511), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(G210), .B1(G237), .B2(G902), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n511), .A2(new_n523), .A3(new_n521), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n476), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(G221), .ZN(new_n528));
  XOR2_X1   g342(.A(KEYINPUT9), .B(G234), .Z(new_n529));
  AOI21_X1  g343(.A(new_n528), .B1(new_n529), .B2(new_n237), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n474), .A2(new_n527), .A3(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT93), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n278), .A2(new_n280), .ZN(new_n535));
  OR2_X1    g349(.A1(KEYINPUT89), .A2(G143), .ZN(new_n536));
  NAND2_X1  g350(.A1(KEYINPUT89), .A2(G143), .ZN(new_n537));
  AOI22_X1  g351(.A1(new_n536), .A2(new_n537), .B1(new_n339), .B2(G214), .ZN(new_n538));
  INV_X1    g352(.A(G237), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n539), .A2(new_n231), .A3(G214), .ZN(new_n540));
  NOR2_X1   g354(.A1(KEYINPUT89), .A2(G143), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n535), .B1(new_n538), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n537), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n540), .B1(new_n544), .B2(new_n541), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n278), .A2(new_n280), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n536), .A2(G214), .A3(new_n339), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT17), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n543), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  OAI211_X1 g364(.A(KEYINPUT17), .B(new_n535), .C1(new_n538), .C2(new_n542), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n217), .A2(new_n550), .A3(new_n218), .A4(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(G113), .B(G122), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(new_n384), .ZN(new_n554));
  NAND2_X1  g368(.A1(KEYINPUT18), .A2(G131), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n545), .A2(new_n555), .A3(new_n547), .ZN(new_n556));
  OAI211_X1 g370(.A(KEYINPUT18), .B(G131), .C1(new_n538), .C2(new_n542), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n227), .A2(new_n207), .A3(new_n209), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n210), .A2(G146), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n558), .A2(KEYINPUT90), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(KEYINPUT90), .B1(new_n558), .B2(new_n559), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n556), .B(new_n557), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n552), .A2(new_n554), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(KEYINPUT91), .A2(KEYINPUT19), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n224), .A2(new_n564), .ZN(new_n565));
  OR2_X1    g379(.A1(KEYINPUT91), .A2(KEYINPUT19), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n566), .A2(new_n564), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n565), .B(new_n227), .C1(new_n224), .C2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n543), .A2(new_n548), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(new_n569), .A3(new_n218), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n554), .B1(new_n562), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT92), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n563), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AOI211_X1 g387(.A(KEYINPUT92), .B(new_n554), .C1(new_n562), .C2(new_n570), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n534), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT20), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(G475), .A2(G902), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n578), .B1(new_n573), .B2(new_n574), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n562), .A2(new_n570), .ZN(new_n581));
  OAI21_X1  g395(.A(KEYINPUT92), .B1(new_n581), .B2(new_n554), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n571), .A2(new_n572), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n582), .A2(new_n583), .A3(new_n563), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n584), .A2(KEYINPUT93), .A3(new_n576), .A4(new_n578), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n563), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT94), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n552), .A2(new_n562), .ZN(new_n589));
  INV_X1    g403(.A(new_n554), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n589), .A2(new_n588), .A3(new_n590), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n587), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(G475), .B1(new_n594), .B2(G902), .ZN(new_n595));
  INV_X1    g409(.A(G478), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(KEYINPUT15), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT96), .ZN(new_n599));
  XOR2_X1   g413(.A(G116), .B(G122), .Z(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(G107), .ZN(new_n601));
  XNOR2_X1  g415(.A(G116), .B(G122), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n397), .ZN(new_n603));
  XNOR2_X1  g417(.A(G128), .B(G143), .ZN(new_n604));
  AOI22_X1  g418(.A1(new_n601), .A2(new_n603), .B1(new_n271), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(KEYINPUT13), .ZN(new_n606));
  NOR3_X1   g420(.A1(new_n191), .A2(KEYINPUT13), .A3(G143), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n607), .A2(new_n271), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT95), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n606), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n609), .B1(new_n606), .B2(new_n608), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n605), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n604), .B(new_n271), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n261), .A2(KEYINPUT14), .A3(G122), .ZN(new_n614));
  OAI211_X1 g428(.A(G107), .B(new_n614), .C1(new_n600), .C2(KEYINPUT14), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n613), .A2(new_n603), .A3(new_n615), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n529), .A2(new_n231), .A3(new_n243), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n612), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n617), .B1(new_n612), .B2(new_n616), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n599), .B1(new_n620), .B2(G902), .ZN(new_n621));
  OAI211_X1 g435(.A(KEYINPUT96), .B(new_n237), .C1(new_n618), .C2(new_n619), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n598), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n231), .A2(G952), .ZN(new_n624));
  NAND2_X1  g438(.A1(G234), .A2(G237), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n625), .A2(G902), .A3(G953), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(KEYINPUT21), .B(G898), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n627), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n620), .A2(G902), .A3(new_n597), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n623), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n586), .A2(new_n595), .A3(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n379), .A2(new_n533), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(KEYINPUT97), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G101), .ZN(G3));
  NAND2_X1  g452(.A1(new_n358), .A2(new_n237), .ZN(new_n639));
  AOI22_X1  g453(.A1(new_n639), .A2(G472), .B1(new_n358), .B2(new_n359), .ZN(new_n640));
  INV_X1    g454(.A(new_n254), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n640), .A2(new_n531), .A3(new_n474), .A4(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n631), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n621), .A2(new_n622), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n596), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT98), .ZN(new_n646));
  OAI21_X1  g460(.A(KEYINPUT33), .B1(new_n618), .B2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(new_n620), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n648), .A2(G478), .A3(new_n237), .ZN(new_n649));
  AOI22_X1  g463(.A1(new_n586), .A2(new_n595), .B1(new_n645), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n527), .A2(new_n643), .A3(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n642), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(KEYINPUT34), .B(G104), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G6));
  XNOR2_X1  g468(.A(new_n579), .B(new_n576), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n623), .A2(new_n632), .ZN(new_n656));
  INV_X1    g470(.A(G475), .ZN(new_n657));
  INV_X1    g471(.A(new_n593), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n563), .B1(new_n658), .B2(new_n591), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n657), .B1(new_n659), .B2(new_n237), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n655), .A2(new_n656), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n527), .A2(new_n643), .A3(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n642), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT35), .B(G107), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G9));
  AOI21_X1  g479(.A(new_n246), .B1(new_n239), .B2(KEYINPUT25), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT99), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n667), .B1(new_n220), .B2(new_n229), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n235), .A2(KEYINPUT36), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n220), .A2(new_n667), .A3(new_n229), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n229), .ZN(new_n673));
  AOI211_X1 g487(.A(KEYINPUT99), .B(new_n673), .C1(new_n200), .C2(new_n219), .ZN(new_n674));
  OAI22_X1  g488(.A1(new_n668), .A2(new_n674), .B1(KEYINPUT36), .B2(new_n235), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  AOI22_X1  g490(.A1(new_n666), .A2(new_n242), .B1(new_n676), .B2(new_n250), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n634), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n640), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n679), .A2(new_n532), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT37), .B(G110), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G12));
  NAND2_X1  g496(.A1(new_n358), .A2(new_n359), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT32), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n358), .A2(KEYINPUT32), .A3(new_n359), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n378), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n474), .A2(new_n531), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n676), .A2(new_n250), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n248), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n523), .B1(new_n511), .B2(new_n521), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n511), .A2(new_n523), .A3(new_n521), .ZN(new_n693));
  OAI211_X1 g507(.A(new_n691), .B(new_n475), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT100), .B(G900), .Z(new_n695));
  AOI21_X1  g509(.A(new_n627), .B1(new_n629), .B2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n661), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n689), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G128), .ZN(G30));
  XOR2_X1   g515(.A(new_n696), .B(KEYINPUT39), .Z(new_n702));
  NAND2_X1  g516(.A1(new_n688), .A2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT40), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n363), .A2(new_n343), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n372), .A2(new_n351), .A3(new_n337), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n237), .ZN(new_n708));
  OAI21_X1  g522(.A(G472), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n685), .A2(new_n709), .A3(new_n686), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n693), .A2(new_n692), .ZN(new_n711));
  XOR2_X1   g525(.A(new_n711), .B(KEYINPUT38), .Z(new_n712));
  INV_X1    g526(.A(new_n585), .ZN(new_n713));
  AOI22_X1  g527(.A1(new_n575), .A2(new_n576), .B1(new_n584), .B2(new_n578), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n595), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n656), .A2(new_n476), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n677), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n705), .A2(new_n710), .A3(new_n712), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(KEYINPUT101), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G143), .ZN(G45));
  NAND2_X1  g534(.A1(new_n649), .A2(new_n645), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n715), .A2(new_n721), .A3(new_n697), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n694), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n689), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G146), .ZN(G48));
  INV_X1    g539(.A(KEYINPUT102), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n685), .A2(new_n686), .ZN(new_n727));
  INV_X1    g541(.A(G472), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n728), .B1(new_n369), .B2(new_n376), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n641), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n459), .A2(new_n460), .A3(new_n237), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n460), .B1(new_n459), .B2(new_n237), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n731), .A2(new_n732), .A3(new_n530), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n475), .B(new_n643), .C1(new_n693), .C2(new_n692), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n715), .A2(new_n721), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n726), .B1(new_n730), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n459), .A2(new_n237), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(G469), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n531), .A3(new_n461), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n741), .A2(new_n651), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n379), .A2(new_n742), .A3(KEYINPUT102), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n738), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(KEYINPUT41), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G113), .ZN(G15));
  NOR2_X1   g560(.A1(new_n741), .A2(new_n662), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n379), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G116), .ZN(G18));
  AND4_X1   g563(.A1(new_n527), .A2(new_n740), .A3(new_n531), .A4(new_n461), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n687), .A2(new_n750), .A3(new_n678), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G119), .ZN(G21));
  OAI211_X1 g566(.A(new_n715), .B(new_n716), .C1(new_n693), .C2(new_n692), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n753), .A2(new_n631), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n733), .ZN(new_n755));
  INV_X1    g569(.A(new_n359), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n373), .A2(new_n370), .ZN(new_n757));
  INV_X1    g571(.A(new_n371), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n351), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n345), .A2(new_n357), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n756), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n728), .B1(new_n358), .B2(new_n237), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n763), .A2(new_n641), .A3(new_n765), .ZN(new_n766));
  OAI21_X1  g580(.A(KEYINPUT103), .B1(new_n755), .B2(new_n766), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n762), .A2(new_n254), .A3(new_n764), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT103), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n768), .A2(new_n769), .A3(new_n733), .A4(new_n754), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G122), .ZN(G24));
  NOR3_X1   g586(.A1(new_n762), .A2(new_n764), .A3(new_n677), .ZN(new_n773));
  INV_X1    g587(.A(new_n722), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n750), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G125), .ZN(G27));
  OAI21_X1  g590(.A(G469), .B1(new_n472), .B2(G902), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n461), .A2(new_n777), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n693), .A2(new_n692), .A3(new_n476), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n778), .A2(new_n531), .A3(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n379), .A2(new_n774), .A3(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT42), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT104), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n729), .B1(new_n783), .B2(new_n685), .ZN(new_n784));
  OAI21_X1  g598(.A(KEYINPUT104), .B1(new_n360), .B2(new_n361), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n254), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n530), .B1(new_n461), .B2(new_n777), .ZN(new_n787));
  AND4_X1   g601(.A1(KEYINPUT42), .A2(new_n787), .A3(new_n774), .A4(new_n779), .ZN(new_n788));
  AOI22_X1  g602(.A1(new_n781), .A2(new_n782), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(new_n277), .ZN(G33));
  INV_X1    g604(.A(new_n698), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n687), .A2(new_n780), .A3(new_n641), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(KEYINPUT105), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT105), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n379), .A2(new_n794), .A3(new_n791), .A4(new_n780), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G134), .ZN(G36));
  INV_X1    g611(.A(new_n779), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n472), .A2(KEYINPUT45), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n472), .A2(KEYINPUT45), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n799), .A2(G469), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(G469), .A2(G902), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT46), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n731), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n805), .B1(new_n804), .B2(new_n803), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(new_n531), .A3(new_n702), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT44), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n586), .A2(new_n721), .A3(new_n595), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT106), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n809), .A2(new_n810), .A3(KEYINPUT43), .ZN(new_n811));
  AOI21_X1  g625(.A(KEYINPUT43), .B1(new_n809), .B2(new_n810), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n640), .A2(new_n677), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT107), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n814), .A2(new_n815), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n813), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AOI211_X1 g633(.A(new_n798), .B(new_n807), .C1(new_n808), .C2(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n820), .B1(new_n808), .B2(new_n819), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(G137), .ZN(G39));
  INV_X1    g636(.A(KEYINPUT47), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n806), .A2(new_n823), .A3(new_n531), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n823), .B1(new_n806), .B2(new_n531), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n774), .A2(new_n254), .A3(new_n779), .ZN(new_n826));
  OR4_X1    g640(.A1(new_n687), .A2(new_n824), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(G140), .ZN(G42));
  NOR4_X1   g642(.A1(new_n809), .A2(new_n254), .A3(new_n476), .A4(new_n530), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n830), .A2(KEYINPUT108), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n831), .A2(new_n710), .A3(new_n712), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n740), .A2(new_n461), .ZN(new_n833));
  AOI22_X1  g647(.A1(new_n830), .A2(KEYINPUT108), .B1(KEYINPUT49), .B2(new_n833), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n832), .B(new_n834), .C1(KEYINPUT49), .C2(new_n833), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n710), .A2(new_n254), .A3(new_n626), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n741), .A2(new_n798), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n624), .B1(new_n838), .B2(new_n735), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n811), .A2(new_n812), .A3(new_n626), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n786), .A2(new_n840), .A3(new_n837), .ZN(new_n841));
  XOR2_X1   g655(.A(new_n841), .B(KEYINPUT48), .Z(new_n842));
  AND2_X1   g656(.A1(new_n840), .A2(new_n768), .ZN(new_n843));
  AOI211_X1 g657(.A(new_n839), .B(new_n842), .C1(new_n750), .C2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n840), .A2(new_n773), .A3(new_n837), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(KEYINPUT116), .ZN(new_n846));
  OR3_X1    g660(.A1(new_n838), .A2(new_n715), .A3(new_n721), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n712), .A2(new_n475), .A3(new_n741), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n843), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT50), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n849), .A2(KEYINPUT115), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n850), .B1(new_n849), .B2(KEYINPUT115), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n846), .B(new_n847), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n531), .B1(new_n833), .B2(KEYINPUT114), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n854), .B1(KEYINPUT114), .B2(new_n833), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n855), .B1(new_n824), .B2(new_n825), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n856), .A2(new_n779), .A3(new_n843), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n853), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n844), .B1(new_n859), .B2(KEYINPUT51), .ZN(new_n860));
  OR2_X1    g674(.A1(new_n851), .A2(new_n852), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n846), .A2(new_n847), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n861), .A2(KEYINPUT51), .A3(new_n857), .A4(new_n862), .ZN(new_n863));
  OR2_X1    g677(.A1(new_n863), .A2(KEYINPUT117), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(KEYINPUT117), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n860), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT113), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n868));
  INV_X1    g682(.A(new_n678), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n869), .B1(new_n362), .B2(new_n378), .ZN(new_n870));
  AOI22_X1  g684(.A1(new_n870), .A2(new_n750), .B1(new_n379), .B2(new_n747), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n744), .A2(new_n771), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n735), .B1(new_n715), .B2(new_n656), .ZN(new_n873));
  INV_X1    g687(.A(new_n734), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI22_X1  g689(.A1(new_n642), .A2(new_n875), .B1(new_n679), .B2(new_n532), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT109), .B1(new_n877), .B2(new_n636), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n872), .A2(new_n878), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n687), .B(new_n688), .C1(new_n699), .C2(new_n723), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n696), .B(KEYINPUT111), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT112), .B1(new_n677), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n882), .A2(new_n753), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n677), .A2(KEYINPUT112), .A3(new_n881), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n883), .A2(new_n710), .A3(new_n787), .A4(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n880), .A2(new_n775), .A3(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT52), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n880), .A2(KEYINPUT52), .A3(new_n775), .A4(new_n885), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n789), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n877), .A2(KEYINPUT109), .A3(new_n636), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n879), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n655), .A2(new_n660), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n691), .A2(new_n893), .A3(new_n656), .A4(new_n697), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n798), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n687), .A2(new_n688), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n780), .A2(new_n773), .A3(new_n774), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI211_X1 g712(.A(KEYINPUT110), .B(new_n898), .C1(new_n795), .C2(new_n793), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT110), .ZN(new_n900));
  INV_X1    g714(.A(new_n898), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n900), .B1(new_n796), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n868), .B1(new_n892), .B2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT54), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n898), .B1(new_n793), .B2(new_n795), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(new_n900), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n730), .A2(new_n532), .A3(new_n634), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT109), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n908), .A2(new_n876), .A3(new_n909), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n872), .A2(new_n878), .A3(new_n910), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n907), .A2(new_n911), .A3(KEYINPUT53), .A4(new_n890), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n904), .A2(new_n905), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n905), .B1(new_n904), .B2(new_n912), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n867), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n888), .A2(new_n889), .ZN(new_n916));
  INV_X1    g730(.A(new_n789), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n748), .A2(new_n751), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n919), .B1(new_n770), .B2(new_n767), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n909), .B1(new_n908), .B2(new_n876), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n920), .A2(new_n744), .A3(new_n891), .A4(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n918), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(KEYINPUT53), .B1(new_n923), .B2(new_n907), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n892), .A2(new_n903), .A3(new_n868), .ZN(new_n925));
  OAI21_X1  g739(.A(KEYINPUT54), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n904), .A2(new_n905), .A3(new_n912), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n926), .A2(KEYINPUT113), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n866), .A2(new_n915), .A3(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT118), .ZN(new_n930));
  OAI22_X1  g744(.A1(new_n929), .A2(new_n930), .B1(G952), .B2(G953), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n929), .A2(new_n930), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n835), .B1(new_n931), .B2(new_n932), .ZN(G75));
  NAND2_X1  g747(.A1(new_n515), .A2(new_n520), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(new_n518), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT55), .Z(new_n936));
  AOI21_X1  g750(.A(new_n237), .B1(new_n904), .B2(new_n912), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n937), .A2(G210), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n936), .B1(new_n938), .B2(KEYINPUT56), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n231), .A2(G952), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n937), .A2(G210), .ZN(new_n941));
  XOR2_X1   g755(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n942));
  NOR2_X1   g756(.A1(new_n936), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n940), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n939), .A2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT120), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(G51));
  NAND2_X1  g761(.A1(new_n926), .A2(new_n927), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n802), .B(KEYINPUT57), .Z(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n459), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n937), .A2(G469), .A3(new_n800), .A4(new_n799), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n940), .B1(new_n951), .B2(new_n952), .ZN(G54));
  NAND3_X1  g767(.A1(new_n937), .A2(KEYINPUT58), .A3(G475), .ZN(new_n954));
  INV_X1    g768(.A(new_n584), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n954), .A2(new_n955), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n956), .A2(new_n957), .A3(new_n940), .ZN(G60));
  NAND2_X1  g772(.A1(G478), .A2(G902), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT59), .Z(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n913), .A2(new_n914), .A3(new_n867), .ZN(new_n962));
  AOI21_X1  g776(.A(KEYINPUT113), .B1(new_n926), .B2(new_n927), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT122), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n648), .B(KEYINPUT121), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n964), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n960), .B1(new_n915), .B2(new_n928), .ZN(new_n969));
  OAI21_X1  g783(.A(KEYINPUT122), .B1(new_n969), .B2(new_n966), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n967), .A2(new_n960), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n940), .B1(new_n948), .B2(new_n971), .ZN(new_n972));
  AND3_X1   g786(.A1(new_n968), .A2(new_n970), .A3(new_n972), .ZN(G63));
  NAND2_X1  g787(.A1(G217), .A2(G902), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT60), .Z(new_n975));
  OAI21_X1  g789(.A(new_n975), .B1(new_n924), .B2(new_n925), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n940), .B1(new_n976), .B2(new_n249), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n676), .B(KEYINPUT123), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n977), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT61), .Z(G66));
  NAND2_X1  g794(.A1(G224), .A2(G953), .ZN(new_n981));
  OAI22_X1  g795(.A1(new_n922), .A2(G953), .B1(new_n630), .B2(new_n981), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT124), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n934), .B1(G898), .B2(new_n231), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n983), .B(new_n984), .ZN(G69));
  AND2_X1   g799(.A1(new_n880), .A2(new_n775), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n719), .A2(new_n986), .ZN(new_n987));
  OR2_X1    g801(.A1(new_n987), .A2(KEYINPUT62), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(KEYINPUT62), .ZN(new_n989));
  INV_X1    g803(.A(new_n703), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n990), .A2(new_n379), .A3(new_n779), .A4(new_n873), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n821), .A2(new_n827), .A3(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n988), .A2(new_n989), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(new_n231), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n224), .A2(new_n567), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n995), .B1(new_n224), .B2(new_n564), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n356), .B(new_n996), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(KEYINPUT125), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n994), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n231), .B1(G227), .B2(G900), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT127), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(new_n753), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n786), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n986), .B1(new_n807), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n1006), .A2(new_n789), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n821), .A2(new_n796), .A3(new_n827), .A4(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1008), .A2(new_n231), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n231), .A2(G900), .ZN(new_n1010));
  XOR2_X1   g824(.A(new_n1010), .B(KEYINPUT126), .Z(new_n1011));
  NAND2_X1  g825(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(new_n997), .ZN(new_n1013));
  AOI22_X1  g827(.A1(new_n1012), .A2(new_n1013), .B1(new_n1001), .B2(new_n1000), .ZN(new_n1014));
  AND3_X1   g828(.A1(new_n999), .A2(new_n1003), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1003), .B1(new_n999), .B2(new_n1014), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n1015), .A2(new_n1016), .ZN(G72));
  INV_X1    g831(.A(new_n706), .ZN(new_n1018));
  OR2_X1    g832(.A1(new_n993), .A2(new_n922), .ZN(new_n1019));
  NAND2_X1  g833(.A1(G472), .A2(G902), .ZN(new_n1020));
  XOR2_X1   g834(.A(new_n1020), .B(KEYINPUT63), .Z(new_n1021));
  AOI21_X1  g835(.A(new_n1018), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n363), .A2(new_n343), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1024));
  AOI211_X1 g838(.A(new_n1023), .B(new_n1024), .C1(new_n904), .C2(new_n912), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1021), .B1(new_n1008), .B2(new_n922), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1026), .A2(new_n1023), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1027), .B1(G952), .B2(new_n231), .ZN(new_n1028));
  NOR3_X1   g842(.A1(new_n1022), .A2(new_n1025), .A3(new_n1028), .ZN(G57));
endmodule


