//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 1 0 1 0 0 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1 1 1 0 1 0 1 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n999, new_n1000, new_n1001, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1024, new_n1025;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT16), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(G1gat), .B2(new_n202), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(G8gat), .ZN(new_n207));
  INV_X1    g006(.A(G43gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G50gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT15), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n208), .A2(G50gat), .ZN(new_n212));
  NOR3_X1   g011(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT89), .B(KEYINPUT15), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT90), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n212), .B1(new_n216), .B2(new_n209), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n208), .A2(KEYINPUT90), .A3(G50gat), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n215), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT14), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(G29gat), .B2(G36gat), .ZN(new_n221));
  INV_X1    g020(.A(G29gat), .ZN(new_n222));
  INV_X1    g021(.A(G36gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(new_n223), .A3(KEYINPUT14), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT88), .B(G36gat), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n221), .B(new_n224), .C1(new_n225), .C2(new_n222), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n214), .B1(new_n219), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n224), .A2(new_n221), .ZN(new_n228));
  INV_X1    g027(.A(new_n225), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n228), .B1(new_n229), .B2(G29gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(new_n213), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n207), .B1(new_n232), .B2(KEYINPUT17), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT91), .ZN(new_n234));
  INV_X1    g033(.A(G50gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n216), .B1(new_n235), .B2(G43gat), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n236), .B(new_n218), .C1(new_n208), .C2(G50gat), .ZN(new_n237));
  INV_X1    g036(.A(new_n215), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n213), .B1(new_n230), .B2(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n214), .A2(new_n226), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n234), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n227), .A2(KEYINPUT91), .A3(new_n231), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT17), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n233), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(G229gat), .A2(G233gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n242), .A2(new_n243), .A3(new_n207), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT92), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(KEYINPUT18), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT18), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n249), .A2(KEYINPUT92), .A3(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n247), .B(KEYINPUT13), .Z(new_n254));
  NAND2_X1  g053(.A1(new_n242), .A2(new_n243), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n256), .A2(new_n207), .ZN(new_n257));
  INV_X1    g056(.A(new_n248), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n254), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n251), .A2(new_n253), .A3(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G113gat), .B(G141gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n261), .B(G197gat), .ZN(new_n262));
  XOR2_X1   g061(.A(KEYINPUT11), .B(G169gat), .Z(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(KEYINPUT12), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n251), .A2(new_n253), .A3(new_n265), .A4(new_n259), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G155gat), .ZN(new_n271));
  INV_X1    g070(.A(G162gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(G155gat), .A2(G162gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G148gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(G141gat), .ZN(new_n277));
  INV_X1    g076(.A(G141gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(G148gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT2), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n275), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT77), .ZN(new_n283));
  AND3_X1   g082(.A1(new_n277), .A2(new_n279), .A3(KEYINPUT76), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT76), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n285), .A2(new_n276), .A3(G141gat), .ZN(new_n286));
  NOR3_X1   g085(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n287));
  INV_X1    g086(.A(new_n274), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n283), .B1(new_n284), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n274), .B1(new_n273), .B2(KEYINPUT2), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n277), .A2(new_n279), .A3(KEYINPUT76), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n291), .A2(new_n292), .A3(KEYINPUT77), .A4(new_n286), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n282), .B1(new_n290), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT3), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT29), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(G197gat), .B(G204gat), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT22), .ZN(new_n298));
  INV_X1    g097(.A(G211gat), .ZN(new_n299));
  INV_X1    g098(.A(G218gat), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(G211gat), .B(G218gat), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n303), .A2(new_n297), .A3(new_n301), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n305), .A2(KEYINPUT74), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT74), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n302), .A2(new_n308), .A3(new_n304), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n296), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT29), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n307), .A2(new_n313), .A3(new_n309), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n294), .B1(new_n314), .B2(new_n295), .ZN(new_n315));
  NAND2_X1  g114(.A1(G228gat), .A2(G233gat), .ZN(new_n316));
  NOR3_X1   g115(.A1(new_n312), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n305), .A2(new_n306), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT3), .B1(new_n319), .B2(new_n313), .ZN(new_n320));
  OAI22_X1  g119(.A1(new_n296), .A2(new_n311), .B1(new_n294), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT81), .ZN(new_n322));
  XOR2_X1   g121(.A(new_n316), .B(KEYINPUT80), .Z(new_n323));
  NAND3_X1  g122(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n322), .B1(new_n321), .B2(new_n323), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n318), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  XOR2_X1   g126(.A(KEYINPUT31), .B(G50gat), .Z(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G78gat), .B(G106gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(G22gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n321), .A2(new_n323), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT81), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(new_n324), .ZN(new_n334));
  INV_X1    g133(.A(new_n328), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n334), .A2(new_n335), .A3(new_n318), .ZN(new_n336));
  AND3_X1   g135(.A1(new_n329), .A2(new_n331), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n331), .B1(new_n329), .B2(new_n336), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(G169gat), .A2(G176gat), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NOR2_X1   g140(.A1(G169gat), .A2(G176gat), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n341), .B1(new_n343), .B2(KEYINPUT26), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n344), .B1(KEYINPUT26), .B2(new_n343), .ZN(new_n345));
  NAND2_X1  g144(.A1(G183gat), .A2(G190gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT27), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n349), .A2(G183gat), .ZN(new_n350));
  INV_X1    g149(.A(G183gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n351), .A2(KEYINPUT27), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT28), .ZN(new_n353));
  NOR4_X1   g152(.A1(new_n350), .A2(new_n352), .A3(new_n353), .A4(G190gat), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT68), .B1(new_n350), .B2(new_n352), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n351), .A2(KEYINPUT27), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT68), .ZN(new_n358));
  AOI21_X1  g157(.A(G190gat), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT28), .B1(new_n356), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n355), .B1(new_n360), .B2(KEYINPUT69), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n349), .A2(G183gat), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n358), .B1(new_n357), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n358), .B1(new_n349), .B2(G183gat), .ZN(new_n364));
  INV_X1    g163(.A(G190gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI211_X1 g165(.A(KEYINPUT69), .B(new_n353), .C1(new_n363), .C2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n348), .B1(new_n361), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT25), .ZN(new_n370));
  INV_X1    g169(.A(G169gat), .ZN(new_n371));
  INV_X1    g170(.A(G176gat), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n371), .A2(new_n372), .A3(KEYINPUT23), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(new_n340), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT65), .B1(new_n342), .B2(KEYINPUT23), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT65), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT23), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n376), .B(new_n377), .C1(G169gat), .C2(G176gat), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n374), .B1(new_n375), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT67), .ZN(new_n381));
  OR2_X1    g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n346), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n380), .A2(new_n381), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n382), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n370), .B1(new_n379), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n384), .A2(new_n380), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(new_n370), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n375), .A2(new_n378), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n377), .A2(G176gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n371), .A2(KEYINPUT64), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT64), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(G169gat), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n391), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n390), .A2(new_n340), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT66), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n389), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n390), .A2(KEYINPUT66), .A3(new_n340), .A4(new_n395), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n387), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT29), .B1(new_n369), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(G226gat), .A2(G233gat), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(KEYINPUT75), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n402), .B1(new_n369), .B2(new_n400), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n375), .A2(new_n378), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n395), .A2(new_n340), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n397), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n389), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(new_n399), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n387), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n353), .B1(new_n363), .B2(new_n366), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT69), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n354), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n347), .B1(new_n415), .B2(new_n367), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n313), .B1(new_n412), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n405), .B1(new_n402), .B2(new_n417), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n311), .B(new_n404), .C1(new_n418), .C2(KEYINPUT75), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n403), .B1(new_n412), .B2(new_n416), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n420), .B1(new_n401), .B2(new_n403), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n310), .ZN(new_n422));
  XNOR2_X1  g221(.A(G8gat), .B(G36gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(G64gat), .B(G92gat), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n423), .B(new_n424), .Z(new_n425));
  NAND3_X1  g224(.A1(new_n419), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT30), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n419), .A2(KEYINPUT30), .A3(new_n422), .A4(new_n425), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n419), .A2(new_n422), .ZN(new_n430));
  INV_X1    g229(.A(new_n425), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n428), .A2(new_n429), .A3(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT79), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n290), .A2(new_n293), .ZN(new_n436));
  INV_X1    g235(.A(new_n282), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n438), .A2(KEYINPUT78), .A3(KEYINPUT3), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT78), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n440), .B1(new_n294), .B2(new_n295), .ZN(new_n441));
  XOR2_X1   g240(.A(G127gat), .B(G134gat), .Z(new_n442));
  XNOR2_X1  g241(.A(G113gat), .B(G120gat), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n442), .B1(KEYINPUT1), .B2(new_n443), .ZN(new_n444));
  XOR2_X1   g243(.A(G113gat), .B(G120gat), .Z(new_n445));
  INV_X1    g244(.A(KEYINPUT1), .ZN(new_n446));
  XNOR2_X1  g245(.A(G127gat), .B(G134gat), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  AND2_X1   g247(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n449), .B1(new_n294), .B2(new_n295), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n439), .A2(new_n441), .A3(new_n450), .ZN(new_n451));
  AND4_X1   g250(.A1(KEYINPUT4), .A2(new_n436), .A3(new_n437), .A4(new_n449), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT4), .B1(new_n294), .B2(new_n449), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(G225gat), .A2(G233gat), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n451), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT5), .ZN(new_n457));
  INV_X1    g256(.A(new_n449), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n438), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n294), .A2(new_n449), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n455), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n457), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n456), .A2(new_n463), .ZN(new_n464));
  XOR2_X1   g263(.A(G1gat), .B(G29gat), .Z(new_n465));
  XNOR2_X1  g264(.A(new_n465), .B(KEYINPUT0), .ZN(new_n466));
  XNOR2_X1  g265(.A(G57gat), .B(G85gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n466), .B(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n451), .A2(new_n454), .A3(new_n457), .A4(new_n455), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n464), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT6), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n468), .B1(new_n464), .B2(new_n469), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n435), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n473), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n475), .A2(KEYINPUT79), .A3(new_n471), .A4(new_n470), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n464), .A2(new_n469), .ZN(new_n477));
  INV_X1    g276(.A(new_n468), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(KEYINPUT6), .A3(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n474), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n339), .B1(new_n434), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n458), .B1(new_n412), .B2(new_n416), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n369), .A2(new_n400), .A3(new_n449), .ZN(new_n483));
  INV_X1    g282(.A(G227gat), .ZN(new_n484));
  INV_X1    g283(.A(G233gat), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n482), .A2(new_n483), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(KEYINPUT72), .A2(KEYINPUT34), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  OR2_X1    g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g290(.A1(KEYINPUT72), .A2(KEYINPUT34), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n488), .B1(new_n492), .B2(new_n490), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  XOR2_X1   g293(.A(G71gat), .B(G99gat), .Z(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(KEYINPUT71), .ZN(new_n496));
  XNOR2_X1  g295(.A(G15gat), .B(G43gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n497), .B(KEYINPUT70), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n496), .B(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n487), .B1(new_n482), .B2(new_n483), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n499), .B1(new_n500), .B2(KEYINPUT33), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT32), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n482), .A2(new_n483), .ZN(new_n505));
  AOI221_X4 g304(.A(new_n502), .B1(KEYINPUT33), .B2(new_n499), .C1(new_n505), .C2(new_n486), .ZN(new_n506));
  OAI211_X1 g305(.A(KEYINPUT73), .B(new_n494), .C1(new_n504), .C2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NOR3_X1   g307(.A1(new_n412), .A2(new_n416), .A3(new_n458), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n449), .B1(new_n369), .B2(new_n400), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n486), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT32), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT33), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n512), .A2(new_n514), .A3(new_n499), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n501), .A2(new_n503), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n494), .B1(new_n517), .B2(KEYINPUT73), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT36), .B1(new_n508), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n494), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n515), .A2(new_n494), .A3(new_n516), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT36), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n481), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n426), .A2(new_n479), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n310), .B(new_n404), .C1(new_n418), .C2(KEYINPUT75), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n529), .B(KEYINPUT37), .C1(new_n418), .C2(new_n310), .ZN(new_n530));
  OR2_X1    g329(.A1(new_n425), .A2(KEYINPUT38), .ZN(new_n531));
  XOR2_X1   g330(.A(KEYINPUT86), .B(KEYINPUT37), .Z(new_n532));
  AND2_X1   g331(.A1(new_n422), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n531), .B1(new_n533), .B2(new_n419), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n528), .B1(new_n530), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n419), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(new_n431), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT37), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n538), .B1(new_n419), .B2(new_n422), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT38), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n477), .A2(KEYINPUT84), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT84), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n464), .A2(new_n542), .A3(new_n469), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n468), .B(KEYINPUT82), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n541), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n472), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n545), .A2(KEYINPUT85), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT85), .B1(new_n545), .B2(new_n546), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n535), .B(new_n540), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n331), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n335), .B1(new_n334), .B2(new_n318), .ZN(new_n551));
  AOI211_X1 g350(.A(new_n328), .B(new_n317), .C1(new_n333), .C2(new_n324), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n329), .A2(new_n331), .A3(new_n336), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n455), .B1(new_n451), .B2(new_n454), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n459), .A2(new_n455), .A3(new_n460), .ZN(new_n557));
  AND3_X1   g356(.A1(new_n557), .A2(KEYINPUT83), .A3(KEYINPUT39), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT83), .B1(new_n557), .B2(KEYINPUT39), .ZN(new_n559));
  NOR3_X1   g358(.A1(new_n556), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT39), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n544), .B1(new_n556), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n561), .A2(KEYINPUT40), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT40), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n556), .A2(new_n562), .ZN(new_n566));
  INV_X1    g365(.A(new_n544), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n565), .B1(new_n568), .B2(new_n560), .ZN(new_n569));
  AND3_X1   g368(.A1(new_n545), .A2(new_n564), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n555), .B1(new_n570), .B2(new_n433), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n549), .A2(new_n571), .A3(KEYINPUT87), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT87), .B1(new_n549), .B2(new_n571), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n527), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n522), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n494), .B1(new_n515), .B2(new_n516), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NOR4_X1   g376(.A1(new_n577), .A2(new_n555), .A3(new_n433), .A4(KEYINPUT35), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n479), .B1(new_n547), .B2(new_n548), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n508), .A2(new_n518), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n580), .A2(new_n434), .A3(new_n339), .A4(new_n480), .ZN(new_n581));
  AOI22_X1  g380(.A1(new_n578), .A2(new_n579), .B1(new_n581), .B2(KEYINPUT35), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n270), .B1(new_n574), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n480), .ZN(new_n585));
  INV_X1    g384(.A(G92gat), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n586), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT7), .ZN(new_n588));
  INV_X1    g387(.A(G85gat), .ZN(new_n589));
  OAI21_X1  g388(.A(G92gat), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n587), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT8), .ZN(new_n593));
  NAND2_X1  g392(.A1(G99gat), .A2(G106gat), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT95), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n596), .B1(new_n595), .B2(new_n594), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(G99gat), .B(G106gat), .Z(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n599), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n601), .A2(new_n592), .A3(new_n597), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n600), .A2(KEYINPUT96), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT96), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n601), .A2(new_n592), .A3(new_n597), .A4(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n606), .A2(new_n242), .A3(new_n243), .ZN(new_n607));
  INV_X1    g406(.A(G232gat), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n608), .A2(new_n485), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(KEYINPUT41), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT97), .ZN(new_n612));
  AND3_X1   g411(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n240), .A2(new_n241), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n605), .B(new_n603), .C1(new_n614), .C2(new_n244), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n612), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n606), .B1(KEYINPUT17), .B2(new_n232), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n617), .A2(KEYINPUT97), .A3(new_n245), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n611), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G190gat), .B(G218gat), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(KEYINPUT98), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n609), .A2(KEYINPUT41), .ZN(new_n623));
  XNOR2_X1  g422(.A(G134gat), .B(G162gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n619), .A2(new_n621), .ZN(new_n627));
  AOI211_X1 g426(.A(new_n620), .B(new_n611), .C1(new_n616), .C2(new_n618), .ZN(new_n628));
  OAI22_X1  g427(.A1(new_n622), .A2(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n616), .A2(new_n618), .ZN(new_n630));
  INV_X1    g429(.A(new_n611), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n620), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n619), .A2(new_n621), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n633), .A2(KEYINPUT98), .A3(new_n634), .A4(new_n625), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n629), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G57gat), .B(G64gat), .ZN(new_n637));
  AOI21_X1  g436(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(G71gat), .B(G78gat), .Z(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n639), .B(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(KEYINPUT21), .ZN(new_n643));
  XNOR2_X1  g442(.A(G127gat), .B(G155gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n207), .B1(KEYINPUT21), .B2(new_n642), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n645), .B(new_n646), .Z(new_n647));
  XNOR2_X1  g446(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT94), .ZN(new_n649));
  NAND2_X1  g448(.A1(G231gat), .A2(G233gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT93), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n649), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(G183gat), .B(G211gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n647), .B(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n636), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n639), .B(new_n640), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n603), .A2(new_n605), .A3(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n642), .A2(new_n602), .A3(new_n600), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(G230gat), .A2(G233gat), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT10), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n658), .A2(new_n664), .A3(new_n659), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT99), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n658), .A2(new_n659), .A3(KEYINPUT99), .A4(new_n664), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n657), .A2(new_n664), .ZN(new_n669));
  AOI22_X1  g468(.A1(new_n667), .A2(new_n668), .B1(new_n606), .B2(new_n669), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n661), .B(KEYINPUT100), .Z(new_n671));
  OAI21_X1  g470(.A(new_n663), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(G120gat), .B(G148gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(G176gat), .B(G204gat), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n673), .B(new_n674), .Z(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n667), .A2(new_n668), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n669), .A2(new_n606), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(new_n661), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n676), .B1(new_n660), .B2(new_n662), .ZN(new_n681));
  AOI22_X1  g480(.A1(new_n672), .A2(new_n676), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n656), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n584), .A2(new_n585), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g485(.A1(new_n584), .A2(new_n684), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(new_n434), .ZN(new_n688));
  XOR2_X1   g487(.A(KEYINPUT16), .B(G8gat), .Z(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(G8gat), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n690), .B1(new_n691), .B2(new_n688), .ZN(new_n692));
  MUX2_X1   g491(.A(new_n690), .B(new_n692), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g492(.A(new_n687), .ZN(new_n694));
  OAI21_X1  g493(.A(KEYINPUT73), .B1(new_n504), .B2(new_n506), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(new_n520), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n524), .B1(new_n696), .B2(new_n507), .ZN(new_n697));
  AOI21_X1  g496(.A(KEYINPUT36), .B1(new_n521), .B2(new_n522), .ZN(new_n698));
  OAI21_X1  g497(.A(KEYINPUT102), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT102), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n519), .A2(new_n700), .A3(new_n525), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n694), .A2(G15gat), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(G15gat), .B1(new_n694), .B2(new_n523), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT101), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AOI211_X1 g506(.A(KEYINPUT101), .B(G15gat), .C1(new_n694), .C2(new_n523), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n704), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT103), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n704), .B(KEYINPUT103), .C1(new_n707), .C2(new_n708), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(G1326gat));
  NAND3_X1  g512(.A1(new_n584), .A2(new_n555), .A3(new_n684), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT43), .B(G22gat), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1327gat));
  NAND4_X1  g515(.A1(new_n584), .A2(new_n636), .A3(new_n655), .A4(new_n682), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n718), .A2(new_n222), .A3(new_n585), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT45), .ZN(new_n720));
  INV_X1    g519(.A(new_n636), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OR2_X1    g522(.A1(new_n481), .A2(new_n526), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n549), .A2(new_n571), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT87), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n549), .A2(new_n571), .A3(KEYINPUT87), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n724), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n723), .B1(new_n729), .B2(new_n582), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n655), .A2(new_n682), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n270), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n481), .B1(new_n699), .B2(new_n701), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n733), .B1(new_n572), .B2(new_n573), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n721), .B1(new_n734), .B2(new_n583), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n730), .B(new_n732), .C1(new_n735), .C2(KEYINPUT44), .ZN(new_n736));
  OAI21_X1  g535(.A(G29gat), .B1(new_n736), .B2(new_n480), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n720), .A2(new_n737), .ZN(G1328gat));
  INV_X1    g537(.A(KEYINPUT104), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(KEYINPUT46), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n718), .A2(new_n225), .A3(new_n433), .A4(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n739), .A2(KEYINPUT46), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n229), .B1(new_n736), .B2(new_n434), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(G1329gat));
  OAI21_X1  g544(.A(G43gat), .B1(new_n736), .B2(new_n702), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT105), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT47), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n718), .A2(new_n208), .A3(new_n523), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n748), .B(new_n750), .ZN(G1330gat));
  NAND2_X1  g550(.A1(new_n734), .A2(new_n583), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(new_n636), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n574), .A2(new_n583), .ZN(new_n754));
  AOI22_X1  g553(.A1(new_n753), .A2(new_n722), .B1(new_n754), .B2(new_n723), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n755), .A2(KEYINPUT106), .A3(new_n555), .A4(new_n732), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT106), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n757), .B1(new_n736), .B2(new_n339), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n756), .A2(new_n758), .A3(G50gat), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n339), .A2(G50gat), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(KEYINPUT48), .B1(new_n717), .B2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n727), .A2(new_n728), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n582), .B1(new_n765), .B2(new_n733), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n722), .B1(new_n766), .B2(new_n721), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n767), .A2(new_n555), .A3(new_n730), .A4(new_n732), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(G50gat), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n718), .A2(new_n760), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT48), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT107), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n764), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n235), .B1(new_n768), .B2(new_n757), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n762), .B1(new_n775), .B2(new_n756), .ZN(new_n776));
  OAI21_X1  g575(.A(KEYINPUT107), .B1(new_n776), .B2(new_n771), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n774), .A2(new_n777), .ZN(G1331gat));
  INV_X1    g577(.A(new_n682), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n656), .A2(new_n270), .A3(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n766), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n585), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(G57gat), .ZN(G1332gat));
  NOR3_X1   g582(.A1(new_n766), .A2(new_n434), .A3(new_n780), .ZN(new_n784));
  NOR2_X1   g583(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n785));
  AND2_X1   g584(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n787), .B1(new_n784), .B2(new_n785), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(KEYINPUT108), .ZN(G1333gat));
  INV_X1    g588(.A(G71gat), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n781), .A2(new_n790), .A3(new_n523), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n766), .A2(new_n702), .A3(new_n780), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n791), .B1(new_n792), .B2(new_n790), .ZN(new_n793));
  XNOR2_X1  g592(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n793), .B(new_n794), .ZN(G1334gat));
  NAND2_X1  g594(.A1(new_n781), .A2(new_n555), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(G78gat), .ZN(G1335gat));
  INV_X1    g596(.A(new_n655), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n798), .A2(new_n269), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n752), .A2(new_n636), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n735), .A2(KEYINPUT51), .A3(new_n799), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n802), .A2(KEYINPUT110), .A3(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT110), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n800), .A2(new_n805), .A3(new_n801), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n585), .A2(new_n589), .A3(new_n779), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(KEYINPUT111), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n269), .A2(new_n798), .A3(new_n682), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n730), .B(new_n811), .C1(new_n735), .C2(KEYINPUT44), .ZN(new_n812));
  OAI21_X1  g611(.A(G85gat), .B1(new_n812), .B2(new_n480), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n810), .A2(new_n813), .ZN(G1336gat));
  NOR3_X1   g613(.A1(new_n434), .A2(G92gat), .A3(new_n682), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n804), .A2(new_n806), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(KEYINPUT112), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT112), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n804), .A2(new_n818), .A3(new_n806), .A4(new_n815), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n767), .A2(new_n433), .A3(new_n730), .A4(new_n811), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(KEYINPUT113), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT113), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n586), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT52), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n820), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n802), .A2(new_n803), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n815), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n829), .B1(new_n822), .B2(new_n586), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(KEYINPUT52), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n827), .A2(new_n831), .ZN(G1337gat));
  INV_X1    g631(.A(G99gat), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n755), .A2(new_n703), .A3(new_n811), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT114), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n836), .B1(new_n835), .B2(new_n834), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n807), .A2(new_n833), .A3(new_n523), .A4(new_n779), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(G1338gat));
  OR3_X1    g638(.A1(new_n339), .A2(G106gat), .A3(new_n682), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n804), .A2(new_n806), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(KEYINPUT116), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n804), .A2(new_n844), .A3(new_n806), .A4(new_n841), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n767), .A2(new_n555), .A3(new_n730), .A4(new_n811), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n847), .A2(G106gat), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n848), .A2(KEYINPUT53), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  AOI22_X1  g649(.A1(new_n828), .A2(new_n841), .B1(new_n847), .B2(G106gat), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT53), .ZN(new_n852));
  OAI21_X1  g651(.A(KEYINPUT115), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n840), .B1(new_n802), .B2(new_n803), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n854), .B(KEYINPUT53), .C1(new_n848), .C2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n850), .A2(new_n857), .ZN(G1339gat));
  NOR2_X1   g657(.A1(new_n683), .A2(new_n269), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n860));
  INV_X1    g659(.A(new_n671), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n679), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(KEYINPUT54), .B1(new_n670), .B2(new_n662), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n677), .A2(new_n671), .A3(new_n678), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n862), .B(new_n676), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT55), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n269), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n670), .A2(new_n671), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n680), .A2(KEYINPUT54), .A3(new_n869), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n870), .A2(KEYINPUT55), .A3(new_n676), .A4(new_n862), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n680), .A2(new_n681), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n257), .A2(new_n258), .A3(new_n254), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n247), .B1(new_n246), .B2(new_n248), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n264), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n268), .A2(new_n876), .ZN(new_n877));
  OAI22_X1  g676(.A1(new_n868), .A2(new_n873), .B1(new_n682), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n721), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n871), .A2(new_n872), .ZN(new_n880));
  AOI22_X1  g679(.A1(new_n629), .A2(new_n635), .B1(new_n865), .B2(new_n866), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT117), .ZN(new_n882));
  INV_X1    g681(.A(new_n877), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n880), .A2(new_n881), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n880), .A2(new_n881), .A3(new_n883), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(KEYINPUT117), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n879), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n859), .B1(new_n887), .B2(new_n655), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n888), .A2(new_n480), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n580), .A2(new_n339), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n890), .A2(new_n433), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(G113gat), .B1(new_n893), .B2(new_n269), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n888), .A2(new_n555), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n480), .A2(new_n433), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n895), .A2(new_n523), .A3(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(G113gat), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n897), .A2(new_n898), .A3(new_n270), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n894), .A2(new_n899), .ZN(G1340gat));
  OAI21_X1  g699(.A(G120gat), .B1(new_n897), .B2(new_n682), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(KEYINPUT118), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n682), .A2(G120gat), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n902), .B1(new_n892), .B2(new_n903), .ZN(G1341gat));
  OR3_X1    g703(.A1(new_n892), .A2(G127gat), .A3(new_n655), .ZN(new_n905));
  OAI21_X1  g704(.A(G127gat), .B1(new_n897), .B2(new_n655), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(G1342gat));
  OR3_X1    g706(.A1(new_n892), .A2(G134gat), .A3(new_n721), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n908), .A2(KEYINPUT56), .ZN(new_n909));
  OAI21_X1  g708(.A(G134gat), .B1(new_n897), .B2(new_n721), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(KEYINPUT56), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(G1343gat));
  NOR3_X1   g711(.A1(new_n703), .A2(new_n433), .A3(new_n339), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n889), .A2(new_n913), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n914), .A2(G141gat), .A3(new_n270), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n915), .A2(KEYINPUT58), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT57), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n917), .B1(new_n888), .B2(new_n339), .ZN(new_n918));
  AOI22_X1  g717(.A1(new_n878), .A2(new_n721), .B1(new_n885), .B2(KEYINPUT117), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n798), .B1(new_n919), .B2(new_n884), .ZN(new_n920));
  OAI211_X1 g719(.A(KEYINPUT57), .B(new_n555), .C1(new_n920), .C2(new_n859), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n702), .A2(new_n896), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(G141gat), .B1(new_n925), .B2(new_n270), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n916), .A2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT119), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n922), .A2(KEYINPUT119), .A3(new_n924), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n929), .A2(new_n269), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n915), .B1(new_n931), .B2(G141gat), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT58), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n927), .B1(new_n932), .B2(new_n933), .ZN(G1344gat));
  INV_X1    g733(.A(new_n914), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(new_n276), .A3(new_n779), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n936), .B(KEYINPUT120), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT59), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n924), .A2(new_n779), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n636), .A2(new_n872), .A3(new_n871), .A4(new_n867), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n883), .B1(new_n940), .B2(KEYINPUT121), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT121), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n942), .B1(new_n880), .B2(new_n881), .ZN(new_n943));
  AOI22_X1  g742(.A1(new_n267), .A2(new_n268), .B1(new_n865), .B2(new_n866), .ZN(new_n944));
  AOI22_X1  g743(.A1(new_n880), .A2(new_n944), .B1(new_n779), .B2(new_n883), .ZN(new_n945));
  OAI22_X1  g744(.A1(new_n941), .A2(new_n943), .B1(new_n945), .B2(new_n636), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT122), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n798), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  OAI211_X1 g747(.A(new_n879), .B(KEYINPUT122), .C1(new_n943), .C2(new_n941), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n859), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n917), .B1(new_n950), .B2(new_n339), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n939), .B1(new_n951), .B2(new_n921), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n276), .B1(new_n952), .B2(KEYINPUT123), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT123), .ZN(new_n954));
  INV_X1    g753(.A(new_n921), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n946), .A2(new_n947), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n956), .A2(new_n655), .A3(new_n949), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n555), .B1(new_n957), .B2(new_n859), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n955), .B1(new_n958), .B2(new_n917), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n954), .B1(new_n959), .B2(new_n939), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n938), .B1(new_n953), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n938), .A2(G148gat), .ZN(new_n962));
  AOI21_X1  g761(.A(KEYINPUT119), .B1(new_n922), .B2(new_n924), .ZN(new_n963));
  AOI211_X1 g762(.A(new_n928), .B(new_n923), .C1(new_n918), .C2(new_n921), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n962), .B1(new_n965), .B2(new_n779), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n937), .B1(new_n961), .B2(new_n966), .ZN(G1345gat));
  NAND3_X1  g766(.A1(new_n935), .A2(new_n271), .A3(new_n798), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n963), .A2(new_n964), .A3(new_n655), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n968), .B1(new_n969), .B2(new_n271), .ZN(G1346gat));
  NOR2_X1   g769(.A1(new_n721), .A2(new_n272), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n965), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g771(.A(G162gat), .B1(new_n935), .B2(new_n636), .ZN(new_n973));
  INV_X1    g772(.A(new_n973), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n972), .A2(KEYINPUT124), .A3(new_n974), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT124), .ZN(new_n976));
  INV_X1    g775(.A(new_n971), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n963), .A2(new_n964), .A3(new_n977), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n976), .B1(new_n978), .B2(new_n973), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n975), .A2(new_n979), .ZN(G1347gat));
  NOR2_X1   g779(.A1(new_n585), .A2(new_n434), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(new_n523), .ZN(new_n982));
  XOR2_X1   g781(.A(new_n982), .B(KEYINPUT125), .Z(new_n983));
  NAND2_X1  g782(.A1(new_n895), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g783(.A(G169gat), .B1(new_n984), .B2(new_n270), .ZN(new_n985));
  INV_X1    g784(.A(new_n981), .ZN(new_n986));
  NOR3_X1   g785(.A1(new_n888), .A2(new_n890), .A3(new_n986), .ZN(new_n987));
  NAND4_X1  g786(.A1(new_n987), .A2(new_n269), .A3(new_n392), .A4(new_n394), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n985), .A2(new_n988), .ZN(G1348gat));
  OAI21_X1  g788(.A(G176gat), .B1(new_n984), .B2(new_n682), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n987), .A2(new_n372), .A3(new_n779), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n991), .ZN(G1349gat));
  OAI21_X1  g791(.A(G183gat), .B1(new_n984), .B2(new_n655), .ZN(new_n993));
  NAND4_X1  g792(.A1(new_n987), .A2(new_n357), .A3(new_n362), .A4(new_n798), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT60), .ZN(new_n995));
  AOI22_X1  g794(.A1(new_n993), .A2(new_n994), .B1(KEYINPUT126), .B2(new_n995), .ZN(new_n996));
  NOR2_X1   g795(.A1(new_n995), .A2(KEYINPUT126), .ZN(new_n997));
  XNOR2_X1  g796(.A(new_n996), .B(new_n997), .ZN(G1350gat));
  OAI21_X1  g797(.A(G190gat), .B1(new_n984), .B2(new_n721), .ZN(new_n999));
  XNOR2_X1  g798(.A(new_n999), .B(KEYINPUT61), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n987), .A2(new_n365), .A3(new_n636), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1000), .A2(new_n1001), .ZN(G1351gat));
  NOR2_X1   g801(.A1(new_n888), .A2(new_n339), .ZN(new_n1003));
  NOR2_X1   g802(.A1(new_n703), .A2(new_n986), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g804(.A(new_n1005), .ZN(new_n1006));
  AOI21_X1  g805(.A(G197gat), .B1(new_n1006), .B2(new_n269), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n951), .A2(new_n921), .ZN(new_n1008));
  AND2_X1   g807(.A1(new_n1008), .A2(new_n1004), .ZN(new_n1009));
  AND2_X1   g808(.A1(new_n269), .A2(G197gat), .ZN(new_n1010));
  AOI21_X1  g809(.A(new_n1007), .B1(new_n1009), .B2(new_n1010), .ZN(G1352gat));
  XNOR2_X1  g810(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1012));
  INV_X1    g811(.A(G204gat), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n779), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g813(.A(new_n1012), .B1(new_n1005), .B2(new_n1014), .ZN(new_n1015));
  OR3_X1    g814(.A1(new_n1005), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1016));
  AND2_X1   g815(.A1(new_n1009), .A2(new_n779), .ZN(new_n1017));
  OAI211_X1 g816(.A(new_n1015), .B(new_n1016), .C1(new_n1017), .C2(new_n1013), .ZN(G1353gat));
  NAND3_X1  g817(.A1(new_n1006), .A2(new_n299), .A3(new_n798), .ZN(new_n1019));
  NAND3_X1  g818(.A1(new_n1008), .A2(new_n798), .A3(new_n1004), .ZN(new_n1020));
  AND3_X1   g819(.A1(new_n1020), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1021));
  AOI21_X1  g820(.A(KEYINPUT63), .B1(new_n1020), .B2(G211gat), .ZN(new_n1022));
  OAI21_X1  g821(.A(new_n1019), .B1(new_n1021), .B2(new_n1022), .ZN(G1354gat));
  NAND3_X1  g822(.A1(new_n1006), .A2(new_n300), .A3(new_n636), .ZN(new_n1024));
  AND2_X1   g823(.A1(new_n1009), .A2(new_n636), .ZN(new_n1025));
  OAI21_X1  g824(.A(new_n1024), .B1(new_n1025), .B2(new_n300), .ZN(G1355gat));
endmodule


