

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589;

  XNOR2_X1 U322 ( .A(n301), .B(n300), .ZN(n306) );
  XNOR2_X1 U323 ( .A(n299), .B(n298), .ZN(n300) );
  INV_X1 U324 ( .A(G15GAT), .ZN(n292) );
  XNOR2_X1 U325 ( .A(n293), .B(n292), .ZN(n294) );
  INV_X1 U326 ( .A(KEYINPUT33), .ZN(n434) );
  XNOR2_X1 U327 ( .A(n346), .B(n294), .ZN(n295) );
  XNOR2_X1 U328 ( .A(n435), .B(n434), .ZN(n436) );
  INV_X1 U329 ( .A(KEYINPUT37), .ZN(n414) );
  NOR2_X1 U330 ( .A1(n377), .A2(n376), .ZN(n486) );
  XNOR2_X1 U331 ( .A(n437), .B(n436), .ZN(n439) );
  XNOR2_X1 U332 ( .A(n414), .B(KEYINPUT98), .ZN(n415) );
  XNOR2_X1 U333 ( .A(n416), .B(n415), .ZN(n521) );
  NOR2_X1 U334 ( .A1(n480), .A2(n479), .ZN(n569) );
  XNOR2_X1 U335 ( .A(n444), .B(KEYINPUT38), .ZN(n506) );
  XNOR2_X1 U336 ( .A(n481), .B(G190GAT), .ZN(n482) );
  XNOR2_X1 U337 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U338 ( .A(n483), .B(n482), .ZN(G1351GAT) );
  XNOR2_X1 U339 ( .A(n448), .B(n447), .ZN(G1330GAT) );
  XOR2_X1 U340 ( .A(G127GAT), .B(KEYINPUT0), .Z(n291) );
  XNOR2_X1 U341 ( .A(G113GAT), .B(G134GAT), .ZN(n290) );
  XNOR2_X1 U342 ( .A(n291), .B(n290), .ZN(n346) );
  NAND2_X1 U343 ( .A1(G227GAT), .A2(G233GAT), .ZN(n293) );
  XOR2_X1 U344 ( .A(G120GAT), .B(G71GAT), .Z(n441) );
  XOR2_X1 U345 ( .A(n295), .B(n441), .Z(n301) );
  XOR2_X1 U346 ( .A(G176GAT), .B(KEYINPUT20), .Z(n297) );
  XNOR2_X1 U347 ( .A(G169GAT), .B(KEYINPUT77), .ZN(n296) );
  XNOR2_X1 U348 ( .A(n297), .B(n296), .ZN(n299) );
  XNOR2_X1 U349 ( .A(G43GAT), .B(G99GAT), .ZN(n298) );
  XOR2_X1 U350 ( .A(KEYINPUT76), .B(KEYINPUT19), .Z(n303) );
  XNOR2_X1 U351 ( .A(G183GAT), .B(KEYINPUT18), .ZN(n302) );
  XNOR2_X1 U352 ( .A(n303), .B(n302), .ZN(n305) );
  XOR2_X1 U353 ( .A(G190GAT), .B(KEYINPUT17), .Z(n304) );
  XNOR2_X1 U354 ( .A(n305), .B(n304), .ZN(n362) );
  XNOR2_X1 U355 ( .A(n306), .B(n362), .ZN(n479) );
  INV_X1 U356 ( .A(n479), .ZN(n535) );
  XNOR2_X1 U357 ( .A(G22GAT), .B(G197GAT), .ZN(n307) );
  XNOR2_X1 U358 ( .A(n307), .B(G141GAT), .ZN(n417) );
  XOR2_X1 U359 ( .A(KEYINPUT78), .B(n417), .Z(n309) );
  NAND2_X1 U360 ( .A1(G228GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U361 ( .A(n309), .B(n308), .ZN(n328) );
  XNOR2_X1 U362 ( .A(G211GAT), .B(KEYINPUT21), .ZN(n310) );
  XNOR2_X1 U363 ( .A(n310), .B(KEYINPUT80), .ZN(n359) );
  XOR2_X1 U364 ( .A(n359), .B(KEYINPUT79), .Z(n312) );
  XOR2_X1 U365 ( .A(G218GAT), .B(G162GAT), .Z(n391) );
  XNOR2_X1 U366 ( .A(G50GAT), .B(n391), .ZN(n311) );
  XNOR2_X1 U367 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U368 ( .A(KEYINPUT81), .B(KEYINPUT24), .Z(n314) );
  XNOR2_X1 U369 ( .A(KEYINPUT22), .B(KEYINPUT23), .ZN(n313) );
  XNOR2_X1 U370 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U371 ( .A(n316), .B(n315), .Z(n326) );
  XNOR2_X1 U372 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n317) );
  XNOR2_X1 U373 ( .A(n317), .B(KEYINPUT2), .ZN(n345) );
  XNOR2_X1 U374 ( .A(G106GAT), .B(G204GAT), .ZN(n323) );
  INV_X1 U375 ( .A(G148GAT), .ZN(n318) );
  NAND2_X1 U376 ( .A1(G78GAT), .A2(n318), .ZN(n321) );
  INV_X1 U377 ( .A(G78GAT), .ZN(n319) );
  NAND2_X1 U378 ( .A1(n319), .A2(G148GAT), .ZN(n320) );
  NAND2_X1 U379 ( .A1(n321), .A2(n320), .ZN(n322) );
  XNOR2_X1 U380 ( .A(n323), .B(n322), .ZN(n430) );
  BUF_X1 U381 ( .A(n430), .Z(n324) );
  XNOR2_X1 U382 ( .A(n345), .B(n324), .ZN(n325) );
  XNOR2_X1 U383 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U384 ( .A(n328), .B(n327), .Z(n476) );
  XNOR2_X1 U385 ( .A(n476), .B(KEYINPUT67), .ZN(n329) );
  XNOR2_X1 U386 ( .A(n329), .B(KEYINPUT28), .ZN(n538) );
  XOR2_X1 U387 ( .A(G85GAT), .B(G162GAT), .Z(n331) );
  XNOR2_X1 U388 ( .A(G29GAT), .B(G141GAT), .ZN(n330) );
  XNOR2_X1 U389 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U390 ( .A(KEYINPUT84), .B(G148GAT), .Z(n333) );
  XNOR2_X1 U391 ( .A(G1GAT), .B(G120GAT), .ZN(n332) );
  XNOR2_X1 U392 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U393 ( .A(n335), .B(n334), .Z(n340) );
  XOR2_X1 U394 ( .A(KEYINPUT82), .B(G57GAT), .Z(n337) );
  NAND2_X1 U395 ( .A1(G225GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U396 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U397 ( .A(KEYINPUT6), .B(n338), .ZN(n339) );
  XNOR2_X1 U398 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U399 ( .A(KEYINPUT1), .B(KEYINPUT5), .Z(n342) );
  XNOR2_X1 U400 ( .A(KEYINPUT83), .B(KEYINPUT4), .ZN(n341) );
  XNOR2_X1 U401 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U402 ( .A(n344), .B(n343), .Z(n348) );
  XNOR2_X1 U403 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U404 ( .A(n348), .B(n347), .ZN(n522) );
  XOR2_X1 U405 ( .A(G169GAT), .B(G8GAT), .Z(n425) );
  XOR2_X1 U406 ( .A(G218GAT), .B(G204GAT), .Z(n350) );
  XNOR2_X1 U407 ( .A(G36GAT), .B(G197GAT), .ZN(n349) );
  XNOR2_X1 U408 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U409 ( .A(n425), .B(n351), .Z(n353) );
  NAND2_X1 U410 ( .A1(G226GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U411 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U412 ( .A(KEYINPUT87), .B(KEYINPUT85), .Z(n355) );
  XNOR2_X1 U413 ( .A(KEYINPUT86), .B(KEYINPUT88), .ZN(n354) );
  XNOR2_X1 U414 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U415 ( .A(n357), .B(n356), .Z(n361) );
  XNOR2_X1 U416 ( .A(G176GAT), .B(G92GAT), .ZN(n358) );
  XNOR2_X1 U417 ( .A(n358), .B(G64GAT), .ZN(n440) );
  XNOR2_X1 U418 ( .A(n359), .B(n440), .ZN(n360) );
  XNOR2_X1 U419 ( .A(n361), .B(n360), .ZN(n363) );
  XOR2_X1 U420 ( .A(n363), .B(n362), .Z(n524) );
  XNOR2_X1 U421 ( .A(n524), .B(KEYINPUT27), .ZN(n367) );
  NAND2_X1 U422 ( .A1(n522), .A2(n367), .ZN(n533) );
  NOR2_X1 U423 ( .A1(n538), .A2(n533), .ZN(n364) );
  XNOR2_X1 U424 ( .A(n364), .B(KEYINPUT89), .ZN(n365) );
  NOR2_X1 U425 ( .A1(n535), .A2(n365), .ZN(n377) );
  NOR2_X1 U426 ( .A1(n476), .A2(n535), .ZN(n366) );
  XNOR2_X1 U427 ( .A(n366), .B(KEYINPUT26), .ZN(n571) );
  NAND2_X1 U428 ( .A1(n367), .A2(n571), .ZN(n368) );
  XOR2_X1 U429 ( .A(KEYINPUT90), .B(n368), .Z(n374) );
  INV_X1 U430 ( .A(n524), .ZN(n471) );
  NOR2_X1 U431 ( .A1(n471), .A2(n479), .ZN(n369) );
  XNOR2_X1 U432 ( .A(KEYINPUT91), .B(n369), .ZN(n370) );
  NAND2_X1 U433 ( .A1(n370), .A2(n476), .ZN(n371) );
  XNOR2_X1 U434 ( .A(n371), .B(KEYINPUT92), .ZN(n372) );
  XNOR2_X1 U435 ( .A(n372), .B(KEYINPUT25), .ZN(n373) );
  NOR2_X1 U436 ( .A1(n374), .A2(n373), .ZN(n375) );
  NOR2_X1 U437 ( .A1(n522), .A2(n375), .ZN(n376) );
  XNOR2_X1 U438 ( .A(KEYINPUT36), .B(KEYINPUT97), .ZN(n395) );
  XNOR2_X1 U439 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n378) );
  XNOR2_X1 U440 ( .A(n378), .B(G29GAT), .ZN(n379) );
  XOR2_X1 U441 ( .A(n379), .B(KEYINPUT8), .Z(n381) );
  XNOR2_X1 U442 ( .A(G43GAT), .B(G50GAT), .ZN(n380) );
  XNOR2_X1 U443 ( .A(n381), .B(n380), .ZN(n429) );
  XOR2_X1 U444 ( .A(G99GAT), .B(G85GAT), .Z(n438) );
  XOR2_X1 U445 ( .A(G92GAT), .B(n438), .Z(n383) );
  NAND2_X1 U446 ( .A1(G232GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U447 ( .A(n383), .B(n382), .ZN(n387) );
  XOR2_X1 U448 ( .A(KEYINPUT11), .B(G106GAT), .Z(n385) );
  XNOR2_X1 U449 ( .A(G190GAT), .B(G134GAT), .ZN(n384) );
  XNOR2_X1 U450 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U451 ( .A(n387), .B(n386), .Z(n393) );
  XOR2_X1 U452 ( .A(KEYINPUT10), .B(KEYINPUT72), .Z(n389) );
  XNOR2_X1 U453 ( .A(KEYINPUT9), .B(KEYINPUT71), .ZN(n388) );
  XNOR2_X1 U454 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U455 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U456 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U457 ( .A(n429), .B(n394), .ZN(n559) );
  XNOR2_X1 U458 ( .A(n395), .B(n559), .ZN(n587) );
  NOR2_X1 U459 ( .A1(n486), .A2(n587), .ZN(n413) );
  XOR2_X1 U460 ( .A(G211GAT), .B(G78GAT), .Z(n397) );
  XNOR2_X1 U461 ( .A(G22GAT), .B(G155GAT), .ZN(n396) );
  XNOR2_X1 U462 ( .A(n397), .B(n396), .ZN(n401) );
  XOR2_X1 U463 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n399) );
  XNOR2_X1 U464 ( .A(G8GAT), .B(KEYINPUT12), .ZN(n398) );
  XNOR2_X1 U465 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U466 ( .A(n401), .B(n400), .Z(n403) );
  XOR2_X1 U467 ( .A(G15GAT), .B(G1GAT), .Z(n424) );
  XOR2_X1 U468 ( .A(G57GAT), .B(KEYINPUT13), .Z(n433) );
  XNOR2_X1 U469 ( .A(n424), .B(n433), .ZN(n402) );
  XNOR2_X1 U470 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U471 ( .A(KEYINPUT73), .B(KEYINPUT75), .Z(n405) );
  NAND2_X1 U472 ( .A1(G231GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U473 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U474 ( .A(n407), .B(n406), .Z(n412) );
  XOR2_X1 U475 ( .A(G64GAT), .B(G127GAT), .Z(n409) );
  XNOR2_X1 U476 ( .A(G183GAT), .B(G71GAT), .ZN(n408) );
  XNOR2_X1 U477 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U478 ( .A(n410), .B(KEYINPUT74), .ZN(n411) );
  XOR2_X1 U479 ( .A(n412), .B(n411), .Z(n583) );
  INV_X1 U480 ( .A(n583), .ZN(n484) );
  NAND2_X1 U481 ( .A1(n413), .A2(n484), .ZN(n416) );
  XOR2_X1 U482 ( .A(n417), .B(KEYINPUT68), .Z(n419) );
  NAND2_X1 U483 ( .A1(G229GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U484 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U485 ( .A(KEYINPUT30), .B(KEYINPUT69), .Z(n421) );
  XNOR2_X1 U486 ( .A(G113GAT), .B(KEYINPUT29), .ZN(n420) );
  XNOR2_X1 U487 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U488 ( .A(n423), .B(n422), .Z(n427) );
  XNOR2_X1 U489 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U490 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U491 ( .A(n429), .B(n428), .Z(n508) );
  XOR2_X1 U492 ( .A(KEYINPUT70), .B(n508), .Z(n561) );
  XNOR2_X1 U493 ( .A(n430), .B(KEYINPUT31), .ZN(n432) );
  AND2_X1 U494 ( .A1(G230GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U495 ( .A(n432), .B(n431), .ZN(n437) );
  XNOR2_X1 U496 ( .A(n433), .B(KEYINPUT32), .ZN(n435) );
  XNOR2_X1 U497 ( .A(n439), .B(n438), .ZN(n443) );
  XOR2_X1 U498 ( .A(n441), .B(n440), .Z(n442) );
  XNOR2_X1 U499 ( .A(n443), .B(n442), .ZN(n577) );
  NAND2_X1 U500 ( .A1(n561), .A2(n577), .ZN(n489) );
  NOR2_X1 U501 ( .A1(n521), .A2(n489), .ZN(n444) );
  NAND2_X1 U502 ( .A1(n506), .A2(n535), .ZN(n448) );
  XOR2_X1 U503 ( .A(KEYINPUT40), .B(KEYINPUT101), .Z(n446) );
  XNOR2_X1 U504 ( .A(G43GAT), .B(KEYINPUT102), .ZN(n445) );
  XOR2_X1 U505 ( .A(KEYINPUT120), .B(KEYINPUT55), .Z(n478) );
  XNOR2_X1 U506 ( .A(n577), .B(KEYINPUT64), .ZN(n449) );
  XNOR2_X1 U507 ( .A(n449), .B(KEYINPUT41), .ZN(n566) );
  INV_X1 U508 ( .A(n508), .ZN(n573) );
  NAND2_X1 U509 ( .A1(n566), .A2(n573), .ZN(n452) );
  XOR2_X1 U510 ( .A(KEYINPUT46), .B(KEYINPUT110), .Z(n450) );
  XNOR2_X1 U511 ( .A(KEYINPUT109), .B(n450), .ZN(n451) );
  XNOR2_X1 U512 ( .A(n452), .B(n451), .ZN(n454) );
  NOR2_X1 U513 ( .A1(n559), .A2(n583), .ZN(n453) );
  NAND2_X1 U514 ( .A1(n454), .A2(n453), .ZN(n456) );
  INV_X1 U515 ( .A(KEYINPUT47), .ZN(n455) );
  XNOR2_X1 U516 ( .A(n456), .B(n455), .ZN(n459) );
  INV_X1 U517 ( .A(n459), .ZN(n457) );
  NAND2_X1 U518 ( .A1(n457), .A2(KEYINPUT111), .ZN(n461) );
  INV_X1 U519 ( .A(KEYINPUT111), .ZN(n458) );
  NAND2_X1 U520 ( .A1(n459), .A2(n458), .ZN(n460) );
  NAND2_X1 U521 ( .A1(n461), .A2(n460), .ZN(n468) );
  XOR2_X1 U522 ( .A(KEYINPUT112), .B(KEYINPUT45), .Z(n462) );
  XNOR2_X1 U523 ( .A(KEYINPUT66), .B(n462), .ZN(n464) );
  NOR2_X1 U524 ( .A1(n587), .A2(n484), .ZN(n463) );
  XNOR2_X1 U525 ( .A(n464), .B(n463), .ZN(n465) );
  NOR2_X1 U526 ( .A1(n561), .A2(n465), .ZN(n466) );
  NAND2_X1 U527 ( .A1(n466), .A2(n577), .ZN(n467) );
  NAND2_X1 U528 ( .A1(n468), .A2(n467), .ZN(n470) );
  XNOR2_X1 U529 ( .A(KEYINPUT113), .B(KEYINPUT48), .ZN(n469) );
  XNOR2_X1 U530 ( .A(n470), .B(n469), .ZN(n534) );
  NOR2_X1 U531 ( .A1(n471), .A2(n534), .ZN(n473) );
  INV_X1 U532 ( .A(KEYINPUT54), .ZN(n472) );
  XNOR2_X1 U533 ( .A(n473), .B(n472), .ZN(n474) );
  NOR2_X1 U534 ( .A1(n522), .A2(n474), .ZN(n475) );
  XOR2_X1 U535 ( .A(KEYINPUT65), .B(n475), .Z(n572) );
  NAND2_X1 U536 ( .A1(n572), .A2(n476), .ZN(n477) );
  XNOR2_X1 U537 ( .A(n478), .B(n477), .ZN(n480) );
  NAND2_X1 U538 ( .A1(n569), .A2(n559), .ZN(n483) );
  XOR2_X1 U539 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n481) );
  NOR2_X1 U540 ( .A1(n484), .A2(n559), .ZN(n485) );
  XNOR2_X1 U541 ( .A(n485), .B(KEYINPUT16), .ZN(n488) );
  INV_X1 U542 ( .A(n486), .ZN(n487) );
  NAND2_X1 U543 ( .A1(n488), .A2(n487), .ZN(n509) );
  NOR2_X1 U544 ( .A1(n489), .A2(n509), .ZN(n497) );
  NAND2_X1 U545 ( .A1(n497), .A2(n522), .ZN(n492) );
  XOR2_X1 U546 ( .A(G1GAT), .B(KEYINPUT34), .Z(n490) );
  XNOR2_X1 U547 ( .A(KEYINPUT93), .B(n490), .ZN(n491) );
  XNOR2_X1 U548 ( .A(n492), .B(n491), .ZN(G1324GAT) );
  NAND2_X1 U549 ( .A1(n524), .A2(n497), .ZN(n493) );
  XNOR2_X1 U550 ( .A(n493), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U551 ( .A(KEYINPUT94), .B(KEYINPUT35), .Z(n495) );
  NAND2_X1 U552 ( .A1(n497), .A2(n535), .ZN(n494) );
  XNOR2_X1 U553 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U554 ( .A(G15GAT), .B(n496), .ZN(G1326GAT) );
  XOR2_X1 U555 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n499) );
  NAND2_X1 U556 ( .A1(n497), .A2(n538), .ZN(n498) );
  XNOR2_X1 U557 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U558 ( .A(G22GAT), .B(n500), .ZN(G1327GAT) );
  NAND2_X1 U559 ( .A1(n506), .A2(n522), .ZN(n503) );
  XNOR2_X1 U560 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n501) );
  XNOR2_X1 U561 ( .A(n501), .B(KEYINPUT99), .ZN(n502) );
  XNOR2_X1 U562 ( .A(n503), .B(n502), .ZN(G1328GAT) );
  XNOR2_X1 U563 ( .A(G36GAT), .B(KEYINPUT100), .ZN(n505) );
  NAND2_X1 U564 ( .A1(n524), .A2(n506), .ZN(n504) );
  XNOR2_X1 U565 ( .A(n505), .B(n504), .ZN(G1329GAT) );
  NAND2_X1 U566 ( .A1(n506), .A2(n538), .ZN(n507) );
  XNOR2_X1 U567 ( .A(n507), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT42), .B(KEYINPUT103), .Z(n511) );
  NAND2_X1 U569 ( .A1(n508), .A2(n566), .ZN(n520) );
  NOR2_X1 U570 ( .A1(n520), .A2(n509), .ZN(n516) );
  NAND2_X1 U571 ( .A1(n516), .A2(n522), .ZN(n510) );
  XNOR2_X1 U572 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U573 ( .A(G57GAT), .B(n512), .ZN(G1332GAT) );
  NAND2_X1 U574 ( .A1(n524), .A2(n516), .ZN(n513) );
  XNOR2_X1 U575 ( .A(n513), .B(KEYINPUT104), .ZN(n514) );
  XNOR2_X1 U576 ( .A(G64GAT), .B(n514), .ZN(G1333GAT) );
  NAND2_X1 U577 ( .A1(n516), .A2(n535), .ZN(n515) );
  XNOR2_X1 U578 ( .A(n515), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT43), .B(KEYINPUT105), .Z(n518) );
  NAND2_X1 U580 ( .A1(n516), .A2(n538), .ZN(n517) );
  XNOR2_X1 U581 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U582 ( .A(G78GAT), .B(n519), .Z(G1335GAT) );
  NOR2_X1 U583 ( .A1(n521), .A2(n520), .ZN(n529) );
  NAND2_X1 U584 ( .A1(n522), .A2(n529), .ZN(n523) );
  XNOR2_X1 U585 ( .A(G85GAT), .B(n523), .ZN(G1336GAT) );
  NAND2_X1 U586 ( .A1(n524), .A2(n529), .ZN(n525) );
  XNOR2_X1 U587 ( .A(n525), .B(KEYINPUT106), .ZN(n526) );
  XNOR2_X1 U588 ( .A(G92GAT), .B(n526), .ZN(G1337GAT) );
  XOR2_X1 U589 ( .A(G99GAT), .B(KEYINPUT107), .Z(n528) );
  NAND2_X1 U590 ( .A1(n529), .A2(n535), .ZN(n527) );
  XNOR2_X1 U591 ( .A(n528), .B(n527), .ZN(G1338GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT44), .B(KEYINPUT108), .Z(n531) );
  NAND2_X1 U593 ( .A1(n529), .A2(n538), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U595 ( .A(G106GAT), .B(n532), .Z(G1339GAT) );
  NOR2_X1 U596 ( .A1(n534), .A2(n533), .ZN(n547) );
  NAND2_X1 U597 ( .A1(n535), .A2(n547), .ZN(n536) );
  XNOR2_X1 U598 ( .A(KEYINPUT114), .B(n536), .ZN(n537) );
  NOR2_X1 U599 ( .A1(n538), .A2(n537), .ZN(n544) );
  NAND2_X1 U600 ( .A1(n561), .A2(n544), .ZN(n539) );
  XNOR2_X1 U601 ( .A(G113GAT), .B(n539), .ZN(G1340GAT) );
  XOR2_X1 U602 ( .A(G120GAT), .B(KEYINPUT49), .Z(n541) );
  NAND2_X1 U603 ( .A1(n544), .A2(n566), .ZN(n540) );
  XNOR2_X1 U604 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  NAND2_X1 U605 ( .A1(n583), .A2(n544), .ZN(n542) );
  XNOR2_X1 U606 ( .A(n542), .B(KEYINPUT50), .ZN(n543) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(n543), .ZN(G1342GAT) );
  XOR2_X1 U608 ( .A(G134GAT), .B(KEYINPUT51), .Z(n546) );
  NAND2_X1 U609 ( .A1(n544), .A2(n559), .ZN(n545) );
  XNOR2_X1 U610 ( .A(n546), .B(n545), .ZN(G1343GAT) );
  XNOR2_X1 U611 ( .A(G141GAT), .B(KEYINPUT116), .ZN(n550) );
  NAND2_X1 U612 ( .A1(n571), .A2(n547), .ZN(n548) );
  XNOR2_X1 U613 ( .A(n548), .B(KEYINPUT115), .ZN(n558) );
  NAND2_X1 U614 ( .A1(n558), .A2(n573), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n550), .B(n549), .ZN(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT52), .B(KEYINPUT53), .Z(n552) );
  NAND2_X1 U617 ( .A1(n558), .A2(n566), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(n554) );
  XOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT117), .Z(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(G1345GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n556) );
  NAND2_X1 U622 ( .A1(n558), .A2(n583), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U624 ( .A(G155GAT), .B(n557), .ZN(G1346GAT) );
  NAND2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n569), .ZN(n562) );
  XNOR2_X1 U628 ( .A(G169GAT), .B(n562), .ZN(G1348GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n564) );
  XNOR2_X1 U630 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n565) );
  XOR2_X1 U632 ( .A(KEYINPUT121), .B(n565), .Z(n568) );
  NAND2_X1 U633 ( .A1(n569), .A2(n566), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1349GAT) );
  NAND2_X1 U635 ( .A1(n583), .A2(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n575) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n586) );
  INV_X1 U639 ( .A(n586), .ZN(n582) );
  NAND2_X1 U640 ( .A1(n582), .A2(n573), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(n576), .ZN(G1352GAT) );
  NOR2_X1 U643 ( .A1(n586), .A2(n577), .ZN(n581) );
  XOR2_X1 U644 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n579) );
  XNOR2_X1 U645 ( .A(G204GAT), .B(KEYINPUT125), .ZN(n578) );
  XNOR2_X1 U646 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(G1353GAT) );
  NAND2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n584), .B(KEYINPUT126), .ZN(n585) );
  XNOR2_X1 U650 ( .A(G211GAT), .B(n585), .ZN(G1354GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U652 ( .A(KEYINPUT62), .B(n588), .Z(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

