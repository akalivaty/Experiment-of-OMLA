//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 0 1 0 1 1 1 1 1 1 1 0 0 0 1 0 1 0 1 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n547, new_n548, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n606, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1150, new_n1151, new_n1152, new_n1153, new_n1155,
    new_n1156;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT65), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT67), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  OAI21_X1  g036(.A(KEYINPUT69), .B1(new_n461), .B2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n461), .A2(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n462), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT68), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  AND3_X1   g048(.A1(new_n468), .A2(G137), .A3(new_n473), .ZN(new_n474));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G125), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n473), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n464), .A2(G2105), .ZN(new_n479));
  AND2_X1   g054(.A1(new_n479), .A2(G101), .ZN(new_n480));
  NOR3_X1   g055(.A1(new_n474), .A2(new_n478), .A3(new_n480), .ZN(G160));
  NOR2_X1   g056(.A1(new_n467), .A2(new_n473), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n464), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI221_X1 g061(.A(new_n486), .B1(new_n485), .B2(new_n484), .C1(new_n473), .C2(G112), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n467), .A2(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G136), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n493), .B1(new_n494), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  AND2_X1   g071(.A1(G126), .A2(G2105), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n462), .A2(new_n465), .A3(new_n466), .A4(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT71), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n498), .A2(new_n499), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n496), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n470), .A2(new_n472), .A3(G138), .ZN(new_n503));
  OR3_X1    g078(.A1(new_n467), .A2(new_n503), .A3(KEYINPUT72), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT72), .B1(new_n467), .B2(new_n503), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n504), .A2(KEYINPUT4), .A3(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n473), .A2(new_n475), .A3(new_n507), .A4(G138), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n502), .B1(new_n506), .B2(new_n508), .ZN(G164));
  NAND2_X1  g084(.A1(KEYINPUT73), .A2(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(KEYINPUT73), .A2(KEYINPUT5), .A3(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT6), .B(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(G543), .ZN(new_n521));
  INV_X1    g096(.A(G50), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n517), .A2(new_n523), .ZN(G166));
  NAND3_X1  g099(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  INV_X1    g102(.A(G51), .ZN(new_n528));
  OAI211_X1 g103(.A(new_n525), .B(new_n527), .C1(new_n521), .C2(new_n528), .ZN(new_n529));
  AND3_X1   g104(.A1(new_n514), .A2(G89), .A3(new_n518), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(G168));
  AOI22_X1  g106(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n516), .ZN(new_n533));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  INV_X1    g109(.A(G52), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n519), .A2(new_n534), .B1(new_n521), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n533), .A2(new_n536), .ZN(G171));
  INV_X1    g112(.A(new_n519), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G81), .ZN(new_n539));
  INV_X1    g114(.A(new_n521), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G43), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  OAI211_X1 g117(.A(new_n539), .B(new_n541), .C1(new_n516), .C2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  NAND4_X1  g120(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(G188));
  INV_X1    g124(.A(G91), .ZN(new_n550));
  OR3_X1    g125(.A1(new_n519), .A2(KEYINPUT75), .A3(new_n550), .ZN(new_n551));
  OAI21_X1  g126(.A(KEYINPUT75), .B1(new_n519), .B2(new_n550), .ZN(new_n552));
  NAND2_X1  g127(.A1(KEYINPUT74), .A2(KEYINPUT9), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n540), .A2(G53), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(G53), .ZN(new_n555));
  OAI211_X1 g130(.A(KEYINPUT74), .B(KEYINPUT9), .C1(new_n521), .C2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n551), .A2(new_n552), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(G65), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n558), .B1(new_n512), .B2(new_n513), .ZN(new_n559));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  OR3_X1    g136(.A1(new_n559), .A2(KEYINPUT76), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT76), .B1(new_n559), .B2(new_n561), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n562), .A2(G651), .A3(new_n563), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n564), .A2(KEYINPUT77), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT77), .ZN(new_n566));
  AND2_X1   g141(.A1(new_n563), .A2(G651), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n566), .B1(new_n567), .B2(new_n562), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n557), .B1(new_n565), .B2(new_n568), .ZN(G299));
  INV_X1    g144(.A(G171), .ZN(G301));
  INV_X1    g145(.A(G168), .ZN(G286));
  INV_X1    g146(.A(G166), .ZN(G303));
  AOI22_X1  g147(.A1(new_n538), .A2(G87), .B1(new_n540), .B2(G49), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(G288));
  AOI22_X1  g150(.A1(new_n514), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n576));
  OR2_X1    g151(.A1(new_n576), .A2(new_n516), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n540), .A2(G48), .ZN(new_n578));
  AND2_X1   g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n538), .A2(G86), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(G305));
  AOI22_X1  g156(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n516), .ZN(new_n583));
  INV_X1    g158(.A(G85), .ZN(new_n584));
  INV_X1    g159(.A(G47), .ZN(new_n585));
  OAI22_X1  g160(.A1(new_n519), .A2(new_n584), .B1(new_n521), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  AND3_X1   g164(.A1(new_n514), .A2(G92), .A3(new_n518), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT10), .ZN(new_n591));
  INV_X1    g166(.A(G54), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n592), .B1(new_n521), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n594), .B1(new_n593), .B2(new_n521), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n514), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n596), .A2(new_n516), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n591), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n589), .B1(new_n599), .B2(G868), .ZN(G284));
  OAI21_X1  g175(.A(new_n589), .B1(new_n599), .B2(G868), .ZN(G321));
  NAND2_X1  g176(.A1(G286), .A2(G868), .ZN(new_n602));
  INV_X1    g177(.A(G299), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(G868), .ZN(G297));
  OAI21_X1  g179(.A(new_n602), .B1(new_n603), .B2(G868), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n599), .B1(new_n606), .B2(G860), .ZN(G148));
  OR3_X1    g182(.A1(new_n598), .A2(KEYINPUT79), .A3(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(KEYINPUT79), .B1(new_n598), .B2(G559), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n608), .A2(G868), .A3(new_n609), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n543), .A2(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g187(.A(KEYINPUT80), .B(KEYINPUT11), .Z(new_n613));
  XNOR2_X1  g188(.A(new_n612), .B(new_n613), .ZN(G282));
  INV_X1    g189(.A(new_n612), .ZN(G323));
  NAND2_X1  g190(.A1(new_n475), .A2(new_n479), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT12), .Z(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT13), .Z(new_n618));
  INV_X1    g193(.A(G2100), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT81), .Z(new_n621));
  NAND2_X1  g196(.A1(new_n482), .A2(G123), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n489), .A2(G135), .ZN(new_n623));
  OAI221_X1 g198(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n473), .C2(G111), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(G2096), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n618), .A2(new_n619), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT82), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n621), .A2(new_n627), .A3(new_n629), .ZN(G156));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2435), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2427), .B(G2430), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(KEYINPUT14), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT83), .Z(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(new_n632), .B2(new_n633), .ZN(new_n637));
  XOR2_X1   g212(.A(G2443), .B(G2446), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2451), .B(G2454), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT16), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n639), .A2(new_n642), .ZN(new_n644));
  XNOR2_X1  g219(.A(G1341), .B(G1348), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n643), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT84), .ZN(new_n648));
  INV_X1    g223(.A(G14), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n643), .A2(new_n644), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n649), .B1(new_n650), .B2(new_n645), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(G401));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT85), .Z(new_n656));
  XOR2_X1   g231(.A(G2072), .B(G2078), .Z(new_n657));
  AOI21_X1  g232(.A(new_n654), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n658), .A2(KEYINPUT86), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(KEYINPUT86), .ZN(new_n660));
  XOR2_X1   g235(.A(KEYINPUT87), .B(KEYINPUT17), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n657), .B(new_n661), .ZN(new_n662));
  OAI211_X1 g237(.A(new_n659), .B(new_n660), .C1(new_n656), .C2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n657), .ZN(new_n664));
  AND3_X1   g239(.A1(new_n664), .A2(new_n654), .A3(new_n655), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n665), .A2(KEYINPUT18), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(KEYINPUT18), .ZN(new_n667));
  AND2_X1   g242(.A1(new_n656), .A2(new_n654), .ZN(new_n668));
  AOI22_X1  g243(.A1(new_n666), .A2(new_n667), .B1(new_n668), .B2(new_n662), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n663), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(new_n626), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT88), .B(G2100), .ZN(new_n672));
  AND2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(G227));
  XOR2_X1   g250(.A(G1971), .B(G1976), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT19), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1956), .B(G2474), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1961), .B(G1966), .ZN(new_n679));
  AND2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n678), .A2(new_n679), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n677), .A2(new_n682), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n685));
  OAI221_X1 g260(.A(new_n681), .B1(new_n683), .B2(new_n677), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(new_n684), .B2(new_n685), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1981), .B(G1986), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n691), .B(new_n692), .Z(G229));
  INV_X1    g268(.A(KEYINPUT36), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n694), .A2(KEYINPUT93), .ZN(new_n695));
  MUX2_X1   g270(.A(G6), .B(G305), .S(G16), .Z(new_n696));
  XOR2_X1   g271(.A(KEYINPUT32), .B(G1981), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G22), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G166), .B2(new_n699), .ZN(new_n701));
  INV_X1    g276(.A(G1971), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n699), .A2(G23), .ZN(new_n704));
  INV_X1    g279(.A(G288), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n704), .B1(new_n705), .B2(new_n699), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT33), .B(G1976), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n698), .A2(new_n703), .A3(new_n708), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n709), .A2(KEYINPUT34), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(KEYINPUT34), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n712), .A2(KEYINPUT90), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(KEYINPUT90), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G25), .ZN(new_n717));
  OAI221_X1 g292(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n473), .C2(G107), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n718), .A2(KEYINPUT91), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(KEYINPUT91), .ZN(new_n720));
  AOI22_X1  g295(.A1(new_n719), .A2(new_n720), .B1(G119), .B2(new_n482), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n489), .A2(G131), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n717), .B1(new_n724), .B2(new_n716), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT35), .B(G1991), .Z(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n725), .A2(new_n727), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n699), .A2(G24), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n587), .B2(new_n699), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1986), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n710), .A2(new_n711), .A3(new_n728), .A4(new_n733), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n694), .A2(KEYINPUT92), .ZN(new_n735));
  AOI211_X1 g310(.A(new_n695), .B(new_n734), .C1(KEYINPUT93), .C2(new_n735), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n734), .A2(new_n735), .ZN(new_n737));
  INV_X1    g312(.A(G19), .ZN(new_n738));
  OR3_X1    g313(.A1(new_n738), .A2(KEYINPUT94), .A3(G16), .ZN(new_n739));
  OAI21_X1  g314(.A(KEYINPUT94), .B1(new_n738), .B2(G16), .ZN(new_n740));
  OAI211_X1 g315(.A(new_n739), .B(new_n740), .C1(new_n544), .C2(new_n699), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT95), .B(G1341), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(G168), .A2(new_n699), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n699), .B2(G21), .ZN(new_n745));
  INV_X1    g320(.A(G1966), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT31), .B(G11), .Z(new_n748));
  INV_X1    g323(.A(G28), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n749), .A2(KEYINPUT30), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT100), .ZN(new_n751));
  AOI21_X1  g326(.A(G29), .B1(new_n749), .B2(KEYINPUT30), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n748), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n747), .B(new_n753), .C1(new_n625), .C2(new_n716), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT24), .B(G34), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n716), .A2(new_n755), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT98), .Z(new_n757));
  INV_X1    g332(.A(G160), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n757), .B1(new_n758), .B2(new_n712), .ZN(new_n759));
  INV_X1    g334(.A(G2084), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(G171), .A2(new_n699), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G5), .B2(new_n699), .ZN(new_n763));
  INV_X1    g338(.A(G1961), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OAI22_X1  g340(.A1(new_n746), .A2(new_n745), .B1(new_n763), .B2(new_n764), .ZN(new_n766));
  NOR4_X1   g341(.A1(new_n754), .A2(new_n761), .A3(new_n765), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n599), .A2(G16), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G4), .B2(G16), .ZN(new_n769));
  INV_X1    g344(.A(G1348), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n716), .A2(G35), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT102), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n491), .B2(new_n715), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT29), .B(G2090), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  AND4_X1   g351(.A1(new_n743), .A2(new_n767), .A3(new_n771), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n699), .A2(G20), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT23), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n603), .B2(new_n699), .ZN(new_n780));
  INV_X1    g355(.A(G1956), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n712), .A2(G33), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n475), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n784), .A2(new_n473), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT97), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n489), .A2(G139), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT25), .Z(new_n789));
  NAND3_X1  g364(.A1(new_n786), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n783), .B1(new_n790), .B2(G29), .ZN(new_n791));
  INV_X1    g366(.A(G2072), .ZN(new_n792));
  OAI22_X1  g367(.A1(new_n769), .A2(new_n770), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n792), .B2(new_n791), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n715), .A2(G27), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G164), .B2(new_n715), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT101), .B(G2078), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n796), .B(new_n797), .Z(new_n798));
  AND2_X1   g373(.A1(new_n712), .A2(G32), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n489), .A2(G141), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT99), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n482), .A2(G129), .ZN(new_n802));
  NAND3_X1  g377(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT26), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n479), .A2(G105), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n801), .A2(new_n802), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n799), .B1(new_n806), .B2(G29), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT27), .B(G1996), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n716), .A2(G26), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT96), .B(KEYINPUT28), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n482), .A2(G128), .ZN(new_n813));
  OAI221_X1 g388(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n473), .C2(G116), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(G140), .B2(new_n489), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n812), .B1(new_n816), .B2(new_n712), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(G2067), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n807), .A2(new_n808), .ZN(new_n819));
  NOR4_X1   g394(.A1(new_n798), .A2(new_n809), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n777), .A2(new_n782), .A3(new_n794), .A4(new_n820), .ZN(new_n821));
  NOR3_X1   g396(.A1(new_n736), .A2(new_n737), .A3(new_n821), .ZN(G311));
  INV_X1    g397(.A(G311), .ZN(G150));
  AOI22_X1  g398(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n824), .A2(new_n516), .ZN(new_n825));
  INV_X1    g400(.A(G93), .ZN(new_n826));
  INV_X1    g401(.A(G55), .ZN(new_n827));
  OAI22_X1  g402(.A1(new_n519), .A2(new_n826), .B1(new_n827), .B2(new_n521), .ZN(new_n828));
  OR3_X1    g403(.A1(new_n825), .A2(new_n828), .A3(KEYINPUT103), .ZN(new_n829));
  OAI21_X1  g404(.A(KEYINPUT103), .B1(new_n825), .B2(new_n828), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n544), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NOR3_X1   g406(.A1(new_n543), .A2(new_n825), .A3(new_n828), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT38), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n599), .A2(G559), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n836), .A2(KEYINPUT39), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n836), .A2(KEYINPUT39), .ZN(new_n838));
  NOR3_X1   g413(.A1(new_n837), .A2(new_n838), .A3(G860), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n829), .A2(new_n830), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(G860), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT37), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n839), .A2(new_n842), .ZN(G145));
  NAND2_X1  g418(.A1(new_n482), .A2(G130), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n489), .A2(G142), .ZN(new_n845));
  OAI221_X1 g420(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n473), .C2(G118), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n723), .A2(new_n617), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n723), .A2(new_n617), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n847), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n850), .ZN(new_n852));
  INV_X1    g427(.A(new_n847), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n852), .A2(new_n853), .A3(new_n848), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT104), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(KEYINPUT104), .B1(new_n851), .B2(new_n854), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n860));
  NOR3_X1   g435(.A1(new_n467), .A2(new_n503), .A3(KEYINPUT72), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n508), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n501), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n498), .A2(new_n499), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n495), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n816), .B(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n806), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n790), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n859), .B(new_n869), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n491), .B(new_n625), .Z(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(G160), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n859), .A2(new_n869), .ZN(new_n874));
  INV_X1    g449(.A(new_n872), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n874), .B(new_n875), .C1(new_n869), .C2(new_n855), .ZN(new_n876));
  XOR2_X1   g451(.A(KEYINPUT105), .B(G37), .Z(new_n877));
  NAND3_X1  g452(.A1(new_n873), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g454(.A(new_n564), .B(KEYINPUT77), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n880), .A2(new_n557), .A3(new_n598), .ZN(new_n881));
  NAND2_X1  g456(.A1(G299), .A2(new_n599), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT41), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n881), .A2(new_n882), .A3(KEYINPUT106), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT106), .ZN(new_n886));
  NAND3_X1  g461(.A1(G299), .A2(new_n886), .A3(new_n599), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n884), .B1(new_n888), .B2(new_n883), .ZN(new_n889));
  INV_X1    g464(.A(new_n833), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n608), .A2(new_n609), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n890), .B(new_n891), .ZN(new_n892));
  MUX2_X1   g467(.A(new_n889), .B(new_n888), .S(new_n892), .Z(new_n893));
  OR2_X1    g468(.A1(new_n893), .A2(KEYINPUT42), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(KEYINPUT42), .ZN(new_n895));
  XNOR2_X1  g470(.A(G305), .B(new_n587), .ZN(new_n896));
  XNOR2_X1  g471(.A(G288), .B(G166), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n896), .B(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n894), .A2(new_n895), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n899), .B1(new_n894), .B2(new_n895), .ZN(new_n901));
  OAI21_X1  g476(.A(G868), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n840), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n902), .B1(G868), .B2(new_n903), .ZN(G295));
  OAI21_X1  g479(.A(new_n902), .B1(G868), .B2(new_n903), .ZN(G331));
  INV_X1    g480(.A(new_n888), .ZN(new_n906));
  XNOR2_X1  g481(.A(G168), .B(G171), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n840), .A2(new_n543), .ZN(new_n909));
  INV_X1    g484(.A(new_n832), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(KEYINPUT109), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT109), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n833), .A2(new_n913), .A3(new_n908), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n907), .B1(new_n831), .B2(new_n832), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT108), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n916), .A2(new_n917), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n906), .A2(new_n915), .A3(new_n918), .A4(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n911), .A2(new_n916), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n884), .B(new_n921), .C1(new_n888), .C2(new_n883), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n898), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  OR3_X1    g498(.A1(new_n923), .A2(KEYINPUT110), .A3(G37), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT110), .B1(new_n923), .B2(G37), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT43), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n920), .A2(new_n898), .A3(new_n922), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n924), .A2(new_n925), .A3(new_n926), .A4(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT111), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n913), .B1(new_n833), .B2(new_n908), .ZN(new_n931));
  NOR4_X1   g506(.A1(new_n831), .A2(new_n907), .A3(KEYINPUT109), .A4(new_n832), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n919), .B(new_n918), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n881), .A2(new_n882), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(KEYINPUT41), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n888), .B1(new_n936), .B2(new_n921), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n883), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n899), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n927), .A2(new_n877), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n930), .B1(new_n941), .B2(KEYINPUT43), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n929), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n928), .A2(KEYINPUT111), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n939), .A2(new_n940), .A3(new_n926), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n924), .A2(new_n927), .A3(new_n925), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n945), .B1(KEYINPUT43), .B2(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n948));
  OAI22_X1  g523(.A1(new_n943), .A2(new_n944), .B1(new_n947), .B2(new_n948), .ZN(G397));
  INV_X1    g524(.A(G2067), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n816), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n806), .B(G1996), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n816), .B(new_n950), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n724), .A2(new_n726), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n951), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(G1384), .ZN(new_n958));
  AOI21_X1  g533(.A(KEYINPUT45), .B1(new_n866), .B2(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(KEYINPUT112), .B(G40), .ZN(new_n960));
  NOR4_X1   g535(.A1(new_n474), .A2(new_n478), .A3(new_n480), .A4(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n957), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT47), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT46), .ZN(new_n966));
  OR3_X1    g541(.A1(new_n962), .A2(new_n966), .A3(G1996), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n963), .B1(new_n953), .B2(new_n806), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n966), .B1(new_n962), .B2(G1996), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n723), .A2(new_n727), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n954), .A2(new_n956), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n963), .ZN(new_n973));
  XOR2_X1   g548(.A(new_n973), .B(KEYINPUT126), .Z(new_n974));
  INV_X1    g549(.A(G1986), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n587), .A2(new_n975), .ZN(new_n976));
  XOR2_X1   g551(.A(new_n976), .B(KEYINPUT113), .Z(new_n977));
  NOR2_X1   g552(.A1(new_n977), .A2(new_n962), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n978), .B(KEYINPUT48), .ZN(new_n979));
  OAI221_X1 g554(.A(new_n964), .B1(new_n965), .B2(new_n970), .C1(new_n974), .C2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n980), .B1(new_n965), .B2(new_n970), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n982));
  AOI21_X1  g557(.A(G1384), .B1(new_n862), .B2(new_n865), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT50), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n982), .A2(new_n985), .A3(new_n961), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n764), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT45), .ZN(new_n988));
  AOI211_X1 g563(.A(new_n988), .B(G1384), .C1(new_n862), .C2(new_n865), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n959), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G2078), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n990), .A2(KEYINPUT53), .A3(new_n991), .A4(new_n961), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n988), .B1(G164), .B2(G1384), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n866), .A2(KEYINPUT45), .A3(new_n958), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n993), .A2(new_n961), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT115), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n993), .A2(KEYINPUT115), .A3(new_n994), .A4(new_n961), .ZN(new_n998));
  AOI21_X1  g573(.A(G2078), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n987), .B(new_n992), .C1(new_n999), .C2(KEYINPUT53), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(G171), .ZN(new_n1001));
  XNOR2_X1  g576(.A(KEYINPUT116), .B(G8), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n995), .A2(new_n746), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n982), .A2(new_n985), .A3(new_n760), .A4(new_n961), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1002), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(G168), .A2(new_n1002), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1006), .A2(KEYINPUT51), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1010), .B1(new_n1005), .B2(G286), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1006), .ZN(new_n1012));
  INV_X1    g587(.A(new_n986), .ZN(new_n1013));
  AOI22_X1  g588(.A1(new_n1013), .A2(new_n760), .B1(new_n995), .B2(new_n746), .ZN(new_n1014));
  INV_X1    g589(.A(G8), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1012), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1009), .B1(new_n1011), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1001), .B1(new_n1017), .B2(KEYINPUT62), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT125), .ZN(new_n1019));
  INV_X1    g594(.A(G1981), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n579), .A2(new_n1020), .A3(new_n580), .ZN(new_n1021));
  XOR2_X1   g596(.A(KEYINPUT117), .B(G86), .Z(new_n1022));
  NAND2_X1  g597(.A1(new_n538), .A2(new_n1022), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n577), .A2(new_n578), .A3(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1021), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT49), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1002), .B1(new_n983), .B2(new_n961), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1021), .B(KEYINPUT49), .C1(new_n1020), .C2(new_n1024), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n705), .A2(G1976), .ZN(new_n1031));
  INV_X1    g606(.A(G1976), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT52), .B1(G288), .B2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1028), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1030), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT52), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1035), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n997), .A2(new_n702), .A3(new_n998), .ZN(new_n1040));
  OR2_X1    g615(.A1(new_n986), .A2(G2090), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1002), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(G303), .A2(G8), .ZN(new_n1043));
  XNOR2_X1  g618(.A(new_n1043), .B(KEYINPUT55), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1039), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1046));
  AOI211_X1 g621(.A(new_n1015), .B(new_n1044), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1019), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1002), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n1044), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1049), .A2(G8), .A3(new_n1045), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1052), .A2(KEYINPUT125), .A3(new_n1053), .A4(new_n1039), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1007), .B1(new_n1014), .B2(new_n1002), .ZN(new_n1055));
  AOI21_X1  g630(.A(G1966), .B1(new_n990), .B2(new_n961), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1004), .ZN(new_n1057));
  OAI211_X1 g632(.A(G286), .B(new_n1050), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT51), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1006), .B1(new_n1060), .B2(G8), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1055), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT62), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1018), .A2(new_n1048), .A3(new_n1054), .A4(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1049), .A2(G8), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n1044), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT118), .B1(new_n1035), .B2(new_n1038), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1030), .A2(new_n1037), .A3(new_n1069), .A4(new_n1034), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n1005), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1067), .A2(new_n1071), .A3(new_n1053), .A4(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1005), .A2(G168), .ZN(new_n1074));
  NOR3_X1   g649(.A1(new_n1046), .A2(new_n1047), .A3(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g650(.A(KEYINPUT119), .B(KEYINPUT63), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1073), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1030), .A2(new_n1032), .A3(new_n705), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n1021), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1071), .A2(new_n1047), .B1(new_n1028), .B2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1065), .A2(new_n1077), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT61), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT120), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n1086));
  NAND3_X1  g661(.A1(G299), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n880), .A2(new_n1083), .A3(new_n1084), .A4(new_n557), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  XNOR2_X1  g664(.A(KEYINPUT56), .B(G2072), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n990), .A2(new_n961), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n986), .A2(new_n781), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1089), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1089), .B1(new_n1092), .B2(new_n1091), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1082), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n983), .A2(new_n961), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT121), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n983), .A2(KEYINPUT121), .A3(new_n961), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT58), .B(G1341), .Z(new_n1101));
  NAND3_X1  g676(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(G1996), .B2(new_n995), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(new_n544), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1104), .A2(KEYINPUT59), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1104), .A2(KEYINPUT59), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1096), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1089), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT122), .ZN(new_n1110));
  AND3_X1   g685(.A1(new_n1108), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1110), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1093), .A2(KEYINPUT61), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n1111), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT123), .B1(new_n1107), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1112), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1095), .A2(new_n1110), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1116), .A2(new_n1117), .A3(KEYINPUT61), .A4(new_n1093), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1104), .B(KEYINPUT59), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT123), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .A4(new_n1096), .ZN(new_n1121));
  AOI21_X1  g696(.A(G2067), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1122), .B1(new_n770), .B2(new_n986), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1123), .A2(KEYINPUT60), .A3(new_n598), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n598), .B1(new_n1123), .B2(KEYINPUT60), .ZN(new_n1125));
  OAI22_X1  g700(.A1(new_n1124), .A2(new_n1125), .B1(KEYINPUT60), .B2(new_n1123), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1115), .A2(new_n1121), .A3(new_n1126), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1116), .B(new_n1117), .C1(new_n598), .C2(new_n1123), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n1093), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1048), .A2(new_n1054), .ZN(new_n1131));
  AND2_X1   g706(.A1(KEYINPUT124), .A2(G2078), .ZN(new_n1132));
  NOR2_X1   g707(.A1(KEYINPUT124), .A2(G2078), .ZN(new_n1133));
  OAI211_X1 g708(.A(KEYINPUT53), .B(G40), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n758), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n990), .A2(new_n1135), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n987), .B(new_n1136), .C1(new_n999), .C2(KEYINPUT53), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1137), .A2(G171), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT54), .B1(new_n1000), .B2(G171), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1017), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  OR2_X1    g715(.A1(new_n1137), .A2(G171), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT54), .B1(new_n1141), .B2(new_n1001), .ZN(new_n1142));
  NOR3_X1   g717(.A1(new_n1131), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1081), .B1(new_n1130), .B2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n977), .B1(new_n975), .B2(new_n587), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n963), .B1(new_n972), .B2(new_n1145), .ZN(new_n1146));
  XOR2_X1   g721(.A(new_n1146), .B(KEYINPUT114), .Z(new_n1147));
  OAI21_X1  g722(.A(new_n981), .B1(new_n1144), .B2(new_n1147), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g723(.A(G229), .B1(new_n648), .B2(new_n651), .ZN(new_n1150));
  OAI21_X1  g724(.A(G319), .B1(new_n673), .B2(new_n674), .ZN(new_n1151));
  XNOR2_X1  g725(.A(new_n1151), .B(KEYINPUT127), .ZN(new_n1152));
  NAND3_X1  g726(.A1(new_n878), .A2(new_n1150), .A3(new_n1152), .ZN(new_n1153));
  NOR2_X1   g727(.A1(new_n1153), .A2(new_n947), .ZN(G308));
  NAND2_X1  g728(.A1(new_n946), .A2(KEYINPUT43), .ZN(new_n1155));
  OAI21_X1  g729(.A(new_n1155), .B1(KEYINPUT43), .B2(new_n941), .ZN(new_n1156));
  NAND4_X1  g730(.A1(new_n1156), .A2(new_n878), .A3(new_n1152), .A4(new_n1150), .ZN(G225));
endmodule


