//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 0 0 0 0 0 1 0 1 0 1 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 0 1 1 0 1 0 0 1 1 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n488, new_n489,
    new_n490, new_n491, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n507, new_n508, new_n509, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n553, new_n555, new_n556, new_n557, new_n558, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n628, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  INV_X1    g031(.A(G2104), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(KEYINPUT3), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n457), .A2(G2105), .ZN(new_n463));
  AOI22_X1  g038(.A1(new_n462), .A2(G137), .B1(G101), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n465), .B1(new_n461), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(G160));
  NAND2_X1  g045(.A1(new_n462), .A2(G136), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n461), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G124), .ZN(new_n474));
  OR2_X1    g049(.A1(G100), .A2(G2105), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n475), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n471), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G162));
  NOR2_X1   g053(.A1(new_n472), .A2(G114), .ZN(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n480));
  OAI21_X1  g055(.A(KEYINPUT65), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  OR3_X1    g056(.A1(new_n479), .A2(new_n480), .A3(KEYINPUT65), .ZN(new_n482));
  AOI22_X1  g057(.A1(new_n481), .A2(new_n482), .B1(new_n473), .B2(G126), .ZN(new_n483));
  NAND4_X1  g058(.A1(new_n458), .A2(new_n460), .A3(G138), .A4(new_n472), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT4), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G164));
  INV_X1    g062(.A(KEYINPUT5), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G543), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT67), .ZN(new_n490));
  INV_X1    g065(.A(G543), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(KEYINPUT5), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n488), .A2(KEYINPUT67), .A3(G543), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n489), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G651), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(KEYINPUT6), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT66), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT6), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(G651), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n495), .A2(KEYINPUT66), .A3(KEYINPUT6), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n496), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n494), .A2(new_n501), .A3(G88), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n501), .A2(G50), .A3(G543), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n494), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n502), .B(new_n503), .C1(new_n504), .C2(new_n495), .ZN(G303));
  INV_X1    g080(.A(G303), .ZN(G166));
  NAND3_X1  g081(.A1(new_n494), .A2(new_n501), .A3(G89), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n501), .A2(G51), .A3(G543), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT68), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n491), .A2(KEYINPUT5), .ZN(new_n511));
  AND3_X1   g086(.A1(new_n488), .A2(KEYINPUT67), .A3(G543), .ZN(new_n512));
  AOI21_X1  g087(.A(KEYINPUT67), .B1(new_n488), .B2(G543), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(G63), .A2(G651), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n510), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AOI221_X4 g091(.A(new_n515), .B1(KEYINPUT5), .B2(new_n491), .C1(new_n492), .C2(new_n493), .ZN(new_n517));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT69), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT69), .ZN(new_n520));
  NAND4_X1  g095(.A1(new_n520), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT7), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT7), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n519), .A2(new_n524), .A3(new_n521), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n517), .A2(KEYINPUT68), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  AND3_X1   g101(.A1(new_n509), .A2(new_n516), .A3(new_n526), .ZN(G168));
  NAND3_X1  g102(.A1(new_n494), .A2(new_n501), .A3(G90), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n501), .A2(G52), .A3(G543), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n530));
  AND3_X1   g105(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n530), .B1(new_n528), .B2(new_n529), .ZN(new_n532));
  AND2_X1   g107(.A1(G77), .A2(G543), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n533), .B1(new_n494), .B2(G64), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT70), .ZN(new_n535));
  OAI21_X1  g110(.A(G651), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AOI211_X1 g111(.A(KEYINPUT70), .B(new_n533), .C1(new_n494), .C2(G64), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n531), .A2(new_n532), .B1(new_n536), .B2(new_n537), .ZN(G301));
  INV_X1    g113(.A(G301), .ZN(G171));
  NAND3_X1  g114(.A1(new_n494), .A2(new_n501), .A3(G81), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n501), .A2(G43), .A3(G543), .ZN(new_n541));
  AND2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g117(.A(G56), .B(new_n511), .C1(new_n512), .C2(new_n513), .ZN(new_n543));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n495), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  AOI21_X1  g121(.A(KEYINPUT72), .B1(new_n542), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n540), .A2(new_n541), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT72), .ZN(new_n549));
  NOR3_X1   g124(.A1(new_n548), .A2(new_n545), .A3(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  AND3_X1   g127(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G36), .ZN(G176));
  XOR2_X1   g129(.A(KEYINPUT73), .B(KEYINPUT8), .Z(new_n555));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n555), .B(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  XOR2_X1   g133(.A(new_n558), .B(KEYINPUT74), .Z(G188));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n560), .A2(KEYINPUT75), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n501), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G53), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n561), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n501), .A2(G53), .A3(G543), .A4(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n494), .A2(new_n501), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G91), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT76), .ZN(new_n572));
  XNOR2_X1  g147(.A(KEYINPUT77), .B(G65), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n514), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G651), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n567), .A2(new_n570), .A3(new_n575), .ZN(G299));
  NAND3_X1  g151(.A1(new_n509), .A2(new_n516), .A3(new_n526), .ZN(G286));
  OAI21_X1  g152(.A(G651), .B1(new_n494), .B2(G74), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n494), .A2(new_n501), .A3(G87), .ZN(new_n579));
  AND2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n499), .A2(new_n500), .ZN(new_n581));
  INV_X1    g156(.A(new_n496), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(G49), .A2(G543), .ZN(new_n584));
  OAI21_X1  g159(.A(KEYINPUT78), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT78), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n501), .A2(new_n586), .A3(G49), .A4(G543), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n580), .A2(new_n588), .ZN(G288));
  NAND3_X1  g164(.A1(new_n494), .A2(new_n501), .A3(G86), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n501), .A2(G48), .A3(G543), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  OAI211_X1 g168(.A(G61), .B(new_n511), .C1(new_n512), .C2(new_n513), .ZN(new_n594));
  NAND2_X1  g169(.A1(G73), .A2(G543), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(KEYINPUT79), .B1(new_n596), .B2(G651), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT79), .ZN(new_n598));
  AOI211_X1 g173(.A(new_n598), .B(new_n495), .C1(new_n594), .C2(new_n595), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n593), .B1(new_n597), .B2(new_n599), .ZN(G305));
  NAND3_X1  g175(.A1(new_n494), .A2(new_n501), .A3(G85), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n501), .A2(G47), .A3(G543), .ZN(new_n602));
  AND2_X1   g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(G72), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n605), .B1(new_n494), .B2(G60), .ZN(new_n606));
  OAI21_X1  g181(.A(G651), .B1(new_n606), .B2(KEYINPUT80), .ZN(new_n607));
  OAI211_X1 g182(.A(G60), .B(new_n511), .C1(new_n512), .C2(new_n513), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(new_n604), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT80), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n603), .B1(new_n607), .B2(new_n611), .ZN(G290));
  NAND2_X1  g187(.A1(G301), .A2(G868), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n494), .A2(new_n501), .A3(G92), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT10), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(G79), .A2(G543), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT81), .ZN(new_n618));
  INV_X1    g193(.A(G66), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n514), .B2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(new_n562), .ZN(new_n621));
  AOI22_X1  g196(.A1(G651), .A2(new_n620), .B1(new_n621), .B2(G54), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n616), .A2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n613), .B1(new_n624), .B2(G868), .ZN(G284));
  OAI21_X1  g200(.A(new_n613), .B1(new_n624), .B2(G868), .ZN(G321));
  NAND2_X1  g201(.A1(G286), .A2(G868), .ZN(new_n627));
  INV_X1    g202(.A(G299), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(G868), .ZN(G297));
  OAI21_X1  g204(.A(new_n627), .B1(new_n628), .B2(G868), .ZN(G280));
  INV_X1    g205(.A(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n624), .B1(new_n631), .B2(G860), .ZN(G148));
  INV_X1    g207(.A(KEYINPUT82), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n624), .A2(new_n631), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n633), .B1(new_n634), .B2(G868), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(G868), .B2(new_n551), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n634), .A2(new_n633), .A3(G868), .ZN(new_n637));
  AND2_X1   g212(.A1(new_n636), .A2(new_n637), .ZN(G323));
  XNOR2_X1  g213(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g214(.A1(new_n462), .A2(G2104), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT12), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT13), .ZN(new_n642));
  INV_X1    g217(.A(G2100), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n462), .A2(G135), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n473), .A2(G123), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n472), .A2(G111), .ZN(new_n648));
  OAI21_X1  g223(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n649));
  OAI211_X1 g224(.A(new_n646), .B(new_n647), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(G2096), .Z(new_n651));
  NAND3_X1  g226(.A1(new_n644), .A2(new_n645), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT83), .Z(G156));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2435), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2438), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2427), .B(G2430), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  XOR2_X1   g233(.A(KEYINPUT85), .B(KEYINPUT14), .Z(new_n659));
  NAND3_X1  g234(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G1341), .B(G1348), .Z(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n660), .B(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2451), .B(G2454), .Z(new_n665));
  XNOR2_X1  g240(.A(G2443), .B(G2446), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n664), .A2(new_n667), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n668), .A2(G14), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT86), .Z(G401));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g249(.A1(new_n674), .A2(KEYINPUT17), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n672), .A2(new_n673), .ZN(new_n676));
  AOI21_X1  g251(.A(KEYINPUT18), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2072), .B(G2078), .Z(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(new_n674), .B2(KEYINPUT18), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n677), .B(new_n679), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(G2100), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT87), .B(G2096), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n681), .A2(new_n682), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(new_n684), .ZN(G227));
  XOR2_X1   g260(.A(KEYINPUT88), .B(KEYINPUT19), .Z(new_n686));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1956), .B(G2474), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1961), .B(G1966), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n689), .B(new_n690), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n689), .A2(new_n690), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n688), .A2(new_n693), .ZN(new_n694));
  AND2_X1   g269(.A1(new_n694), .A2(KEYINPUT20), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n694), .A2(KEYINPUT20), .ZN(new_n696));
  OAI221_X1 g271(.A(new_n691), .B1(new_n688), .B2(new_n692), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(G1991), .B(G1996), .Z(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n699), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1981), .B(G1986), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n699), .B(new_n700), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(new_n703), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(G229));
  MUX2_X1   g284(.A(G23), .B(G288), .S(G16), .Z(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT33), .B(G1976), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G6), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n494), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n598), .B1(new_n715), .B2(new_n495), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n596), .A2(KEYINPUT79), .A3(G651), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n592), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n714), .B1(new_n718), .B2(new_n713), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT32), .B(G1981), .Z(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT89), .B(G16), .ZN(new_n722));
  MUX2_X1   g297(.A(G303), .B(G22), .S(new_n722), .Z(new_n723));
  INV_X1    g298(.A(G1971), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  AND3_X1   g300(.A1(new_n712), .A2(new_n721), .A3(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT34), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n726), .A2(new_n727), .ZN(new_n729));
  MUX2_X1   g304(.A(G290), .B(G24), .S(new_n722), .Z(new_n730));
  AND2_X1   g305(.A1(new_n730), .A2(G1986), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n730), .A2(G1986), .ZN(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G25), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n462), .A2(G131), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n473), .A2(G119), .ZN(new_n736));
  OR2_X1    g311(.A1(G95), .A2(G2105), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n737), .B(G2104), .C1(G107), .C2(new_n472), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n735), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n734), .B1(new_n740), .B2(new_n733), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT35), .B(G1991), .Z(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n741), .B(new_n743), .ZN(new_n744));
  NOR3_X1   g319(.A1(new_n731), .A2(new_n732), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n728), .A2(new_n729), .A3(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT90), .ZN(new_n747));
  AND2_X1   g322(.A1(new_n747), .A2(KEYINPUT36), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n746), .B(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n733), .A2(G35), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G162), .B2(new_n733), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT29), .Z(new_n752));
  INV_X1    g327(.A(G2090), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(G1348), .ZN(new_n755));
  NOR2_X1   g330(.A1(G4), .A2(G16), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n624), .B2(G16), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n754), .A2(KEYINPUT100), .B1(new_n755), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n722), .A2(G20), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT23), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n628), .B2(new_n713), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT101), .B(G1956), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n759), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n733), .A2(G26), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT28), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n462), .A2(G140), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n473), .A2(G128), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n472), .A2(G116), .ZN(new_n770));
  OAI21_X1  g345(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n768), .B(new_n769), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n767), .B1(new_n772), .B2(G29), .ZN(new_n773));
  INV_X1    g348(.A(G2067), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT31), .B(G11), .Z(new_n776));
  INV_X1    g351(.A(KEYINPUT30), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n733), .B1(new_n777), .B2(G28), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n778), .A2(KEYINPUT98), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n777), .B2(G28), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n778), .A2(KEYINPUT98), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n776), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(G34), .ZN(new_n783));
  AOI21_X1  g358(.A(G29), .B1(new_n783), .B2(KEYINPUT24), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(KEYINPUT24), .B2(new_n783), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n469), .B2(new_n733), .ZN(new_n786));
  INV_X1    g361(.A(G2084), .ZN(new_n787));
  OAI221_X1 g362(.A(new_n782), .B1(new_n733), .B2(new_n650), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n775), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(G27), .A2(G29), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G164), .B2(G29), .ZN(new_n791));
  INV_X1    g366(.A(G2078), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n789), .B(new_n793), .C1(new_n754), .C2(KEYINPUT100), .ZN(new_n794));
  OAI22_X1  g369(.A1(new_n758), .A2(new_n755), .B1(new_n762), .B2(new_n763), .ZN(new_n795));
  OR3_X1    g370(.A1(new_n765), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(G5), .A2(G16), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT99), .Z(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G301), .B2(new_n713), .ZN(new_n799));
  INV_X1    g374(.A(G1961), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT92), .B(KEYINPUT26), .Z(new_n802));
  NAND3_X1  g377(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n463), .A2(G105), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n473), .A2(G129), .ZN(new_n807));
  INV_X1    g382(.A(G141), .ZN(new_n808));
  INV_X1    g383(.A(new_n462), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n806), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n811), .A2(new_n733), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n733), .B2(G32), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT93), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT27), .B(G1996), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT94), .Z(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n814), .A2(new_n817), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n786), .A2(new_n787), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n733), .A2(G33), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT25), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n458), .A2(new_n460), .A3(G127), .ZN(new_n824));
  NAND2_X1  g399(.A1(G115), .A2(G2104), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n472), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AOI211_X1 g401(.A(new_n823), .B(new_n826), .C1(G139), .C2(new_n462), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n821), .B1(new_n827), .B2(new_n733), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n820), .B1(new_n828), .B2(G2072), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(G2072), .B2(new_n828), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n752), .A2(new_n753), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n818), .A2(new_n819), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(G286), .A2(new_n713), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT95), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(G16), .B2(G21), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(KEYINPUT95), .B2(new_n833), .ZN(new_n837));
  XNOR2_X1  g412(.A(KEYINPUT96), .B(G1966), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(new_n800), .B2(new_n799), .ZN(new_n840));
  NOR4_X1   g415(.A1(new_n796), .A2(new_n801), .A3(new_n832), .A4(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n722), .A2(G19), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(new_n551), .B2(new_n722), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT91), .ZN(new_n844));
  INV_X1    g419(.A(G1341), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n837), .A2(new_n838), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT97), .Z(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(new_n845), .B2(new_n844), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n749), .A2(new_n841), .A3(new_n846), .A4(new_n849), .ZN(G150));
  INV_X1    g425(.A(G150), .ZN(G311));
  NAND3_X1  g426(.A1(new_n501), .A2(G55), .A3(G543), .ZN(new_n852));
  INV_X1    g427(.A(G93), .ZN(new_n853));
  AOI22_X1  g428(.A1(new_n494), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n854));
  OAI221_X1 g429(.A(new_n852), .B1(new_n568), .B2(new_n853), .C1(new_n854), .C2(new_n495), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(new_n547), .B2(new_n550), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n852), .B1(new_n568), .B2(new_n853), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n494), .A2(G67), .ZN(new_n858));
  NAND2_X1  g433(.A1(G80), .A2(G543), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n495), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n861), .A2(new_n546), .A3(new_n542), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n856), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT38), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n624), .A2(G559), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT39), .ZN(new_n867));
  AOI21_X1  g442(.A(G860), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n868), .B1(new_n867), .B2(new_n866), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n855), .A2(G860), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(KEYINPUT37), .Z(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT102), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(G145));
  XNOR2_X1  g449(.A(new_n811), .B(new_n772), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n875), .A2(new_n486), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n486), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n827), .B(KEYINPUT103), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT103), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n876), .A2(new_n881), .A3(new_n827), .A4(new_n877), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT105), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n473), .A2(G130), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n472), .A2(G118), .ZN(new_n886));
  OAI21_X1  g461(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n888), .B1(G142), .B2(new_n462), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(new_n641), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(new_n740), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n883), .B1(new_n884), .B2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n650), .B(new_n469), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(new_n477), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n880), .A2(KEYINPUT105), .A3(new_n891), .A4(new_n882), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n893), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(G37), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n880), .A2(new_n882), .A3(new_n891), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(KEYINPUT104), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n891), .B1(new_n880), .B2(new_n882), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT104), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n883), .A2(new_n904), .A3(new_n892), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(new_n895), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n898), .B(new_n899), .C1(new_n903), .C2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g483(.A(KEYINPUT107), .ZN(new_n909));
  NAND2_X1  g484(.A1(G290), .A2(G288), .ZN(new_n910));
  NAND2_X1  g485(.A1(G305), .A2(G166), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n609), .A2(new_n610), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n606), .A2(KEYINPUT80), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(new_n913), .A3(G651), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n914), .A2(new_n588), .A3(new_n580), .A4(new_n603), .ZN(new_n915));
  OAI211_X1 g490(.A(G303), .B(new_n593), .C1(new_n597), .C2(new_n599), .ZN(new_n916));
  AND4_X1   g491(.A1(new_n910), .A2(new_n911), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  AOI22_X1  g492(.A1(new_n911), .A2(new_n916), .B1(new_n910), .B2(new_n915), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n909), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n911), .A2(new_n916), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n910), .A2(new_n915), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n911), .A2(new_n910), .A3(new_n915), .A4(new_n916), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(KEYINPUT107), .A3(new_n923), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n919), .A2(KEYINPUT42), .A3(new_n924), .ZN(new_n925));
  XOR2_X1   g500(.A(new_n925), .B(KEYINPUT108), .Z(new_n926));
  XOR2_X1   g501(.A(new_n863), .B(new_n634), .Z(new_n927));
  NAND2_X1  g502(.A1(new_n623), .A2(G299), .ZN(new_n928));
  AOI22_X1  g503(.A1(G91), .A2(new_n569), .B1(new_n574), .B2(G651), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n616), .A2(new_n929), .A3(new_n622), .A4(new_n567), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT41), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n928), .A2(KEYINPUT41), .A3(new_n930), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n927), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(KEYINPUT106), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n927), .A2(new_n938), .A3(new_n935), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n937), .B(new_n939), .C1(new_n927), .C2(new_n931), .ZN(new_n940));
  XNOR2_X1  g515(.A(KEYINPUT109), .B(KEYINPUT42), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n941), .B1(new_n917), .B2(new_n918), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n926), .A2(new_n940), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n940), .B1(new_n926), .B2(new_n942), .ZN(new_n944));
  OAI21_X1  g519(.A(G868), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n861), .A2(G868), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(G295));
  NAND2_X1  g522(.A1(new_n945), .A2(new_n946), .ZN(G331));
  NOR2_X1   g523(.A1(G301), .A2(G168), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n528), .A2(new_n529), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT71), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n494), .A2(G64), .ZN(new_n954));
  OAI21_X1  g529(.A(KEYINPUT70), .B1(new_n954), .B2(new_n533), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n534), .A2(new_n535), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n955), .A2(G651), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(G286), .B1(new_n953), .B2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n542), .A2(new_n546), .A3(KEYINPUT72), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n549), .B1(new_n548), .B2(new_n545), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n861), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NOR3_X1   g536(.A1(new_n855), .A2(new_n545), .A3(new_n548), .ZN(new_n962));
  OAI22_X1  g537(.A1(new_n949), .A2(new_n958), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(G301), .A2(G168), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n953), .A2(new_n957), .A3(G286), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n856), .A2(new_n964), .A3(new_n862), .A4(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n931), .B1(new_n963), .B2(new_n966), .ZN(new_n967));
  AND4_X1   g542(.A1(new_n856), .A2(new_n964), .A3(new_n862), .A4(new_n965), .ZN(new_n968));
  AOI22_X1  g543(.A1(new_n856), .A2(new_n862), .B1(new_n964), .B2(new_n965), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n967), .B1(new_n935), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n924), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT107), .B1(new_n922), .B2(new_n923), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(G37), .B1(new_n971), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n931), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n976), .B1(new_n968), .B2(new_n969), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n933), .A2(new_n963), .A3(new_n934), .A4(new_n966), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n919), .A2(new_n924), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n975), .A2(new_n981), .ZN(new_n982));
  XOR2_X1   g557(.A(KEYINPUT110), .B(KEYINPUT43), .Z(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n981), .A2(KEYINPUT111), .ZN(new_n986));
  AOI22_X1  g561(.A1(new_n977), .A2(new_n978), .B1(new_n919), .B2(new_n924), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n986), .A2(new_n975), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n985), .B1(new_n984), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT44), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n977), .A2(new_n978), .A3(new_n919), .A4(new_n924), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n899), .B(new_n994), .C1(new_n987), .C2(new_n988), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n981), .A2(KEYINPUT111), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT112), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT113), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT112), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n986), .A2(new_n975), .A3(new_n989), .A4(new_n999), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n997), .A2(new_n998), .A3(KEYINPUT43), .A4(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n982), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n992), .B1(new_n1002), .B2(new_n983), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT43), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1005), .B1(new_n990), .B2(KEYINPUT112), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n998), .B1(new_n1006), .B2(new_n1000), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n993), .B1(new_n1004), .B2(new_n1007), .ZN(G397));
  INV_X1    g583(.A(G1384), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n486), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT45), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n464), .A2(G40), .A3(new_n468), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n772), .B(new_n774), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n1015), .B(KEYINPUT115), .ZN(new_n1016));
  INV_X1    g591(.A(G1996), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n811), .B(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1014), .ZN(new_n1020));
  OR3_X1    g595(.A1(new_n1019), .A2(KEYINPUT116), .A3(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT116), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1022));
  AND4_X1   g597(.A1(new_n742), .A2(new_n1021), .A3(new_n740), .A4(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n772), .A2(G2067), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1014), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n739), .B(new_n743), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1014), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1021), .A2(new_n1022), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT126), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT126), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1021), .A2(new_n1022), .A3(new_n1030), .A4(new_n1027), .ZN(new_n1031));
  OR3_X1    g606(.A1(new_n1020), .A2(G1986), .A3(G290), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n1032), .B(KEYINPUT48), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1029), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n811), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1014), .B1(new_n1016), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT46), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1037), .B1(new_n1020), .B2(G1996), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1014), .A2(KEYINPUT46), .A3(new_n1017), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1036), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  XOR2_X1   g615(.A(KEYINPUT125), .B(KEYINPUT47), .Z(new_n1041));
  XNOR2_X1  g616(.A(new_n1040), .B(new_n1041), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n1025), .A2(new_n1034), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT63), .ZN(new_n1044));
  NAND2_X1  g619(.A1(G168), .A2(G8), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1013), .ZN(new_n1046));
  AOI21_X1  g621(.A(G1384), .B1(new_n483), .B2(new_n485), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1046), .B1(new_n1047), .B2(KEYINPUT45), .ZN(new_n1048));
  AOI211_X1 g623(.A(new_n1011), .B(G1384), .C1(new_n483), .C2(new_n485), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n838), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1010), .A2(KEYINPUT50), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT50), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1047), .A2(new_n1052), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1051), .A2(new_n787), .A3(new_n1046), .A4(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1045), .B1(new_n1050), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(G8), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n724), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1057));
  XOR2_X1   g632(.A(KEYINPUT117), .B(G2090), .Z(new_n1058));
  NAND4_X1  g633(.A1(new_n1051), .A2(new_n1046), .A3(new_n1053), .A4(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1056), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(G303), .A2(G8), .ZN(new_n1061));
  XNOR2_X1  g636(.A(new_n1061), .B(KEYINPUT55), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1044), .B(new_n1055), .C1(new_n1060), .C2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT118), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1065), .A2(new_n1056), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1057), .A2(new_n1059), .A3(KEYINPUT118), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1064), .B1(new_n1068), .B2(new_n1062), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT119), .ZN(new_n1070));
  AOI211_X1 g645(.A(new_n1070), .B(new_n1056), .C1(new_n1047), .C2(new_n1046), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT119), .B1(new_n1072), .B2(G8), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  OR2_X1    g650(.A1(G305), .A2(G1981), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n715), .A2(new_n495), .ZN(new_n1077));
  OAI21_X1  g652(.A(G1981), .B1(new_n1077), .B2(new_n592), .ZN(new_n1078));
  AOI21_X1  g653(.A(KEYINPUT49), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1076), .A2(KEYINPUT49), .A3(new_n1078), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1075), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(G1976), .ZN(new_n1083));
  NOR2_X1   g658(.A1(G288), .A2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT52), .B1(new_n1074), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT52), .B1(G288), .B2(new_n1083), .ZN(new_n1086));
  OAI221_X1 g661(.A(new_n1086), .B1(new_n1083), .B2(G288), .C1(new_n1071), .C2(new_n1073), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1082), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1081), .ZN(new_n1089));
  NOR3_X1   g664(.A1(new_n1089), .A2(new_n1074), .A3(new_n1079), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n580), .A2(new_n588), .A3(new_n1083), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1076), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AOI22_X1  g667(.A1(new_n1069), .A2(new_n1088), .B1(new_n1092), .B2(new_n1075), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT120), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1068), .A2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1082), .A2(new_n1085), .A3(new_n1087), .A4(new_n1055), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1062), .A2(new_n1094), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1097), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1098));
  NOR3_X1   g673(.A1(new_n1095), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1093), .B1(new_n1099), .B2(new_n1044), .ZN(new_n1100));
  INV_X1    g675(.A(G1956), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1046), .B1(new_n1047), .B2(new_n1052), .ZN(new_n1102));
  AOI211_X1 g677(.A(KEYINPUT50), .B(G1384), .C1(new_n483), .C2(new_n485), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1101), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1047), .A2(KEYINPUT45), .ZN(new_n1105));
  XNOR2_X1  g680(.A(KEYINPUT56), .B(G2072), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1012), .A2(new_n1046), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT57), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1110), .B1(new_n929), .B2(new_n567), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1104), .A2(new_n1107), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1114), .A2(new_n1104), .A3(new_n1107), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n755), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1047), .A2(new_n1046), .A3(new_n774), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n623), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1113), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT61), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1114), .A2(new_n1104), .A3(new_n1107), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1120), .B1(new_n1121), .B2(new_n1113), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1104), .A2(new_n1107), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1114), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1125), .A2(KEYINPUT61), .A3(new_n1115), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1116), .A2(new_n1117), .A3(new_n623), .ZN(new_n1127));
  OAI21_X1  g702(.A(KEYINPUT60), .B1(new_n1127), .B2(new_n1118), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1122), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n623), .A2(KEYINPUT60), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1116), .A2(new_n1117), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT59), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1013), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1133), .A2(new_n1017), .A3(new_n1105), .ZN(new_n1134));
  XOR2_X1   g709(.A(KEYINPUT58), .B(G1341), .Z(new_n1135));
  NAND2_X1  g710(.A1(new_n1072), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1132), .B1(new_n1137), .B2(new_n551), .ZN(new_n1138));
  INV_X1    g713(.A(new_n551), .ZN(new_n1139));
  AOI211_X1 g714(.A(KEYINPUT59), .B(new_n1139), .C1(new_n1134), .C2(new_n1136), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1131), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1119), .B1(new_n1129), .B2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1143), .A2(KEYINPUT53), .A3(new_n792), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n800), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(KEYINPUT121), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT121), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1144), .A2(new_n1148), .A3(new_n1145), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT53), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1143), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1150), .B1(new_n1151), .B2(G2078), .ZN(new_n1152));
  XOR2_X1   g727(.A(G301), .B(KEYINPUT54), .Z(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1147), .A2(new_n1149), .A3(new_n1152), .A4(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(KEYINPUT53), .B1(KEYINPUT123), .B2(G2078), .ZN(new_n1156));
  AOI211_X1 g731(.A(new_n1156), .B(new_n1049), .C1(KEYINPUT123), .C2(G2078), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n1133), .A2(KEYINPUT122), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1133), .A2(KEYINPUT122), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1160), .A2(new_n1152), .A3(new_n1145), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(new_n1153), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1050), .A2(new_n1054), .A3(G168), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(G8), .ZN(new_n1164));
  AOI21_X1  g739(.A(G168), .B1(new_n1050), .B2(new_n1054), .ZN(new_n1165));
  OAI21_X1  g740(.A(KEYINPUT51), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT51), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1163), .A2(new_n1167), .A3(G8), .ZN(new_n1168));
  AOI22_X1  g743(.A1(new_n1155), .A2(new_n1162), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1142), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT124), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT62), .ZN(new_n1172));
  AOI22_X1  g747(.A1(new_n1166), .A2(new_n1168), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1174));
  AND2_X1   g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  AND2_X1   g750(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1176));
  AOI21_X1  g751(.A(G301), .B1(new_n1176), .B2(new_n1147), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1177), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1170), .B1(new_n1175), .B2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1088), .B1(new_n1063), .B2(new_n1060), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1068), .A2(new_n1062), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1100), .B1(new_n1179), .B2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1014), .A2(G1986), .A3(G290), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1032), .A2(new_n1184), .ZN(new_n1185));
  XOR2_X1   g760(.A(new_n1185), .B(KEYINPUT114), .Z(new_n1186));
  OR2_X1    g761(.A1(new_n1186), .A2(new_n1028), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1043), .B1(new_n1183), .B2(new_n1187), .ZN(G329));
  assign    G231 = 1'b0;
  NAND4_X1  g763(.A1(new_n683), .A2(G319), .A3(new_n670), .A4(new_n684), .ZN(new_n1190));
  INV_X1    g764(.A(new_n1190), .ZN(new_n1191));
  AOI21_X1  g765(.A(KEYINPUT127), .B1(new_n708), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g766(.A(KEYINPUT127), .ZN(new_n1193));
  AOI211_X1 g767(.A(new_n1193), .B(new_n1190), .C1(new_n705), .C2(new_n707), .ZN(new_n1194));
  OAI211_X1 g768(.A(new_n907), .B(new_n991), .C1(new_n1192), .C2(new_n1194), .ZN(G225));
  INV_X1    g769(.A(G225), .ZN(G308));
endmodule


