//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 0 1 0 0 1 0 1 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n556, new_n557, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n592, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n631, new_n632, new_n635, new_n636, new_n638, new_n639, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1238,
    new_n1239, new_n1240;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT65), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT66), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT67), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(new_n451), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n455), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(G125), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT68), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(new_n466), .A3(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n464), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n465), .A2(G137), .A3(new_n471), .ZN(new_n474));
  AND3_X1   g049(.A1(new_n470), .A2(new_n473), .A3(new_n474), .ZN(G160));
  NOR2_X1   g050(.A1(new_n461), .A2(new_n462), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  XOR2_X1   g053(.A(new_n478), .B(KEYINPUT69), .Z(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(G112), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n480), .B1(new_n481), .B2(G2105), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n476), .A2(new_n471), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(new_n483), .B2(G124), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n479), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  OAI21_X1  g062(.A(G2105), .B1(KEYINPUT70), .B2(G114), .ZN(new_n488));
  AND2_X1   g063(.A1(KEYINPUT70), .A2(G114), .ZN(new_n489));
  OAI211_X1 g064(.A(G2104), .B(new_n487), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  OAI211_X1 g065(.A(G126), .B(G2105), .C1(new_n461), .C2(new_n462), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT71), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n490), .A2(new_n491), .A3(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT72), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n497), .A2(new_n471), .A3(G138), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n496), .B1(new_n476), .B2(new_n498), .ZN(new_n499));
  AND3_X1   g074(.A1(new_n497), .A2(new_n471), .A3(G138), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n465), .A2(new_n500), .A3(KEYINPUT72), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g077(.A(G138), .B(new_n471), .C1(new_n461), .C2(new_n462), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT4), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n493), .A2(new_n495), .B1(new_n502), .B2(new_n504), .ZN(G164));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  OAI21_X1  g083(.A(G62), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(G75), .A2(G543), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g089(.A(G88), .B1(new_n507), .B2(new_n508), .ZN(new_n515));
  NAND2_X1  g090(.A1(G50), .A2(G543), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n511), .A2(new_n517), .ZN(G166));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT6), .B(G651), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT73), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n513), .ZN(new_n523));
  NAND2_X1  g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n523), .A2(KEYINPUT73), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n522), .A2(G51), .A3(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n507), .A2(new_n508), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n527), .A2(new_n514), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G89), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  OR2_X1    g106(.A1(KEYINPUT5), .A2(G543), .ZN(new_n532));
  NAND2_X1  g107(.A1(KEYINPUT5), .A2(G543), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n534), .A2(G63), .A3(G651), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n526), .A2(new_n529), .A3(new_n531), .A4(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G64), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n527), .B2(new_n539), .ZN(new_n540));
  AOI22_X1  g115(.A1(G651), .A2(new_n540), .B1(new_n528), .B2(G90), .ZN(new_n541));
  XOR2_X1   g116(.A(KEYINPUT74), .B(G52), .Z(new_n542));
  NAND3_X1  g117(.A1(new_n522), .A2(new_n525), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n541), .A2(new_n543), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  NAND2_X1  g120(.A1(G68), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G56), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n527), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G651), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n528), .A2(G81), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n520), .A2(new_n521), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n551), .A2(G43), .A3(new_n525), .A4(G543), .ZN(new_n552));
  AND3_X1   g127(.A1(new_n549), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  XNOR2_X1  g133(.A(KEYINPUT76), .B(G65), .ZN(new_n559));
  INV_X1    g134(.A(G78), .ZN(new_n560));
  OAI22_X1  g135(.A1(new_n527), .A2(new_n559), .B1(new_n560), .B2(new_n519), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT77), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI221_X1 g138(.A(KEYINPUT77), .B1(new_n560), .B2(new_n519), .C1(new_n527), .C2(new_n559), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n563), .A2(G651), .A3(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT75), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n528), .A2(new_n566), .A3(G91), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n534), .A2(new_n520), .ZN(new_n568));
  INV_X1    g143(.A(G91), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT75), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n565), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n551), .A2(G53), .A3(new_n525), .A4(G543), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT9), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n573), .B(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT78), .ZN(new_n576));
  NOR3_X1   g151(.A1(new_n572), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  XOR2_X1   g152(.A(KEYINPUT76), .B(G65), .Z(new_n578));
  AOI22_X1  g153(.A1(new_n578), .A2(new_n534), .B1(G78), .B2(G543), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n506), .B1(new_n579), .B2(KEYINPUT77), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(new_n563), .B1(new_n570), .B2(new_n567), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n573), .B(KEYINPUT9), .ZN(new_n582));
  AOI21_X1  g157(.A(KEYINPUT78), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n577), .A2(new_n583), .ZN(G299));
  INV_X1    g159(.A(G88), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n585), .B1(new_n532), .B2(new_n533), .ZN(new_n586));
  INV_X1    g161(.A(new_n516), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n520), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT79), .ZN(new_n589));
  AND2_X1   g164(.A1(new_n509), .A2(new_n510), .ZN(new_n590));
  OAI211_X1 g165(.A(new_n588), .B(new_n589), .C1(new_n590), .C2(new_n506), .ZN(new_n591));
  OAI21_X1  g166(.A(KEYINPUT79), .B1(new_n511), .B2(new_n517), .ZN(new_n592));
  AND2_X1   g167(.A1(new_n591), .A2(new_n592), .ZN(G303));
  INV_X1    g168(.A(G74), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n527), .A2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n528), .A2(G87), .B1(new_n595), .B2(G651), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n522), .A2(G49), .A3(new_n525), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(G288));
  NAND2_X1  g173(.A1(G73), .A2(G543), .ZN(new_n599));
  XOR2_X1   g174(.A(new_n599), .B(KEYINPUT80), .Z(new_n600));
  INV_X1    g175(.A(G61), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n601), .B1(new_n532), .B2(new_n533), .ZN(new_n602));
  OAI21_X1  g177(.A(G651), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(G48), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G86), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n527), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(new_n520), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n603), .A2(new_n607), .ZN(G305));
  NAND2_X1  g183(.A1(new_n528), .A2(G85), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n534), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n522), .A2(new_n525), .ZN(new_n611));
  INV_X1    g186(.A(G47), .ZN(new_n612));
  OAI221_X1 g187(.A(new_n609), .B1(new_n610), .B2(new_n506), .C1(new_n611), .C2(new_n612), .ZN(G290));
  NAND2_X1  g188(.A1(G301), .A2(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(G79), .A2(G543), .ZN(new_n615));
  INV_X1    g190(.A(G66), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n527), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G651), .ZN(new_n618));
  INV_X1    g193(.A(G54), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n611), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(KEYINPUT81), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT81), .ZN(new_n622));
  OAI211_X1 g197(.A(new_n618), .B(new_n622), .C1(new_n611), .C2(new_n619), .ZN(new_n623));
  INV_X1    g198(.A(G92), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n568), .A2(new_n624), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n625), .A2(KEYINPUT10), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(KEYINPUT10), .ZN(new_n627));
  AOI22_X1  g202(.A1(new_n621), .A2(new_n623), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n614), .B1(new_n628), .B2(G868), .ZN(G284));
  OAI21_X1  g204(.A(new_n614), .B1(new_n628), .B2(G868), .ZN(G321));
  INV_X1    g205(.A(G868), .ZN(new_n631));
  NAND2_X1  g206(.A1(G299), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(new_n631), .B2(G168), .ZN(G297));
  OAI21_X1  g208(.A(new_n632), .B1(new_n631), .B2(G168), .ZN(G280));
  INV_X1    g209(.A(G559), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n628), .B1(new_n635), .B2(G860), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT82), .ZN(G148));
  NAND2_X1  g212(.A1(new_n628), .A2(new_n635), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(G868), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(G868), .B2(new_n553), .ZN(G323));
  XNOR2_X1  g215(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g216(.A1(new_n465), .A2(new_n472), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT12), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT13), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n645), .A2(G2100), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n483), .A2(G123), .ZN(new_n647));
  INV_X1    g222(.A(KEYINPUT83), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n650));
  INV_X1    g225(.A(G111), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n650), .B1(new_n651), .B2(G2105), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n652), .B1(new_n477), .B2(G135), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n654), .A2(G2096), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n645), .A2(G2100), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(G2096), .ZN(new_n657));
  NAND4_X1  g232(.A1(new_n646), .A2(new_n655), .A3(new_n656), .A4(new_n657), .ZN(G156));
  XNOR2_X1  g233(.A(KEYINPUT15), .B(G2435), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT84), .B(G2438), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2427), .B(G2430), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n663), .A2(KEYINPUT14), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT85), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n666), .A2(G1341), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(G1341), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(G1348), .ZN(new_n670));
  XOR2_X1   g245(.A(G2451), .B(G2454), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT16), .ZN(new_n672));
  XOR2_X1   g247(.A(G2443), .B(G2446), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(G1348), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n667), .A2(new_n675), .A3(new_n668), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n670), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(G14), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n674), .B1(new_n670), .B2(new_n676), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(G401));
  XNOR2_X1  g255(.A(G2067), .B(G2678), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT87), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G2084), .B(G2090), .Z(new_n684));
  OAI21_X1  g259(.A(KEYINPUT17), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G2072), .B(G2078), .Z(new_n686));
  AOI22_X1  g261(.A1(new_n685), .A2(new_n686), .B1(new_n684), .B2(new_n683), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(new_n686), .B2(new_n685), .ZN(new_n688));
  INV_X1    g263(.A(new_n686), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n689), .A2(new_n684), .A3(new_n681), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT86), .B(KEYINPUT18), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G2096), .B(G2100), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(G227));
  XOR2_X1   g270(.A(G1971), .B(G1976), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT19), .ZN(new_n697));
  XOR2_X1   g272(.A(G1956), .B(G2474), .Z(new_n698));
  XOR2_X1   g273(.A(G1961), .B(G1966), .Z(new_n699));
  AND2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n702));
  OR2_X1    g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n698), .A2(new_n699), .ZN(new_n705));
  OR3_X1    g280(.A1(new_n697), .A2(new_n700), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n697), .A2(new_n705), .ZN(new_n707));
  NAND4_X1  g282(.A1(new_n703), .A2(new_n704), .A3(new_n706), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G1981), .ZN(new_n709));
  INV_X1    g284(.A(G1986), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n709), .A2(new_n710), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT89), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n712), .A2(new_n713), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(G1991), .B(G1996), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n709), .A2(new_n710), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n715), .B1(new_n719), .B2(new_n711), .ZN(new_n720));
  AND3_X1   g295(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n718), .B1(new_n717), .B2(new_n720), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(G229));
  INV_X1    g298(.A(KEYINPUT94), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT36), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n724), .B1(new_n725), .B2(KEYINPUT93), .ZN(new_n726));
  MUX2_X1   g301(.A(G23), .B(G288), .S(G16), .Z(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT33), .B(G1976), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  MUX2_X1   g304(.A(G6), .B(G305), .S(G16), .Z(new_n730));
  XOR2_X1   g305(.A(KEYINPUT32), .B(G1981), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G16), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G22), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G166), .B2(new_n733), .ZN(new_n735));
  INV_X1    g310(.A(G1971), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n729), .A2(new_n732), .A3(new_n737), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n738), .A2(KEYINPUT34), .ZN(new_n739));
  INV_X1    g314(.A(G29), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G25), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT90), .Z(new_n742));
  NAND2_X1  g317(.A1(new_n477), .A2(G131), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n483), .A2(G119), .ZN(new_n744));
  INV_X1    g319(.A(G95), .ZN(new_n745));
  AND3_X1   g320(.A1(new_n745), .A2(new_n471), .A3(KEYINPUT91), .ZN(new_n746));
  AOI21_X1  g321(.A(KEYINPUT91), .B1(new_n745), .B2(new_n471), .ZN(new_n747));
  OAI221_X1 g322(.A(G2104), .B1(G107), .B2(new_n471), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n743), .A2(new_n744), .A3(new_n748), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n749), .A2(KEYINPUT92), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(KEYINPUT92), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n742), .B1(new_n752), .B2(G29), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT35), .B(G1991), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  MUX2_X1   g330(.A(G24), .B(G290), .S(G16), .Z(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G1986), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n738), .A2(KEYINPUT34), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n739), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n724), .A2(new_n725), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n726), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n726), .B2(new_n760), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n740), .A2(G32), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n472), .A2(G105), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n477), .A2(G141), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n483), .A2(G129), .ZN(new_n767));
  NAND3_X1  g342(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT26), .Z(new_n769));
  AND4_X1   g344(.A1(new_n765), .A2(new_n766), .A3(new_n767), .A4(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n764), .B1(new_n770), .B2(new_n740), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT27), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1996), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n477), .A2(G139), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT25), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n780), .A2(new_n471), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n782), .A2(new_n740), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n740), .B2(G33), .ZN(new_n784));
  INV_X1    g359(.A(G2072), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT24), .ZN(new_n787));
  INV_X1    g362(.A(G34), .ZN(new_n788));
  AOI21_X1  g363(.A(G29), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n787), .B2(new_n788), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G160), .B2(new_n740), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(G2084), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n784), .A2(new_n785), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT31), .B(G11), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT30), .B(G28), .Z(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(G29), .ZN(new_n796));
  INV_X1    g371(.A(new_n654), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(G29), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n786), .A2(new_n792), .A3(new_n793), .A4(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n774), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n740), .A2(G26), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT28), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n477), .A2(G140), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n483), .A2(G128), .ZN(new_n804));
  OR2_X1    g379(.A1(G104), .A2(G2105), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n805), .B(G2104), .C1(G116), .C2(new_n471), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n803), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n802), .B1(new_n808), .B2(new_n740), .ZN(new_n809));
  INV_X1    g384(.A(G2067), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(G1341), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n553), .A2(G16), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G16), .B2(G19), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n811), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n812), .B2(new_n814), .ZN(new_n816));
  INV_X1    g391(.A(G35), .ZN(new_n817));
  OR3_X1    g392(.A1(new_n817), .A2(KEYINPUT101), .A3(G29), .ZN(new_n818));
  OAI21_X1  g393(.A(KEYINPUT101), .B1(new_n817), .B2(G29), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n818), .B(new_n819), .C1(G162), .C2(new_n740), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT29), .B(G2090), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n733), .A2(G5), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G171), .B2(new_n733), .ZN(new_n824));
  INV_X1    g399(.A(G1961), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n800), .A2(new_n816), .A3(new_n822), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(G299), .A2(G16), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n733), .A2(G20), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT23), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(G1956), .ZN(new_n832));
  NOR2_X1   g407(.A1(G4), .A2(G16), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT95), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n621), .A2(new_n623), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n626), .A2(new_n627), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n834), .B1(new_n837), .B2(new_n733), .ZN(new_n838));
  XOR2_X1   g413(.A(KEYINPUT96), .B(G1348), .Z(new_n839));
  NOR2_X1   g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT100), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n740), .A2(G27), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT99), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(G164), .B2(new_n740), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(G2078), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n840), .B1(new_n841), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n838), .A2(new_n839), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n846), .B(new_n847), .C1(new_n841), .C2(new_n845), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n791), .A2(G2084), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT98), .Z(new_n850));
  NAND2_X1  g425(.A1(new_n733), .A2(G21), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(G168), .B2(new_n733), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT97), .ZN(new_n853));
  INV_X1    g428(.A(G1966), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  NOR4_X1   g431(.A1(new_n827), .A2(new_n832), .A3(new_n848), .A4(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT102), .ZN(new_n858));
  AND3_X1   g433(.A1(new_n763), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n858), .B1(new_n763), .B2(new_n857), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(G311));
  NAND2_X1  g436(.A1(new_n763), .A2(new_n857), .ZN(G150));
  NAND2_X1  g437(.A1(G80), .A2(G543), .ZN(new_n863));
  INV_X1    g438(.A(G67), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n863), .B1(new_n527), .B2(new_n864), .ZN(new_n865));
  AOI22_X1  g440(.A1(G651), .A2(new_n865), .B1(new_n528), .B2(G93), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n522), .A2(G55), .A3(new_n525), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(G860), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(KEYINPUT37), .Z(new_n870));
  NAND2_X1  g445(.A1(new_n628), .A2(G559), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(KEYINPUT103), .Z(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT38), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n553), .A2(new_n867), .A3(new_n866), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n549), .A2(new_n550), .A3(new_n552), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n868), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n873), .B(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT39), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(G860), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n878), .A2(new_n879), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n870), .B1(new_n882), .B2(new_n883), .ZN(G145));
  NAND2_X1  g459(.A1(new_n770), .A2(new_n808), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n766), .A2(new_n767), .A3(new_n765), .A4(new_n769), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(new_n807), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n492), .B1(new_n502), .B2(new_n504), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR3_X1   g465(.A1(new_n476), .A2(new_n496), .A3(new_n498), .ZN(new_n891));
  AOI21_X1  g466(.A(KEYINPUT72), .B1(new_n465), .B2(new_n500), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n504), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n492), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n885), .A2(new_n887), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n890), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n782), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n890), .A2(new_n782), .A3(new_n896), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT105), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT104), .ZN(new_n903));
  INV_X1    g478(.A(new_n643), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n477), .A2(G142), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n483), .A2(G130), .ZN(new_n906));
  OR2_X1    g481(.A1(G106), .A2(G2105), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n907), .B(G2104), .C1(G118), .C2(new_n471), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n905), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n904), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n643), .A2(new_n905), .A3(new_n906), .A4(new_n908), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n750), .A2(new_n910), .A3(new_n751), .A4(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  AOI22_X1  g488(.A1(new_n751), .A2(new_n750), .B1(new_n910), .B2(new_n911), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n903), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n910), .A2(new_n911), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n752), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n917), .A2(KEYINPUT104), .A3(new_n912), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n901), .A2(new_n902), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n902), .B1(new_n901), .B2(new_n919), .ZN(new_n921));
  OAI22_X1  g496(.A1(new_n920), .A2(new_n921), .B1(new_n901), .B2(new_n919), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n485), .B(G160), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(new_n654), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(G37), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n920), .A2(new_n921), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n913), .A2(new_n914), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n899), .A2(new_n928), .A3(new_n900), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT106), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT106), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n899), .A2(new_n928), .A3(new_n931), .A4(new_n900), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n930), .A2(new_n932), .A3(new_n924), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT107), .ZN(new_n934));
  NOR3_X1   g509(.A1(new_n927), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n930), .A2(new_n932), .A3(new_n924), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n901), .A2(new_n919), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT105), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n901), .A2(new_n902), .A3(new_n919), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(KEYINPUT107), .B1(new_n936), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n926), .B1(new_n935), .B2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n942), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g518(.A(G290), .B(G305), .Z(new_n944));
  XNOR2_X1  g519(.A(G288), .B(G166), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n944), .B(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n946), .B(KEYINPUT42), .ZN(new_n947));
  XOR2_X1   g522(.A(new_n638), .B(new_n877), .Z(new_n948));
  OAI21_X1  g523(.A(new_n837), .B1(new_n577), .B2(new_n583), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n576), .B1(new_n572), .B2(new_n575), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n581), .A2(new_n582), .A3(KEYINPUT78), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(new_n628), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  OR2_X1    g529(.A1(new_n948), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT41), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n950), .A2(new_n628), .A3(new_n951), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n628), .B1(new_n950), .B2(new_n951), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n949), .A2(KEYINPUT41), .A3(new_n952), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n959), .A2(KEYINPUT108), .A3(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT108), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n953), .A2(new_n962), .A3(new_n956), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n961), .A2(new_n948), .A3(new_n963), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n947), .A2(new_n955), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n947), .B1(new_n955), .B2(new_n964), .ZN(new_n966));
  OAI21_X1  g541(.A(G868), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n868), .A2(new_n631), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(G295));
  NAND2_X1  g544(.A1(new_n967), .A2(new_n968), .ZN(G331));
  INV_X1    g545(.A(KEYINPUT43), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT109), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n535), .A2(new_n531), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n973), .B1(G89), .B2(new_n528), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n974), .A2(new_n526), .A3(new_n543), .A4(new_n541), .ZN(new_n975));
  NAND2_X1  g550(.A1(G301), .A2(G286), .ZN(new_n976));
  AND4_X1   g551(.A1(new_n876), .A2(new_n874), .A3(new_n975), .A4(new_n976), .ZN(new_n977));
  AOI22_X1  g552(.A1(new_n876), .A2(new_n874), .B1(new_n975), .B2(new_n976), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n972), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n975), .A2(new_n976), .ZN(new_n980));
  OAI21_X1  g555(.A(KEYINPUT109), .B1(new_n877), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n961), .A2(new_n963), .A3(new_n982), .ZN(new_n983));
  OR2_X1    g558(.A1(new_n977), .A2(new_n978), .ZN(new_n984));
  OR2_X1    g559(.A1(new_n954), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n983), .A2(new_n946), .A3(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G37), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n946), .B1(new_n983), .B2(new_n985), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n971), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n946), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n984), .B1(new_n960), .B2(KEYINPUT110), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n959), .A2(KEYINPUT110), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n992), .B1(new_n993), .B2(new_n960), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT111), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n995), .B1(new_n982), .B2(new_n954), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n953), .A2(new_n979), .A3(KEYINPUT111), .A4(new_n981), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n991), .B1(new_n994), .B2(new_n998), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n999), .A2(KEYINPUT43), .A3(new_n987), .A4(new_n986), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n990), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT44), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT43), .B1(new_n988), .B2(new_n989), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n999), .A2(new_n971), .A3(new_n987), .A4(new_n986), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT44), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1002), .A2(new_n1007), .ZN(G397));
  XNOR2_X1  g583(.A(new_n807), .B(G2067), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1009), .B(KEYINPUT113), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT112), .ZN(new_n1011));
  AOI22_X1  g586(.A1(new_n463), .A2(KEYINPUT68), .B1(G113), .B2(G2104), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n471), .B1(new_n1012), .B2(new_n467), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n474), .A2(G40), .A3(new_n473), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1011), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1014), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n470), .A2(KEYINPUT112), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT45), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1019), .B1(new_n889), .B2(G1384), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1010), .A2(new_n1022), .ZN(new_n1023));
  OR2_X1    g598(.A1(new_n1023), .A2(KEYINPUT114), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(KEYINPUT114), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n886), .B(G1996), .ZN(new_n1026));
  AOI22_X1  g601(.A1(new_n1024), .A2(new_n1025), .B1(new_n1021), .B2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n752), .B(new_n754), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1027), .B1(new_n1022), .B2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g604(.A(G290), .B(G1986), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1029), .B1(new_n1021), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(G1384), .B1(new_n893), .B2(new_n894), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1015), .A2(new_n1017), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n528), .A2(G87), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n595), .A2(G651), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n597), .A2(new_n1034), .A3(G1976), .A4(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT116), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n596), .A2(new_n1038), .A3(G1976), .A4(new_n597), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1033), .A2(new_n1040), .A3(G8), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT52), .ZN(new_n1042));
  INV_X1    g617(.A(G1976), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT52), .B1(G288), .B2(new_n1043), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1033), .A2(new_n1040), .A3(G8), .A4(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT49), .ZN(new_n1046));
  INV_X1    g621(.A(G1981), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n603), .A2(new_n1047), .A3(new_n607), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1047), .B1(new_n603), .B2(new_n607), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1046), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1050), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1052), .A2(KEYINPUT49), .A3(new_n1048), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1051), .A2(new_n1053), .A3(new_n1033), .A4(G8), .ZN(new_n1054));
  AND3_X1   g629(.A1(new_n1042), .A2(new_n1045), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1057));
  INV_X1    g632(.A(G2090), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n1060));
  INV_X1    g635(.A(G1384), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n895), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .A4(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1019), .A2(G1384), .ZN(new_n1064));
  AOI22_X1  g639(.A1(new_n499), .A2(new_n501), .B1(KEYINPUT4), .B2(new_n503), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1064), .B1(new_n1065), .B2(new_n492), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1015), .A2(new_n1017), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n494), .B1(new_n490), .B2(new_n491), .ZN(new_n1068));
  AND3_X1   g643(.A1(new_n490), .A2(new_n494), .A3(new_n491), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n893), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT45), .B1(new_n1070), .B2(new_n1061), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n736), .B1(new_n1067), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1063), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n591), .A2(new_n592), .A3(G8), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT55), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n591), .A2(new_n592), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OR2_X1    g653(.A1(new_n1078), .A2(KEYINPUT115), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(KEYINPUT115), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1073), .A2(new_n1079), .A3(G8), .A4(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1033), .A2(G8), .ZN(new_n1082));
  XNOR2_X1  g657(.A(new_n1048), .B(KEYINPUT117), .ZN(new_n1083));
  NOR2_X1   g658(.A1(G288), .A2(G1976), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1083), .B1(new_n1054), .B2(new_n1084), .ZN(new_n1085));
  OAI22_X1  g660(.A1(new_n1056), .A2(new_n1081), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT63), .ZN(new_n1087));
  INV_X1    g662(.A(G8), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1015), .B(new_n1017), .C1(new_n1032), .C2(new_n1060), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n1091));
  NOR2_X1   g666(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1091), .B1(G164), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1070), .A2(KEYINPUT118), .A3(new_n1092), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1090), .A2(new_n1058), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1088), .B1(new_n1096), .B2(new_n1072), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1081), .B(new_n1055), .C1(new_n1097), .C2(new_n1078), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1069), .A2(new_n1068), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1064), .B1(new_n1099), .B2(new_n1065), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1020), .A2(new_n1100), .A3(new_n1015), .A4(new_n1017), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n854), .ZN(new_n1102));
  INV_X1    g677(.A(G2084), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1057), .A2(new_n1103), .A3(new_n1059), .A4(new_n1062), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1105), .A2(G8), .A3(G168), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1087), .B1(new_n1098), .B2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1106), .A2(new_n1087), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1073), .A2(G8), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1109), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1108), .A2(new_n1081), .A3(new_n1055), .A4(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1086), .B1(new_n1107), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n493), .A2(new_n495), .ZN(new_n1113));
  AOI21_X1  g688(.A(G1384), .B1(new_n1113), .B2(new_n893), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1062), .B1(new_n1114), .B2(new_n1060), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n825), .B1(new_n1115), .B2(new_n1018), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT53), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1118), .A2(G2078), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1020), .A2(new_n1117), .A3(new_n1066), .A4(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1116), .A2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1067), .A2(new_n1071), .ZN(new_n1122));
  INV_X1    g697(.A(G2078), .ZN(new_n1123));
  AOI21_X1  g698(.A(KEYINPUT53), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(G171), .B1(new_n1121), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1019), .B1(G164), .B2(G1384), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1057), .A2(new_n1126), .A3(new_n1066), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1118), .B1(new_n1127), .B2(G2078), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1057), .A2(new_n1119), .A3(new_n1020), .A4(new_n1100), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1128), .A2(G301), .A3(new_n1116), .A4(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1125), .A2(new_n1130), .A3(KEYINPUT54), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(KEYINPUT124), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1125), .A2(new_n1130), .A3(new_n1133), .A4(KEYINPUT54), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT54), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1116), .A2(new_n1129), .ZN(new_n1137));
  OAI21_X1  g712(.A(G171), .B1(new_n1137), .B2(new_n1124), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  NOR3_X1   g714(.A1(new_n1121), .A2(new_n1124), .A3(G171), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1136), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1102), .A2(new_n1104), .A3(G168), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(G8), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1060), .B1(new_n1070), .B2(new_n1061), .ZN(new_n1144));
  NOR3_X1   g719(.A1(new_n889), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1018), .A2(G2084), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1146), .A2(new_n1147), .B1(new_n1101), .B2(new_n854), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1148), .A2(G168), .ZN(new_n1149));
  OAI21_X1  g724(.A(KEYINPUT51), .B1(new_n1143), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1088), .B1(new_n1148), .B2(G168), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT51), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1098), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1135), .A2(new_n1141), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(G1956), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1156), .B1(new_n1157), .B2(new_n1089), .ZN(new_n1158));
  XNOR2_X1  g733(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n1159));
  AND3_X1   g734(.A1(new_n581), .A2(new_n582), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1159), .B1(new_n581), .B2(new_n582), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(KEYINPUT56), .B(G2072), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1057), .A2(new_n1126), .A3(new_n1066), .A4(new_n1163), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1158), .A2(new_n1162), .A3(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1162), .B1(new_n1158), .B2(new_n1164), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n675), .B1(new_n1115), .B2(new_n1018), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1057), .A2(new_n810), .A3(new_n1032), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n628), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1166), .B1(new_n1170), .B2(KEYINPUT120), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT120), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1169), .A2(new_n1172), .A3(new_n628), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1165), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g749(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1175), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1167), .A2(new_n1168), .A3(KEYINPUT60), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1177), .A2(new_n837), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT60), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1169), .A2(new_n1179), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1167), .A2(new_n1168), .A3(KEYINPUT60), .A4(new_n628), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1178), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1158), .A2(new_n1164), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1162), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1158), .A2(new_n1162), .A3(new_n1164), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1185), .A2(new_n1186), .A3(KEYINPUT61), .ZN(new_n1187));
  AND3_X1   g762(.A1(new_n1176), .A2(new_n1182), .A3(new_n1187), .ZN(new_n1188));
  NOR3_X1   g763(.A1(new_n1067), .A2(new_n1071), .A3(G1996), .ZN(new_n1189));
  XNOR2_X1  g764(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1190), .B(G1341), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1033), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(new_n1192), .ZN(new_n1193));
  OAI21_X1  g768(.A(KEYINPUT122), .B1(new_n1189), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT122), .ZN(new_n1195));
  OAI211_X1 g770(.A(new_n1195), .B(new_n1192), .C1(new_n1127), .C2(G1996), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g772(.A(KEYINPUT59), .B1(new_n1197), .B2(new_n553), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT59), .ZN(new_n1199));
  AOI211_X1 g774(.A(new_n1199), .B(new_n875), .C1(new_n1194), .C2(new_n1196), .ZN(new_n1200));
  NOR2_X1   g775(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1174), .B1(new_n1188), .B2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1112), .B1(new_n1155), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1105), .A2(G286), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1152), .B1(new_n1151), .B2(new_n1204), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n1143), .A2(KEYINPUT51), .ZN(new_n1206));
  OAI21_X1  g781(.A(KEYINPUT62), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT62), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1150), .A2(new_n1208), .A3(new_n1153), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1081), .A2(new_n1055), .ZN(new_n1210));
  INV_X1    g785(.A(new_n1032), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1211), .A2(KEYINPUT50), .ZN(new_n1212));
  NAND4_X1  g787(.A1(new_n1057), .A2(new_n1212), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1213));
  OAI21_X1  g788(.A(new_n1072), .B1(new_n1213), .B2(G2090), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1078), .B1(new_n1214), .B2(G8), .ZN(new_n1215));
  NOR3_X1   g790(.A1(new_n1210), .A2(new_n1215), .A3(new_n1138), .ZN(new_n1216));
  NAND3_X1  g791(.A1(new_n1207), .A2(new_n1209), .A3(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1217), .A2(KEYINPUT125), .ZN(new_n1218));
  INV_X1    g793(.A(KEYINPUT125), .ZN(new_n1219));
  NAND4_X1  g794(.A1(new_n1207), .A2(new_n1209), .A3(new_n1216), .A4(new_n1219), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1218), .A2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g796(.A(new_n1031), .B1(new_n1203), .B2(new_n1221), .ZN(new_n1222));
  NAND4_X1  g797(.A1(new_n1027), .A2(new_n754), .A3(new_n751), .A4(new_n750), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n808), .A2(new_n810), .ZN(new_n1224));
  AOI21_X1  g799(.A(new_n1022), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g800(.A(new_n1022), .B1(new_n1010), .B2(new_n770), .ZN(new_n1226));
  OAI21_X1  g801(.A(KEYINPUT46), .B1(new_n1022), .B2(G1996), .ZN(new_n1227));
  OR3_X1    g802(.A1(new_n1022), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1228));
  AOI21_X1  g803(.A(new_n1226), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  XNOR2_X1  g804(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n1230));
  XNOR2_X1  g805(.A(new_n1229), .B(new_n1230), .ZN(new_n1231));
  NOR3_X1   g806(.A1(new_n1022), .A2(G1986), .A3(G290), .ZN(new_n1232));
  XNOR2_X1  g807(.A(new_n1232), .B(KEYINPUT48), .ZN(new_n1233));
  OAI21_X1  g808(.A(new_n1231), .B1(new_n1029), .B2(new_n1233), .ZN(new_n1234));
  NOR2_X1   g809(.A1(new_n1225), .A2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g810(.A1(new_n1222), .A2(new_n1235), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g811(.A1(G227), .A2(new_n459), .ZN(new_n1238));
  OAI21_X1  g812(.A(new_n1238), .B1(new_n678), .B2(new_n679), .ZN(new_n1239));
  NOR2_X1   g813(.A1(G229), .A2(new_n1239), .ZN(new_n1240));
  AND3_X1   g814(.A1(new_n1005), .A2(new_n1240), .A3(new_n942), .ZN(G308));
  NAND3_X1  g815(.A1(new_n1005), .A2(new_n1240), .A3(new_n942), .ZN(G225));
endmodule


