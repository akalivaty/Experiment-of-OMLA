//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 0 1 0 0 1 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 1 1 1 1 1 0 1 1 1 0 0 0 1 0 0 0 1 0 1 0 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015;
  INV_X1    g000(.A(G475), .ZN(new_n187));
  XNOR2_X1  g001(.A(G125), .B(G140), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G140), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G125), .ZN(new_n192));
  INV_X1    g006(.A(G125), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G140), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n192), .A2(new_n194), .A3(KEYINPUT74), .ZN(new_n195));
  OR3_X1    g009(.A1(new_n193), .A2(KEYINPUT74), .A3(G140), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n190), .B1(new_n197), .B2(new_n189), .ZN(new_n198));
  INV_X1    g012(.A(G237), .ZN(new_n199));
  INV_X1    g013(.A(G953), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(G214), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(G237), .A2(G953), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(G143), .A3(G214), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  AOI22_X1  g021(.A1(new_n207), .A2(KEYINPUT89), .B1(KEYINPUT18), .B2(G131), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT89), .ZN(new_n209));
  NAND2_X1  g023(.A1(KEYINPUT18), .A2(G131), .ZN(new_n210));
  NOR3_X1   g024(.A1(new_n206), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n198), .B1(new_n208), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n205), .ZN(new_n213));
  AOI21_X1  g027(.A(G143), .B1(new_n204), .B2(G214), .ZN(new_n214));
  OAI21_X1  g028(.A(G131), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT17), .ZN(new_n216));
  INV_X1    g030(.A(G131), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n203), .A2(new_n217), .A3(new_n205), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n215), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT93), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n215), .A2(KEYINPUT93), .A3(new_n216), .A4(new_n218), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n197), .A2(KEYINPUT16), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT75), .B1(new_n192), .B2(KEYINPUT16), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT75), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT16), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n226), .A2(new_n227), .A3(new_n191), .A4(G125), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n224), .A2(G146), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n227), .B1(new_n195), .B2(new_n196), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n225), .A2(new_n228), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n189), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n206), .A2(KEYINPUT17), .A3(G131), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n230), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n212), .B1(new_n223), .B2(new_n235), .ZN(new_n236));
  XOR2_X1   g050(.A(G113), .B(G122), .Z(new_n237));
  XOR2_X1   g051(.A(KEYINPUT92), .B(G104), .Z(new_n238));
  XOR2_X1   g052(.A(new_n237), .B(new_n238), .Z(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n236), .A2(new_n240), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n239), .B(new_n212), .C1(new_n223), .C2(new_n235), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G902), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n187), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n242), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n195), .A2(new_n196), .A3(KEYINPUT19), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT90), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT19), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n249), .B1(new_n188), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n195), .A2(new_n196), .A3(new_n249), .A4(KEYINPUT19), .ZN(new_n253));
  AOI21_X1  g067(.A(G146), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NOR3_X1   g068(.A1(new_n231), .A2(new_n232), .A3(new_n189), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT91), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n215), .A2(new_n218), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NOR3_X1   g072(.A1(new_n254), .A2(KEYINPUT91), .A3(new_n255), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n212), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n247), .B1(new_n260), .B2(new_n240), .ZN(new_n261));
  NOR2_X1   g075(.A1(G475), .A2(G902), .ZN(new_n262));
  XOR2_X1   g076(.A(new_n262), .B(KEYINPUT94), .Z(new_n263));
  OAI21_X1  g077(.A(KEYINPUT20), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT20), .ZN(new_n265));
  INV_X1    g079(.A(new_n263), .ZN(new_n266));
  INV_X1    g080(.A(new_n259), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(new_n257), .A3(new_n256), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n239), .B1(new_n268), .B2(new_n212), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n265), .B(new_n266), .C1(new_n269), .C2(new_n247), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n264), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT95), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n202), .A2(G128), .ZN(new_n273));
  INV_X1    g087(.A(G128), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G143), .ZN(new_n275));
  INV_X1    g089(.A(G134), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n273), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n276), .B1(new_n273), .B2(new_n275), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n272), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n273), .A2(new_n275), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G134), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(KEYINPUT95), .A3(new_n277), .ZN(new_n283));
  XOR2_X1   g097(.A(G116), .B(G122), .Z(new_n284));
  INV_X1    g098(.A(KEYINPUT14), .ZN(new_n285));
  INV_X1    g099(.A(G116), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n286), .A2(G122), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n284), .B(G107), .C1(new_n285), .C2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(G107), .B1(new_n287), .B2(new_n285), .ZN(new_n289));
  XNOR2_X1  g103(.A(G116), .B(G122), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n280), .A2(new_n283), .A3(new_n288), .A4(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT13), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n273), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n275), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n273), .A2(new_n293), .ZN(new_n296));
  OAI21_X1  g110(.A(G134), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G107), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n284), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n290), .A2(G107), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n297), .A2(new_n299), .A3(new_n300), .A4(new_n277), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT9), .B(G234), .ZN(new_n302));
  INV_X1    g116(.A(G217), .ZN(new_n303));
  NOR3_X1   g117(.A1(new_n302), .A2(new_n303), .A3(G953), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n292), .A2(new_n301), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n304), .B1(new_n292), .B2(new_n301), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n244), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT96), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G478), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n310), .A2(KEYINPUT15), .ZN(new_n311));
  OAI211_X1 g125(.A(KEYINPUT96), .B(new_n244), .C1(new_n305), .C2(new_n306), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n309), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  OR2_X1    g127(.A1(new_n307), .A2(new_n311), .ZN(new_n314));
  AND2_X1   g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n200), .A2(G952), .ZN(new_n316));
  NAND2_X1  g130(.A1(G234), .A2(G237), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  XOR2_X1   g132(.A(new_n318), .B(KEYINPUT97), .Z(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT21), .B(G898), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n317), .A2(G902), .A3(G953), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n320), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  AND4_X1   g139(.A1(new_n246), .A2(new_n271), .A3(new_n315), .A4(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(G214), .B1(G237), .B2(G902), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(G110), .B(G122), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  XOR2_X1   g144(.A(KEYINPUT2), .B(G113), .Z(new_n331));
  XNOR2_X1  g145(.A(G116), .B(G119), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G119), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G116), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n286), .A2(G119), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT2), .B(G113), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n333), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(G104), .ZN(new_n341));
  OAI21_X1  g155(.A(KEYINPUT3), .B1(new_n341), .B2(G107), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT3), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n343), .A2(new_n298), .A3(G104), .ZN(new_n344));
  INV_X1    g158(.A(G101), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n341), .A2(G107), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n342), .A2(new_n344), .A3(new_n345), .A4(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT4), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n342), .A2(new_n344), .A3(new_n346), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n345), .A2(KEYINPUT79), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n349), .A2(KEYINPUT4), .A3(new_n350), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n340), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  AND3_X1   g168(.A1(new_n335), .A2(new_n336), .A3(KEYINPUT5), .ZN(new_n355));
  OAI21_X1  g169(.A(G113), .B1(new_n335), .B2(KEYINPUT5), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n333), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n341), .A2(G107), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n298), .A2(G104), .ZN(new_n359));
  OAI21_X1  g173(.A(G101), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n347), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT81), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT81), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n347), .A2(new_n360), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n357), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n330), .B1(new_n354), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n356), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n332), .A2(KEYINPUT5), .ZN(new_n368));
  AOI22_X1  g182(.A1(new_n367), .A2(new_n368), .B1(new_n332), .B2(new_n331), .ZN(new_n369));
  AND3_X1   g183(.A1(new_n347), .A2(new_n360), .A3(new_n363), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n363), .B1(new_n347), .B2(new_n360), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n369), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n349), .A2(KEYINPUT4), .A3(new_n350), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n373), .B1(new_n351), .B2(new_n348), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n372), .B(new_n329), .C1(new_n374), .C2(new_n340), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n366), .A2(new_n375), .A3(KEYINPUT6), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT6), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n377), .B(new_n330), .C1(new_n354), .C2(new_n365), .ZN(new_n378));
  AND2_X1   g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G224), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n380), .A2(G953), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT84), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n189), .A2(G143), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n202), .A2(G146), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  AND2_X1   g200(.A1(KEYINPUT0), .A2(G128), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(KEYINPUT0), .B(G128), .ZN(new_n389));
  OAI21_X1  g203(.A(KEYINPUT64), .B1(new_n189), .B2(G143), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n383), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n189), .A2(KEYINPUT64), .A3(G143), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n389), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT65), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n388), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT64), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n396), .B1(new_n202), .B2(G146), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n202), .A2(G146), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n392), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n389), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(new_n394), .A3(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(G125), .B1(new_n395), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT1), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n383), .A2(new_n384), .A3(new_n404), .A4(G128), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT1), .B1(new_n202), .B2(G146), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G128), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n406), .B1(new_n399), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(new_n193), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n382), .B1(new_n403), .B2(new_n410), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n189), .A2(KEYINPUT64), .A3(G143), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n412), .B1(new_n383), .B2(new_n390), .ZN(new_n413));
  OAI21_X1  g227(.A(KEYINPUT65), .B1(new_n413), .B2(new_n389), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n414), .A2(new_n401), .A3(new_n388), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT84), .B1(new_n415), .B2(G125), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n381), .B1(new_n411), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n381), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n403), .A2(new_n382), .ZN(new_n419));
  INV_X1    g233(.A(new_n408), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n405), .B1(new_n413), .B2(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n421), .A2(G125), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n422), .B1(G125), .B2(new_n415), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n418), .B(new_n419), .C1(new_n423), .C2(new_n382), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n417), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(G902), .B1(new_n379), .B2(new_n425), .ZN(new_n426));
  XOR2_X1   g240(.A(KEYINPUT86), .B(KEYINPUT7), .Z(new_n427));
  OAI22_X1  g241(.A1(new_n411), .A2(new_n416), .B1(new_n381), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT87), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI221_X1 g244(.A(KEYINPUT87), .B1(new_n381), .B2(new_n427), .C1(new_n411), .C2(new_n416), .ZN(new_n431));
  INV_X1    g245(.A(new_n411), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n432), .A2(KEYINPUT7), .A3(new_n418), .A4(new_n419), .ZN(new_n433));
  INV_X1    g247(.A(new_n375), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT85), .ZN(new_n435));
  INV_X1    g249(.A(new_n361), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n435), .B1(new_n369), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n357), .A2(KEYINPUT85), .A3(new_n361), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n437), .A2(new_n372), .A3(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n329), .B(KEYINPUT8), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n434), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n430), .A2(new_n431), .A3(new_n433), .A4(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n426), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(G210), .B1(G237), .B2(G902), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n444), .B(KEYINPUT88), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n445), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n426), .A2(new_n442), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n328), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(G221), .ZN(new_n450));
  INV_X1    g264(.A(new_n302), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n450), .B1(new_n451), .B2(new_n244), .ZN(new_n452));
  XNOR2_X1  g266(.A(KEYINPUT82), .B(G469), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n352), .A2(new_n353), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n399), .A2(new_n400), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n455), .A2(KEYINPUT65), .B1(new_n387), .B2(new_n386), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n454), .A2(new_n456), .A3(new_n401), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT11), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n458), .B1(new_n276), .B2(G137), .ZN(new_n459));
  INV_X1    g273(.A(G137), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(KEYINPUT11), .A3(G134), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n276), .A2(G137), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n459), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(G131), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n459), .A2(new_n461), .A3(new_n217), .A4(new_n462), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n421), .B(KEYINPUT10), .C1(new_n370), .C2(new_n371), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT10), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT80), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n407), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n383), .A2(KEYINPUT80), .A3(KEYINPUT1), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(G128), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n406), .B1(new_n473), .B2(new_n385), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n469), .B1(new_n474), .B2(new_n361), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n457), .A2(new_n467), .A3(new_n468), .A4(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(G110), .B(G140), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n200), .A2(G227), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n477), .B(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n409), .A2(new_n362), .A3(new_n364), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n404), .B1(G143), .B2(new_n189), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n274), .B1(new_n481), .B2(KEYINPUT80), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n386), .B1(new_n482), .B2(new_n471), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n436), .B1(new_n483), .B2(new_n406), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(KEYINPUT12), .B1(new_n485), .B2(new_n466), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT12), .ZN(new_n487));
  AOI211_X1 g301(.A(new_n487), .B(new_n467), .C1(new_n480), .C2(new_n484), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n476), .B(new_n479), .C1(new_n486), .C2(new_n488), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n475), .B(new_n468), .C1(new_n415), .C2(new_n374), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n466), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n479), .B1(new_n491), .B2(new_n476), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT83), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n489), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AOI211_X1 g308(.A(KEYINPUT83), .B(new_n479), .C1(new_n491), .C2(new_n476), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n244), .B(new_n453), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n476), .B1(new_n486), .B2(new_n488), .ZN(new_n497));
  XOR2_X1   g311(.A(new_n479), .B(KEYINPUT78), .Z(new_n498));
  AND2_X1   g312(.A1(new_n476), .A2(new_n479), .ZN(new_n499));
  AOI22_X1  g313(.A1(new_n497), .A2(new_n498), .B1(new_n499), .B2(new_n491), .ZN(new_n500));
  OAI21_X1  g314(.A(G469), .B1(new_n500), .B2(G902), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n452), .B1(new_n496), .B2(new_n501), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n326), .A2(new_n449), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n340), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n414), .A2(new_n466), .A3(new_n401), .A4(new_n388), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT68), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT68), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n456), .A2(new_n507), .A3(new_n466), .A4(new_n401), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT66), .ZN(new_n509));
  XNOR2_X1  g323(.A(G134), .B(G137), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n509), .B1(new_n510), .B2(new_n217), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n276), .A2(G137), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n460), .A2(G134), .ZN(new_n513));
  OAI211_X1 g327(.A(KEYINPUT66), .B(G131), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n511), .A2(new_n465), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n421), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n506), .A2(new_n508), .A3(KEYINPUT30), .A4(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n505), .A2(new_n516), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT30), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT67), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT67), .ZN(new_n521));
  AOI211_X1 g335(.A(new_n521), .B(KEYINPUT30), .C1(new_n505), .C2(new_n516), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n504), .B(new_n517), .C1(new_n520), .C2(new_n522), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n506), .A2(new_n508), .A3(new_n340), .A4(new_n516), .ZN(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT26), .B(G101), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n204), .A2(G210), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n525), .B(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n528));
  XOR2_X1   g342(.A(new_n527), .B(new_n528), .Z(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n523), .A2(new_n524), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT28), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n532), .B1(new_n518), .B2(new_n504), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n518), .A2(new_n504), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT70), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n340), .B1(new_n505), .B2(new_n516), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT70), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n536), .A2(new_n524), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n534), .B1(new_n540), .B2(KEYINPUT28), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n531), .B1(new_n541), .B2(new_n530), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT29), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT71), .ZN(new_n545));
  OR2_X1    g359(.A1(new_n524), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n506), .A2(new_n508), .A3(new_n516), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n504), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n524), .A2(new_n545), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n546), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(KEYINPUT28), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n551), .A2(KEYINPUT29), .A3(new_n533), .A4(new_n529), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n544), .A2(new_n244), .A3(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(G472), .ZN(new_n554));
  NOR2_X1   g368(.A1(G472), .A2(G902), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT31), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n524), .A2(new_n529), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n523), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n557), .B1(new_n523), .B2(new_n558), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n537), .B(KEYINPUT70), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n532), .B1(new_n562), .B2(new_n524), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n530), .B1(new_n563), .B2(new_n534), .ZN(new_n564));
  AOI211_X1 g378(.A(KEYINPUT32), .B(new_n556), .C1(new_n561), .C2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT32), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n523), .A2(new_n558), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(KEYINPUT31), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n523), .A2(new_n557), .A3(new_n558), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n568), .B(new_n569), .C1(new_n541), .C2(new_n529), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n566), .B1(new_n570), .B2(new_n555), .ZN(new_n571));
  OAI22_X1  g385(.A1(new_n553), .A2(new_n554), .B1(new_n565), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT73), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n573), .B1(new_n334), .B2(G128), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n334), .A2(G128), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(KEYINPUT23), .A3(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(KEYINPUT23), .B1(new_n274), .B2(G119), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n274), .A2(G119), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(new_n573), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(G110), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n575), .A2(new_n578), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT72), .ZN(new_n583));
  INV_X1    g397(.A(G110), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(KEYINPUT24), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT24), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(G110), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n583), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n585), .A2(new_n587), .A3(new_n583), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n582), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n230), .B(new_n190), .C1(new_n581), .C2(new_n591), .ZN(new_n592));
  AND3_X1   g406(.A1(new_n585), .A2(new_n587), .A3(new_n583), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n593), .A2(new_n588), .ZN(new_n594));
  AOI22_X1  g408(.A1(new_n594), .A2(new_n582), .B1(new_n580), .B2(G110), .ZN(new_n595));
  AOI21_X1  g409(.A(G146), .B1(new_n224), .B2(new_n229), .ZN(new_n596));
  OAI211_X1 g410(.A(KEYINPUT76), .B(new_n595), .C1(new_n596), .C2(new_n255), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n230), .A2(new_n233), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT76), .B1(new_n599), .B2(new_n595), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n592), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT22), .B(G137), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n200), .A2(G221), .A3(G234), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n604), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n592), .B(new_n606), .C1(new_n598), .C2(new_n600), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n605), .A2(new_n244), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT25), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n605), .A2(KEYINPUT25), .A3(new_n244), .A4(new_n607), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n303), .B1(G234), .B2(new_n244), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n605), .A2(new_n607), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(KEYINPUT77), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT77), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n605), .A2(new_n616), .A3(new_n607), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n613), .A2(G902), .ZN(new_n619));
  AOI22_X1  g433(.A1(new_n612), .A2(new_n613), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n503), .A2(new_n572), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G101), .ZN(G3));
  NAND2_X1  g436(.A1(new_n449), .A2(new_n325), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n568), .A2(new_n569), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n541), .A2(new_n529), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n555), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(G902), .B1(new_n561), .B2(new_n564), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n626), .B1(new_n627), .B2(new_n554), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n620), .A2(new_n502), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n623), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n271), .A2(new_n246), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n309), .A2(new_n310), .A3(new_n312), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n310), .A2(G902), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n305), .A2(new_n306), .A3(KEYINPUT33), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT33), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n292), .A2(new_n301), .ZN(new_n636));
  INV_X1    g450(.A(new_n304), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n292), .A2(new_n301), .A3(new_n304), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n635), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OAI211_X1 g454(.A(KEYINPUT98), .B(new_n633), .C1(new_n634), .C2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n632), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(KEYINPUT33), .B1(new_n305), .B2(new_n306), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n638), .A2(new_n635), .A3(new_n639), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(KEYINPUT98), .B1(new_n645), .B2(new_n633), .ZN(new_n646));
  OAI21_X1  g460(.A(KEYINPUT99), .B1(new_n642), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n645), .A2(new_n633), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT98), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT99), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n650), .A2(new_n651), .A3(new_n632), .A4(new_n641), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n630), .A2(new_n631), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT34), .B(G104), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G6));
  INV_X1    g470(.A(KEYINPUT100), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n271), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n264), .A2(KEYINPUT100), .A3(new_n270), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n315), .A2(new_n245), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n630), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT35), .B(G107), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G9));
  NOR2_X1   g479(.A1(new_n604), .A2(KEYINPUT36), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n601), .B(new_n666), .ZN(new_n667));
  AOI22_X1  g481(.A1(new_n612), .A2(new_n613), .B1(new_n667), .B2(new_n619), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n628), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n503), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT37), .B(G110), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT101), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n670), .B(new_n672), .ZN(G12));
  INV_X1    g487(.A(new_n502), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n426), .A2(new_n442), .A3(new_n447), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n447), .B1(new_n426), .B2(new_n442), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n327), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n674), .A2(new_n677), .A3(new_n668), .ZN(new_n678));
  INV_X1    g492(.A(G900), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n320), .B1(new_n679), .B2(new_n323), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n661), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n572), .A2(new_n678), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(KEYINPUT102), .B(G128), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G30));
  AND2_X1   g498(.A1(new_n523), .A2(new_n524), .ZN(new_n685));
  OR2_X1    g499(.A1(new_n685), .A2(new_n530), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n244), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n550), .A2(new_n529), .ZN(new_n688));
  OAI21_X1  g502(.A(G472), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n689), .B1(new_n565), .B2(new_n571), .ZN(new_n690));
  XOR2_X1   g504(.A(new_n690), .B(KEYINPUT104), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n680), .B(KEYINPUT39), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n674), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n693), .A2(new_n694), .ZN(new_n696));
  INV_X1    g510(.A(new_n668), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n315), .B1(new_n271), .B2(new_n246), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n697), .A2(new_n699), .A3(new_n328), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n446), .A2(new_n448), .ZN(new_n701));
  XOR2_X1   g515(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n696), .A2(new_n700), .A3(new_n703), .ZN(new_n704));
  OR3_X1    g518(.A1(new_n691), .A2(new_n695), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G143), .ZN(G45));
  INV_X1    g520(.A(new_n680), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n653), .A2(new_n631), .A3(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n572), .A2(new_n678), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G146), .ZN(G48));
  INV_X1    g525(.A(new_n620), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n626), .A2(KEYINPUT32), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n570), .A2(new_n566), .A3(new_n555), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n544), .A2(new_n244), .A3(new_n552), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(G472), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n712), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n244), .B1(new_n494), .B2(new_n495), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(G469), .ZN(new_n720));
  INV_X1    g534(.A(new_n452), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n720), .A2(new_n721), .A3(new_n496), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(KEYINPUT106), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n653), .A2(new_n631), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n623), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n718), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT41), .B(G113), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G15));
  NOR2_X1   g542(.A1(new_n623), .A2(new_n661), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n718), .A2(new_n723), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G116), .ZN(G18));
  NOR3_X1   g545(.A1(new_n722), .A2(new_n677), .A3(new_n668), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n572), .A2(new_n732), .A3(new_n326), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G119), .ZN(G21));
  NAND2_X1  g548(.A1(new_n551), .A2(new_n533), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n530), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n556), .B1(new_n736), .B2(new_n561), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT107), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n738), .B1(new_n627), .B2(new_n554), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n570), .A2(new_n244), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(KEYINPUT107), .A3(G472), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n737), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n623), .A2(new_n699), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n723), .A2(new_n742), .A3(new_n743), .A4(new_n620), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G122), .ZN(G24));
  NAND2_X1  g559(.A1(new_n739), .A2(new_n741), .ZN(new_n746));
  INV_X1    g560(.A(new_n737), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n732), .A2(new_n746), .A3(new_n709), .A4(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G125), .ZN(G27));
  NAND4_X1  g563(.A1(new_n502), .A2(new_n327), .A3(new_n446), .A4(new_n448), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n572), .A2(new_n620), .A3(new_n751), .A4(new_n709), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT42), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT108), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n755), .B1(new_n565), .B2(new_n571), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n713), .A2(KEYINPUT108), .A3(new_n714), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n757), .A3(new_n717), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n750), .A2(new_n753), .A3(new_n708), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(new_n620), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n754), .A2(new_n760), .ZN(new_n761));
  XOR2_X1   g575(.A(KEYINPUT109), .B(G131), .Z(new_n762));
  XNOR2_X1  g576(.A(new_n761), .B(new_n762), .ZN(G33));
  AND4_X1   g577(.A1(new_n572), .A2(new_n620), .A3(new_n681), .A4(new_n751), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(new_n276), .ZN(G36));
  AOI21_X1  g579(.A(new_n245), .B1(new_n264), .B2(new_n270), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n653), .A2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT43), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n769), .A2(new_n628), .A3(new_n697), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT44), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(KEYINPUT111), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT46), .ZN(new_n774));
  OAI21_X1  g588(.A(G469), .B1(new_n500), .B2(KEYINPUT45), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n500), .A2(KEYINPUT45), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n776), .A2(KEYINPUT110), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(KEYINPUT110), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n775), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(G469), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(new_n244), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n774), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n496), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n779), .A2(new_n774), .A3(new_n781), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n721), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(new_n692), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n446), .A2(new_n327), .A3(new_n448), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n788), .B1(new_n770), .B2(new_n771), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n773), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G137), .ZN(G39));
  INV_X1    g605(.A(KEYINPUT47), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n786), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n785), .A2(KEYINPUT47), .A3(new_n721), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR4_X1   g609(.A1(new_n572), .A2(new_n620), .A3(new_n708), .A4(new_n788), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G140), .ZN(G42));
  AOI22_X1  g612(.A1(new_n715), .A2(new_n755), .B1(G472), .B2(new_n716), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n712), .B1(new_n799), .B2(new_n757), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n722), .A2(new_n788), .A3(new_n319), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n769), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  XOR2_X1   g617(.A(new_n803), .B(KEYINPUT48), .Z(new_n804));
  AND2_X1   g618(.A1(new_n720), .A2(new_n496), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n721), .A3(new_n449), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n769), .A2(new_n320), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n742), .A2(new_n620), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n801), .A2(new_n620), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n691), .A2(new_n810), .ZN(new_n811));
  OAI221_X1 g625(.A(new_n316), .B1(new_n806), .B2(new_n809), .C1(new_n811), .C2(new_n724), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n811), .A2(new_n631), .A3(new_n653), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n742), .A2(new_n697), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n813), .B1(new_n802), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n809), .A2(new_n788), .ZN(new_n816));
  INV_X1    g630(.A(new_n805), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n817), .A2(new_n721), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n816), .B1(new_n795), .B2(new_n818), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n703), .A2(new_n327), .A3(new_n722), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n807), .A2(new_n808), .A3(new_n820), .ZN(new_n821));
  XOR2_X1   g635(.A(new_n821), .B(KEYINPUT50), .Z(new_n822));
  NAND3_X1  g636(.A1(new_n815), .A2(new_n819), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT51), .ZN(new_n824));
  AOI211_X1 g638(.A(new_n804), .B(new_n812), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n748), .A2(new_n682), .ZN(new_n826));
  AOI22_X1  g640(.A1(new_n713), .A2(new_n714), .B1(new_n716), .B2(G472), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n697), .A2(new_n502), .A3(new_n449), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n674), .B1(new_n715), .B2(new_n689), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n701), .A2(new_n698), .A3(new_n327), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n612), .A2(new_n613), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n667), .A2(new_n619), .ZN(new_n833));
  XOR2_X1   g647(.A(new_n680), .B(KEYINPUT114), .Z(new_n834));
  NAND3_X1  g648(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT115), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n668), .A2(KEYINPUT115), .A3(new_n834), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n831), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI22_X1  g653(.A1(new_n829), .A2(new_n709), .B1(new_n830), .B2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n826), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n837), .A2(new_n838), .ZN(new_n843));
  INV_X1    g657(.A(new_n831), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n843), .A2(new_n502), .A3(new_n690), .A4(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n845), .A2(new_n748), .A3(new_n682), .A4(new_n710), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT116), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n842), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT52), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n750), .A2(new_n668), .ZN(new_n851));
  AOI211_X1 g665(.A(new_n737), .B(new_n708), .C1(new_n739), .C2(new_n741), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n315), .A2(new_n246), .A3(new_n707), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n658), .A2(new_n853), .A3(new_n659), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n827), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n851), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n764), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT113), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n724), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n653), .A2(new_n631), .A3(KEYINPUT113), .ZN(new_n860));
  OR2_X1    g674(.A1(new_n631), .A2(new_n315), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n628), .A2(new_n629), .ZN(new_n863));
  INV_X1    g677(.A(new_n623), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n503), .B1(new_n718), .B2(new_n669), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n856), .A2(new_n857), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  AOI22_X1  g681(.A1(new_n800), .A2(new_n759), .B1(new_n753), .B2(new_n752), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n726), .A2(new_n744), .A3(new_n730), .A4(new_n733), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n842), .A2(new_n847), .A3(KEYINPUT52), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n850), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(KEYINPUT53), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n849), .B1(new_n826), .B2(new_n840), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n874), .B1(new_n848), .B2(new_n849), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT53), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n875), .A2(new_n876), .A3(new_n870), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n873), .A2(new_n877), .A3(KEYINPUT54), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n868), .A2(new_n869), .ZN(new_n879));
  INV_X1    g693(.A(new_n867), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n871), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT52), .B1(new_n842), .B2(new_n847), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n876), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT54), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n865), .A2(new_n621), .A3(new_n670), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n885), .A2(KEYINPUT53), .A3(new_n857), .A4(new_n856), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT117), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n886), .B1(new_n879), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(KEYINPUT117), .B1(new_n868), .B2(new_n869), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n875), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n883), .A2(new_n884), .A3(new_n890), .ZN(new_n891));
  OR2_X1    g705(.A1(new_n823), .A2(new_n824), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n825), .A2(new_n878), .A3(new_n891), .A4(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n893), .B1(G952), .B2(G953), .ZN(new_n894));
  OR4_X1    g708(.A1(new_n712), .A2(new_n767), .A3(new_n452), .A4(new_n328), .ZN(new_n895));
  AOI211_X1 g709(.A(new_n703), .B(new_n895), .C1(KEYINPUT49), .C2(new_n817), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n817), .A2(KEYINPUT49), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT112), .Z(new_n898));
  NAND3_X1  g712(.A1(new_n896), .A2(new_n691), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n894), .A2(new_n899), .ZN(G75));
  AND3_X1   g714(.A1(new_n744), .A2(new_n726), .A3(new_n733), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n901), .A2(new_n887), .A3(new_n761), .A4(new_n730), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n866), .A2(new_n865), .ZN(new_n903));
  INV_X1    g717(.A(new_n851), .ZN(new_n904));
  INV_X1    g718(.A(new_n854), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n572), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n746), .A2(new_n709), .A3(new_n747), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NOR4_X1   g722(.A1(new_n903), .A2(new_n908), .A3(new_n876), .A4(new_n764), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n889), .A2(new_n902), .A3(new_n909), .ZN(new_n910));
  AOI22_X1  g724(.A1(new_n872), .A2(new_n876), .B1(new_n910), .B2(new_n875), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n911), .A2(new_n244), .A3(new_n447), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n912), .A2(KEYINPUT56), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n379), .B(KEYINPUT118), .Z(new_n914));
  XOR2_X1   g728(.A(new_n425), .B(KEYINPUT55), .Z(new_n915));
  XNOR2_X1  g729(.A(new_n914), .B(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n200), .A2(G952), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  XNOR2_X1  g733(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n919), .B1(new_n912), .B2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n917), .A2(new_n922), .ZN(G51));
  XNOR2_X1  g737(.A(new_n781), .B(KEYINPUT57), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT120), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n883), .A2(new_n890), .A3(new_n925), .A4(new_n884), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n926), .B1(new_n884), .B2(new_n911), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n925), .B1(new_n911), .B2(new_n884), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n924), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  OR2_X1    g743(.A1(new_n494), .A2(new_n495), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n244), .B1(new_n883), .B2(new_n890), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n779), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT121), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n918), .B1(new_n931), .B2(new_n935), .ZN(G54));
  INV_X1    g750(.A(new_n261), .ZN(new_n937));
  AND2_X1   g751(.A1(KEYINPUT58), .A2(G475), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n932), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n937), .B1(new_n932), .B2(new_n938), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n939), .A2(new_n940), .A3(new_n918), .ZN(G60));
  NAND2_X1  g755(.A1(G478), .A2(G902), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT59), .Z(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(new_n878), .B2(new_n891), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n919), .B1(new_n944), .B2(new_n645), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n943), .B1(new_n643), .B2(new_n644), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n946), .B1(new_n927), .B2(new_n928), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(KEYINPUT122), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT122), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n949), .B(new_n946), .C1(new_n927), .C2(new_n928), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n945), .B1(new_n948), .B2(new_n950), .ZN(G63));
  XNOR2_X1  g765(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(G217), .A2(G902), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT60), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n911), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n667), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n919), .B1(new_n956), .B2(new_n618), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n953), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OR2_X1    g774(.A1(new_n956), .A2(new_n618), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n961), .A2(new_n919), .A3(new_n957), .A4(new_n952), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n960), .A2(new_n962), .ZN(G66));
  OAI21_X1  g777(.A(G953), .B1(new_n321), .B2(new_n380), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n869), .A2(new_n903), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n964), .B1(new_n965), .B2(G953), .ZN(new_n966));
  INV_X1    g780(.A(new_n914), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(G898), .B2(new_n200), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n966), .B(new_n968), .ZN(G69));
  AND2_X1   g783(.A1(new_n790), .A2(new_n797), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n826), .A2(new_n710), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT125), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n800), .A2(new_n844), .ZN(new_n974));
  AOI211_X1 g788(.A(new_n764), .B(new_n868), .C1(new_n787), .C2(new_n974), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n970), .A2(new_n200), .A3(new_n973), .A4(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n517), .B1(new_n520), .B2(new_n522), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n252), .A2(new_n253), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n977), .B(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n979), .B1(G900), .B2(G953), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT126), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n200), .B1(G227), .B2(G900), .ZN(new_n982));
  AOI22_X1  g796(.A1(new_n976), .A2(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n982), .A2(new_n981), .ZN(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n973), .A2(new_n705), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(KEYINPUT62), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT62), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n973), .A2(new_n988), .A3(new_n705), .ZN(new_n989));
  INV_X1    g803(.A(new_n862), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n990), .A2(new_n692), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n991), .A2(new_n718), .A3(new_n751), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n987), .A2(new_n970), .A3(new_n989), .A4(new_n992), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n993), .A2(new_n200), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n979), .B(KEYINPUT124), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n983), .B(new_n985), .C1(new_n994), .C2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n976), .A2(new_n980), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n982), .A2(new_n981), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n995), .B1(new_n993), .B2(new_n200), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n984), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  AND2_X1   g815(.A1(new_n996), .A2(new_n1001), .ZN(G72));
  NAND2_X1  g816(.A1(G472), .A2(G902), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1003), .B(KEYINPUT63), .Z(new_n1004));
  XNOR2_X1  g818(.A(new_n1004), .B(KEYINPUT127), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n970), .A2(new_n973), .A3(new_n975), .ZN(new_n1006));
  INV_X1    g820(.A(new_n965), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(new_n531), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n918), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1005), .B1(new_n993), .B2(new_n1007), .ZN(new_n1011));
  INV_X1    g825(.A(new_n686), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  AND2_X1   g827(.A1(new_n531), .A2(new_n1004), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n873), .A2(new_n686), .A3(new_n877), .A4(new_n1014), .ZN(new_n1015));
  AND3_X1   g829(.A1(new_n1010), .A2(new_n1013), .A3(new_n1015), .ZN(G57));
endmodule


