//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 0 1 0 0 1 0 1 0 1 0 1 0 1 0 0 0 1 0 1 0 1 0 0 0 1 1 0 0 0 0 0 1 1 0 0 1 0 0 1 0 0 0 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1288, new_n1289, new_n1290, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI211_X1 g0005(.A(G50), .B(G77), .C1(new_n204), .C2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n204), .A2(new_n205), .ZN(new_n215));
  INV_X1    g0015(.A(G50), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n209), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT65), .Z(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n211), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n214), .B(new_n220), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G226), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  NAND2_X1  g0045(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT8), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G58), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n208), .A2(G20), .ZN(new_n250));
  AND2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n252));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n218), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(KEYINPUT68), .ZN(new_n255));
  AND2_X1   g0055(.A1(new_n253), .A2(new_n218), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT68), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g0058(.A1(new_n251), .A2(new_n252), .A3(new_n255), .A4(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n259), .B1(new_n252), .B2(new_n249), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT76), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n259), .B(KEYINPUT76), .C1(new_n252), .C2(new_n249), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g0064(.A(KEYINPUT3), .B(G33), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT7), .ZN(new_n266));
  NOR3_X1   g0066(.A1(new_n265), .A2(new_n266), .A3(G20), .ZN(new_n267));
  INV_X1    g0067(.A(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT3), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT3), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(KEYINPUT7), .B1(new_n272), .B2(new_n209), .ZN(new_n273));
  OAI21_X1  g0073(.A(G68), .B1(new_n267), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n209), .A2(new_n268), .A3(G159), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT73), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G20), .A2(G33), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT73), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(new_n278), .A3(G159), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G58), .A2(G68), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n204), .A2(new_n205), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n280), .B1(G20), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n274), .A2(new_n283), .A3(KEYINPUT16), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT74), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n266), .B1(new_n265), .B2(G20), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n272), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n203), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n282), .A2(G20), .ZN(new_n290));
  INV_X1    g0090(.A(G159), .ZN(new_n291));
  NOR4_X1   g0091(.A1(new_n291), .A2(KEYINPUT73), .A3(G20), .A4(G33), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n278), .B1(new_n277), .B2(G159), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n290), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n289), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n296), .A2(KEYINPUT74), .A3(KEYINPUT16), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n286), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n272), .A2(new_n209), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT75), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n300), .B1(new_n268), .B2(KEYINPUT3), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n270), .A2(KEYINPUT75), .A3(G33), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n301), .A2(new_n269), .A3(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n266), .A2(G20), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n299), .A2(new_n266), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n283), .B1(new_n305), .B2(new_n203), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT16), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n256), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n264), .B1(new_n298), .B2(new_n308), .ZN(new_n309));
  AND2_X1   g0109(.A1(G1), .A2(G13), .ZN(new_n310));
  NAND2_X1  g0110(.A1(G33), .A2(G41), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G41), .ZN(new_n313));
  INV_X1    g0113(.A(G45), .ZN(new_n314));
  AOI21_X1  g0114(.A(G1), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n312), .A2(G274), .A3(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G232), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n316), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G226), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G1698), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(G223), .B2(G1698), .ZN(new_n323));
  INV_X1    g0123(.A(G87), .ZN(new_n324));
  OAI22_X1  g0124(.A1(new_n323), .A2(new_n272), .B1(new_n268), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n312), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n320), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G179), .ZN(new_n328));
  INV_X1    g0128(.A(G169), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n328), .B1(new_n329), .B2(new_n327), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(KEYINPUT18), .B1(new_n309), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(KEYINPUT74), .B1(new_n296), .B2(KEYINPUT16), .ZN(new_n333));
  NOR4_X1   g0133(.A1(new_n289), .A2(new_n295), .A3(new_n285), .A4(new_n307), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n308), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n262), .A2(new_n263), .ZN(new_n336));
  INV_X1    g0136(.A(G190), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n327), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(G200), .B2(new_n327), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n335), .A2(new_n336), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT17), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n309), .A2(KEYINPUT17), .A3(new_n339), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT18), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n303), .A2(new_n304), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n203), .B1(new_n345), .B2(new_n287), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n307), .B1(new_n346), .B2(new_n295), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n254), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n348), .B1(new_n286), .B2(new_n297), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n344), .B(new_n330), .C1(new_n349), .C2(new_n264), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n332), .A2(new_n342), .A3(new_n343), .A4(new_n350), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n351), .A2(KEYINPUT77), .ZN(new_n352));
  INV_X1    g0152(.A(new_n252), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n203), .ZN(new_n354));
  XNOR2_X1  g0154(.A(new_n354), .B(KEYINPUT12), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n258), .A2(new_n255), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n277), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n357));
  INV_X1    g0157(.A(G77), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n209), .A2(G33), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n356), .A2(KEYINPUT11), .A3(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n353), .A2(new_n254), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n362), .A2(G68), .A3(new_n250), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n355), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(KEYINPUT11), .B1(new_n356), .B2(new_n360), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(G1698), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n321), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n319), .A2(G1698), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n269), .A2(new_n368), .A3(new_n271), .A4(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G33), .A2(G97), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n326), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT13), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n313), .A2(new_n314), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n208), .A2(new_n375), .B1(new_n310), .B2(new_n311), .ZN(new_n376));
  INV_X1    g0176(.A(G274), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n377), .B1(new_n310), .B2(new_n311), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n376), .A2(G238), .B1(new_n378), .B2(new_n315), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n373), .A2(new_n374), .A3(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(G238), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n316), .B1(new_n318), .B2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n312), .B1(new_n370), .B2(new_n371), .ZN(new_n383));
  OAI21_X1  g0183(.A(KEYINPUT13), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n366), .B1(new_n337), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n385), .ZN(new_n387));
  INV_X1    g0187(.A(G200), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n385), .A2(G169), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n391), .A2(KEYINPUT72), .A3(KEYINPUT14), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT72), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n329), .B1(new_n380), .B2(new_n384), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT14), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n394), .A2(new_n395), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n387), .A2(G179), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n392), .A2(new_n396), .A3(new_n397), .A4(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n366), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n390), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n272), .A2(G1698), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(G222), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n272), .A2(G77), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(G223), .ZN(new_n406));
  OAI21_X1  g0206(.A(KEYINPUT67), .B1(new_n272), .B2(new_n367), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT67), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n265), .A2(new_n408), .A3(G1698), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n406), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n326), .B1(new_n405), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n316), .B1(new_n318), .B2(new_n321), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(G190), .A3(new_n413), .ZN(new_n414));
  NOR3_X1   g0214(.A1(new_n272), .A2(KEYINPUT67), .A3(new_n367), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n408), .B1(new_n265), .B2(G1698), .ZN(new_n416));
  OAI21_X1  g0216(.A(G223), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n402), .A2(G222), .B1(G77), .B2(new_n272), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n312), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(G200), .B1(new_n419), .B2(new_n412), .ZN(new_n420));
  XNOR2_X1  g0220(.A(new_n254), .B(new_n257), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n421), .A2(G50), .A3(new_n252), .A4(new_n250), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n209), .B1(new_n215), .B2(new_n216), .ZN(new_n423));
  XNOR2_X1  g0223(.A(KEYINPUT8), .B(G58), .ZN(new_n424));
  INV_X1    g0224(.A(G150), .ZN(new_n425));
  INV_X1    g0225(.A(new_n277), .ZN(new_n426));
  OAI22_X1  g0226(.A1(new_n424), .A2(new_n359), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n356), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n353), .A2(new_n216), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n422), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n430), .A2(KEYINPUT9), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n430), .A2(KEYINPUT9), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n414), .B(new_n420), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n420), .A2(KEYINPUT71), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n433), .A2(KEYINPUT10), .A3(new_n434), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n420), .A2(new_n414), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n388), .B1(new_n411), .B2(new_n413), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT71), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT10), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n436), .B(new_n439), .C1(new_n431), .C2(new_n432), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n435), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(G169), .B1(new_n411), .B2(new_n413), .ZN(new_n442));
  INV_X1    g0242(.A(new_n430), .ZN(new_n443));
  OR3_X1    g0243(.A1(new_n442), .A2(KEYINPUT69), .A3(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(KEYINPUT69), .B1(new_n442), .B2(new_n443), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n411), .A2(new_n413), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n444), .B(new_n445), .C1(G179), .C2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(G238), .B1(new_n415), .B2(new_n416), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n402), .A2(G232), .B1(G107), .B2(new_n272), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n312), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(G244), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n316), .B1(new_n318), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n329), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  OAI22_X1  g0253(.A1(new_n424), .A2(new_n426), .B1(new_n209), .B2(new_n358), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT70), .ZN(new_n455));
  XNOR2_X1  g0255(.A(KEYINPUT15), .B(G87), .ZN(new_n456));
  OAI22_X1  g0256(.A1(new_n454), .A2(new_n455), .B1(new_n359), .B2(new_n456), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n249), .A2(new_n277), .B1(G20), .B2(G77), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(KEYINPUT70), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n254), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n358), .B1(new_n208), .B2(G20), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n362), .A2(new_n461), .B1(new_n358), .B2(new_n353), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n453), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n450), .A2(new_n452), .ZN(new_n465));
  INV_X1    g0265(.A(G179), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n463), .B1(new_n465), .B2(G190), .ZN(new_n469));
  OAI21_X1  g0269(.A(G200), .B1(new_n450), .B2(new_n452), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AND2_X1   g0271(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  AND4_X1   g0272(.A1(new_n401), .A2(new_n441), .A3(new_n447), .A4(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n351), .A2(KEYINPUT77), .ZN(new_n474));
  AND3_X1   g0274(.A1(new_n352), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G116), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n477), .B1(new_n208), .B2(G33), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(KEYINPUT82), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT82), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G116), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n479), .A2(new_n481), .A3(G20), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G13), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(G1), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n362), .A2(new_n478), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G33), .A2(G283), .ZN(new_n487));
  INV_X1    g0287(.A(G97), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n487), .B(new_n209), .C1(G33), .C2(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(KEYINPUT86), .A2(KEYINPUT20), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n482), .A2(new_n254), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n482), .A2(new_n254), .A3(new_n489), .ZN(new_n492));
  XOR2_X1   g0292(.A(KEYINPUT86), .B(KEYINPUT20), .Z(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n486), .A2(new_n491), .A3(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n269), .A2(new_n271), .A3(G257), .A4(new_n367), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n269), .A2(new_n271), .A3(G264), .A4(G1698), .ZN(new_n498));
  INV_X1    g0298(.A(G303), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n497), .B(new_n498), .C1(new_n499), .C2(new_n265), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n326), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT5), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT81), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n502), .B1(new_n503), .B2(G41), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n314), .A2(G1), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n313), .A2(KEYINPUT81), .A3(KEYINPUT5), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n507), .A2(G270), .A3(new_n312), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n378), .A2(new_n504), .A3(new_n505), .A4(new_n506), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT85), .ZN(new_n510));
  AND3_X1   g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n510), .B1(new_n508), .B2(new_n509), .ZN(new_n512));
  OAI211_X1 g0312(.A(G190), .B(new_n501), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n508), .A2(new_n509), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT85), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n515), .A2(new_n516), .B1(new_n326), .B2(new_n500), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n496), .B(new_n513), .C1(new_n517), .C2(new_n388), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT21), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n495), .A2(G169), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n519), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n517), .A2(G179), .A3(new_n495), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n501), .B1(new_n511), .B2(new_n512), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n523), .A2(KEYINPUT21), .A3(G169), .A4(new_n495), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n518), .A2(new_n521), .A3(new_n522), .A4(new_n524), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n269), .A2(new_n271), .A3(new_n209), .A4(G87), .ZN(new_n526));
  NAND2_X1  g0326(.A1(KEYINPUT87), .A2(KEYINPUT22), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n265), .A2(new_n209), .A3(G87), .A4(new_n527), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT24), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n268), .B1(new_n479), .B2(new_n481), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT23), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n209), .B2(G107), .ZN(new_n535));
  INV_X1    g0335(.A(G107), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n536), .A2(KEYINPUT23), .A3(G20), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n533), .A2(new_n209), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n531), .A2(new_n532), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n532), .B1(new_n531), .B2(new_n538), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n254), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  XOR2_X1   g0342(.A(KEYINPUT88), .B(KEYINPUT25), .Z(new_n543));
  NOR2_X1   g0343(.A1(new_n252), .A2(G107), .ZN(new_n544));
  XNOR2_X1  g0344(.A(new_n543), .B(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n208), .A2(G33), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n421), .A2(new_n252), .A3(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n545), .B1(new_n547), .B2(new_n536), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n507), .A2(G264), .A3(new_n312), .ZN(new_n550));
  INV_X1    g0350(.A(G294), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n268), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(G250), .A2(G1698), .ZN(new_n553));
  INV_X1    g0353(.A(G257), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n553), .B1(new_n554), .B2(G1698), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n552), .B1(new_n555), .B2(new_n265), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n550), .B(new_n509), .C1(new_n556), .C2(new_n312), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G169), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n554), .A2(G1698), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(G250), .B2(G1698), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n560), .A2(new_n272), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n326), .B1(new_n561), .B2(new_n552), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n562), .A2(G179), .A3(new_n509), .A4(new_n550), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT89), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n542), .A2(new_n549), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n558), .A2(new_n563), .A3(KEYINPUT89), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n531), .A2(new_n538), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(KEYINPUT24), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n539), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n548), .B1(new_n570), .B2(new_n254), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n557), .A2(new_n388), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n572), .B1(G190), .B2(new_n557), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n566), .A2(new_n567), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n507), .A2(G257), .A3(new_n312), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n509), .ZN(new_n576));
  INV_X1    g0376(.A(new_n487), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n451), .A2(G1698), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n578), .A2(new_n269), .A3(new_n271), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT4), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n577), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n265), .A2(KEYINPUT4), .A3(new_n578), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n269), .A2(new_n271), .A3(G250), .A4(G1698), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(KEYINPUT80), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT80), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n265), .A2(new_n585), .A3(G250), .A4(G1698), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n581), .A2(new_n582), .A3(new_n584), .A4(new_n586), .ZN(new_n587));
  AOI211_X1 g0387(.A(G179), .B(new_n576), .C1(new_n587), .C2(new_n326), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n326), .ZN(new_n589));
  INV_X1    g0389(.A(new_n576), .ZN(new_n590));
  AOI21_X1  g0390(.A(G169), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n345), .A2(new_n287), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(G107), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n536), .A2(G97), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n488), .A2(G107), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g0397(.A(KEYINPUT78), .B(KEYINPUT6), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT6), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n600), .A2(KEYINPUT78), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n600), .A2(KEYINPUT78), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n595), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n599), .A2(new_n603), .A3(G20), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT79), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n277), .A2(G77), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n594), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n605), .B1(new_n604), .B2(new_n606), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n254), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  MUX2_X1   g0410(.A(new_n252), .B(new_n547), .S(G97), .Z(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n592), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n576), .B1(new_n587), .B2(new_n326), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n614), .A2(G200), .ZN(new_n615));
  AOI211_X1 g0415(.A(G190), .B(new_n576), .C1(new_n587), .C2(new_n326), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n610), .B(new_n611), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(G250), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n618), .B1(new_n208), .B2(G45), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n378), .A2(new_n505), .B1(new_n312), .B2(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(G238), .A2(G1698), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n621), .B1(new_n451), .B2(G1698), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n479), .A2(new_n481), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n622), .A2(new_n265), .B1(new_n623), .B2(G33), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n620), .B1(new_n624), .B2(new_n312), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT83), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n625), .A2(new_n626), .A3(G179), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n480), .A2(G116), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n477), .A2(KEYINPUT82), .ZN(new_n629));
  OAI21_X1  g0429(.A(G33), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n381), .A2(new_n367), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n451), .A2(G1698), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n269), .A2(new_n631), .A3(new_n271), .A4(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n312), .B1(new_n630), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n312), .A2(G274), .A3(new_n505), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n312), .A2(new_n619), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(KEYINPUT83), .B1(new_n638), .B2(new_n466), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n627), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n456), .B(KEYINPUT84), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n641), .A2(new_n252), .A3(new_n421), .A4(new_n546), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT19), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n209), .B1(new_n371), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n324), .A2(new_n488), .A3(new_n536), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n269), .A2(new_n271), .A3(new_n209), .A4(G68), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n643), .B1(new_n359), .B2(new_n488), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n649), .A2(new_n254), .B1(new_n353), .B2(new_n456), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n642), .A2(new_n650), .B1(new_n625), .B2(new_n329), .ZN(new_n651));
  OAI21_X1  g0451(.A(G200), .B1(new_n634), .B2(new_n637), .ZN(new_n652));
  OAI211_X1 g0452(.A(G190), .B(new_n620), .C1(new_n624), .C2(new_n312), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n421), .A2(G87), .A3(new_n252), .A4(new_n546), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n653), .A2(new_n654), .A3(new_n650), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n640), .A2(new_n651), .B1(new_n652), .B2(new_n655), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n574), .A2(new_n613), .A3(new_n617), .A4(new_n656), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n476), .A2(new_n525), .A3(new_n657), .ZN(G372));
  INV_X1    g0458(.A(new_n447), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n332), .A2(new_n350), .ZN(new_n660));
  INV_X1    g0460(.A(new_n390), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n467), .A2(new_n463), .A3(new_n453), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n661), .A2(new_n662), .B1(new_n399), .B2(new_n400), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n342), .A2(new_n343), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n660), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n659), .B1(new_n665), .B2(new_n441), .ZN(new_n666));
  INV_X1    g0466(.A(new_n639), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n638), .A2(KEYINPUT83), .A3(new_n466), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(new_n651), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n655), .A2(new_n652), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT26), .B1(new_n613), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n638), .A2(new_n466), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n651), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT90), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n675), .B1(new_n625), .B2(G200), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n675), .B(G200), .C1(new_n634), .C2(new_n637), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n679), .A2(new_n655), .B1(new_n651), .B2(new_n673), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT26), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n680), .A2(new_n681), .A3(new_n612), .A4(new_n592), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n672), .A2(new_n674), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n571), .A2(new_n573), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n613), .A2(new_n684), .A3(new_n617), .A4(new_n680), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n521), .A2(new_n522), .A3(new_n524), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n542), .A2(new_n549), .B1(new_n558), .B2(new_n563), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n683), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n666), .B1(new_n476), .B2(new_n690), .ZN(G369));
  NAND2_X1  g0491(.A1(new_n485), .A2(new_n209), .ZN(new_n692));
  OR2_X1    g0492(.A1(new_n692), .A2(KEYINPUT27), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(KEYINPUT27), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(G213), .A3(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(G343), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n496), .A2(new_n698), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n525), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n686), .A2(new_n699), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT91), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G330), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n574), .B1(new_n571), .B2(new_n698), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n542), .A2(new_n549), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n564), .A2(new_n565), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(new_n708), .A3(new_n567), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n706), .B1(new_n709), .B2(new_n698), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n705), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n686), .A2(new_n698), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n709), .A2(new_n684), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n714), .B1(new_n687), .B2(new_n698), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n711), .A2(new_n715), .ZN(G399));
  INV_X1    g0516(.A(KEYINPUT29), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n717), .B(new_n698), .C1(new_n683), .C2(new_n689), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n684), .A2(new_n680), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n709), .A2(new_n521), .A3(new_n522), .A4(new_n524), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT94), .ZN(new_n721));
  AND3_X1   g0521(.A1(new_n613), .A2(new_n721), .A3(new_n617), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n721), .B1(new_n613), .B2(new_n617), .ZN(new_n723));
  OAI211_X1 g0523(.A(new_n719), .B(new_n720), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n679), .A2(new_n655), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n674), .ZN(new_n726));
  OAI21_X1  g0526(.A(KEYINPUT26), .B1(new_n613), .B2(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n656), .A2(new_n681), .A3(new_n612), .A4(new_n592), .ZN(new_n728));
  AND3_X1   g0528(.A1(new_n727), .A2(new_n674), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n697), .B1(new_n724), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n718), .B1(new_n730), .B2(new_n717), .ZN(new_n731));
  AND3_X1   g0531(.A1(new_n613), .A2(new_n617), .A3(new_n656), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n525), .A2(new_n697), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n732), .A2(new_n733), .A3(new_n574), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT31), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n638), .A2(G179), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n523), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n589), .A2(new_n590), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(new_n557), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT92), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n737), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n738), .A2(KEYINPUT92), .A3(new_n557), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n550), .B1(new_n556), .B2(new_n312), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n625), .A2(new_n743), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n614), .A2(new_n744), .ZN(new_n745));
  OAI211_X1 g0545(.A(G179), .B(new_n501), .C1(new_n511), .C2(new_n512), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT30), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n745), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n614), .A2(new_n744), .ZN(new_n750));
  OAI21_X1  g0550(.A(KEYINPUT30), .B1(new_n750), .B2(new_n746), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n741), .A2(new_n742), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n735), .B1(new_n752), .B2(new_n698), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n697), .A2(KEYINPUT31), .ZN(new_n754));
  OAI21_X1  g0554(.A(KEYINPUT93), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n557), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n740), .B1(new_n614), .B2(new_n756), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n742), .A2(new_n757), .A3(new_n523), .A4(new_n736), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n748), .B1(new_n745), .B2(new_n747), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n750), .A2(new_n746), .A3(KEYINPUT30), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT93), .ZN(new_n762));
  INV_X1    g0562(.A(new_n754), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n734), .A2(new_n753), .A3(new_n755), .A4(new_n764), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n765), .A2(G330), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n731), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(new_n208), .ZN(new_n768));
  INV_X1    g0568(.A(new_n212), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G41), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n645), .A2(G116), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n771), .A2(G1), .A3(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n217), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n773), .B1(new_n774), .B2(new_n771), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT28), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n768), .A2(new_n776), .ZN(G364));
  NOR2_X1   g0577(.A1(new_n484), .A2(G20), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n208), .B1(new_n778), .B2(G45), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n770), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n705), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n782), .B1(G330), .B2(new_n703), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n781), .B(KEYINPUT95), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n769), .A2(new_n272), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G355), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(G116), .B2(new_n212), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n241), .A2(new_n314), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n265), .B(new_n769), .C1(new_n314), .C2(new_n217), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G13), .A2(G33), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(G20), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n218), .B1(G20), .B2(new_n329), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n795), .B(KEYINPUT96), .Z(new_n796));
  OAI21_X1  g0596(.A(new_n784), .B1(new_n790), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n794), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n209), .A2(G190), .ZN(new_n799));
  NOR2_X1   g0599(.A1(G179), .A2(G200), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n291), .ZN(new_n802));
  XNOR2_X1  g0602(.A(KEYINPUT97), .B(KEYINPUT32), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n209), .A2(new_n466), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n804), .A2(G190), .A3(G200), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n802), .A2(new_n803), .B1(new_n216), .B2(new_n805), .ZN(new_n806));
  NOR4_X1   g0606(.A1(new_n209), .A2(new_n466), .A3(new_n388), .A4(G190), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n806), .B1(G68), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n209), .A2(new_n337), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n466), .A2(G200), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n265), .B1(new_n811), .B2(new_n202), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n799), .A2(new_n810), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n812), .B1(G77), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n209), .B1(new_n800), .B2(G190), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n802), .A2(new_n803), .B1(new_n817), .B2(G97), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT98), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n388), .B2(G179), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n466), .A2(KEYINPUT98), .A3(G200), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n820), .A2(new_n809), .A3(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n820), .A2(new_n799), .A3(new_n821), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  AOI22_X1  g0625(.A1(G87), .A2(new_n823), .B1(new_n825), .B2(G107), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n808), .A2(new_n815), .A3(new_n818), .A4(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(G322), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n811), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(G311), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n272), .B1(new_n813), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n801), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n829), .B(new_n831), .C1(G329), .C2(new_n832), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n805), .B(KEYINPUT99), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(G326), .ZN(new_n835));
  XNOR2_X1  g0635(.A(KEYINPUT33), .B(G317), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n807), .A2(new_n836), .B1(new_n817), .B2(G294), .ZN(new_n837));
  AOI22_X1  g0637(.A1(G303), .A2(new_n823), .B1(new_n825), .B2(G283), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n833), .A2(new_n835), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n798), .B1(new_n827), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n797), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n793), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n841), .B1(new_n702), .B2(new_n842), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n783), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(G396));
  NAND3_X1  g0645(.A1(new_n464), .A2(new_n467), .A3(new_n698), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n469), .A2(new_n470), .B1(new_n463), .B2(new_n697), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n846), .B1(new_n847), .B2(new_n662), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n690), .B2(new_n697), .ZN(new_n849));
  INV_X1    g0649(.A(new_n848), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n698), .B(new_n850), .C1(new_n683), .C2(new_n689), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  OR2_X1    g0652(.A1(new_n852), .A2(new_n766), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n766), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n853), .B(new_n854), .C1(new_n770), .C2(new_n780), .ZN(new_n855));
  INV_X1    g0655(.A(new_n784), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n794), .A2(new_n791), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n856), .B1(new_n358), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n805), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n859), .A2(G303), .B1(new_n814), .B2(new_n623), .ZN(new_n860));
  INV_X1    g0660(.A(G283), .ZN(new_n861));
  INV_X1    g0661(.A(new_n807), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(KEYINPUT100), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n272), .B1(new_n822), .B2(new_n536), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n865), .B(KEYINPUT101), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n817), .A2(G97), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n825), .A2(G87), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n832), .A2(G311), .ZN(new_n869));
  INV_X1    g0669(.A(new_n811), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(G294), .ZN(new_n871));
  AND4_X1   g0671(.A1(new_n867), .A2(new_n868), .A3(new_n869), .A4(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n864), .A2(new_n866), .A3(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT102), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n873), .A2(new_n874), .ZN(new_n876));
  AOI22_X1  g0676(.A1(G143), .A2(new_n870), .B1(new_n814), .B2(G159), .ZN(new_n877));
  INV_X1    g0677(.A(G137), .ZN(new_n878));
  OAI221_X1 g0678(.A(new_n877), .B1(new_n878), .B2(new_n805), .C1(new_n425), .C2(new_n862), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT34), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n825), .A2(G68), .ZN(new_n882));
  INV_X1    g0682(.A(G132), .ZN(new_n883));
  OAI221_X1 g0683(.A(new_n265), .B1(new_n816), .B2(new_n202), .C1(new_n883), .C2(new_n801), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(G50), .B2(new_n823), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n881), .A2(new_n882), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n879), .A2(new_n880), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR3_X1   g0688(.A1(new_n875), .A2(new_n876), .A3(new_n888), .ZN(new_n889));
  OAI221_X1 g0689(.A(new_n858), .B1(new_n850), .B2(new_n792), .C1(new_n798), .C2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n855), .A2(new_n890), .ZN(G384));
  NAND2_X1  g0691(.A1(new_n599), .A2(new_n603), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT35), .ZN(new_n893));
  OAI211_X1 g0693(.A(G116), .B(new_n219), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n894), .B1(new_n893), .B2(new_n892), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n895), .B(KEYINPUT36), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n217), .A2(G77), .A3(new_n281), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n216), .A2(G68), .ZN(new_n898));
  AOI211_X1 g0698(.A(new_n208), .B(G13), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n695), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n307), .B1(new_n289), .B2(new_n295), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n356), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n903), .B1(new_n286), .B2(new_n297), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n901), .B1(new_n904), .B2(new_n264), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n351), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n330), .B1(new_n904), .B2(new_n264), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n908), .A2(new_n905), .A3(new_n340), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT37), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n330), .B1(new_n349), .B2(new_n264), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n901), .B1(new_n349), .B2(new_n264), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT37), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n911), .A2(new_n912), .A3(new_n913), .A4(new_n340), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n907), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT38), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n907), .A2(new_n915), .A3(KEYINPUT38), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n613), .A2(new_n656), .A3(new_n617), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n921), .A2(new_n713), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n761), .A2(new_n697), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n922), .A2(new_n733), .B1(new_n923), .B2(new_n735), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n749), .A2(new_n751), .ZN(new_n925));
  AOI211_X1 g0725(.A(KEYINPUT104), .B(new_n754), .C1(new_n925), .C2(new_n758), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT104), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n761), .B2(new_n763), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n924), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n399), .A2(new_n400), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n400), .A2(new_n697), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n931), .A2(new_n661), .A3(new_n932), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n400), .B(new_n697), .C1(new_n399), .C2(new_n390), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n848), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n930), .A2(KEYINPUT105), .A3(new_n935), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n525), .A2(new_n697), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n698), .B1(new_n925), .B2(new_n758), .ZN(new_n938));
  OAI22_X1  g0738(.A1(new_n657), .A2(new_n937), .B1(KEYINPUT31), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(KEYINPUT104), .B1(new_n752), .B2(new_n754), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n761), .A2(new_n927), .A3(new_n763), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n935), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT105), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n920), .A2(new_n936), .A3(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT40), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AND3_X1   g0748(.A1(new_n907), .A2(new_n915), .A3(KEYINPUT38), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n911), .A2(new_n912), .A3(new_n340), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(KEYINPUT37), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n914), .ZN(new_n952));
  INV_X1    g0752(.A(new_n912), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n351), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(KEYINPUT38), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(KEYINPUT40), .B1(new_n949), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n948), .B1(new_n943), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n475), .A2(new_n930), .ZN(new_n958));
  OAI21_X1  g0758(.A(G330), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(new_n957), .B2(new_n958), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n851), .A2(new_n846), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n933), .A2(new_n934), .ZN(new_n962));
  AOI21_X1  g0762(.A(KEYINPUT38), .B1(new_n907), .B2(new_n915), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n961), .B(new_n962), .C1(new_n949), .C2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT103), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n660), .A2(new_n901), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT39), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n949), .B2(new_n955), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n918), .A2(KEYINPUT39), .A3(new_n919), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n931), .A2(new_n697), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n967), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n965), .B1(new_n964), .B2(new_n966), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n731), .A2(new_n475), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n666), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n975), .B(new_n977), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n960), .A2(new_n978), .B1(new_n208), .B2(new_n778), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n960), .A2(new_n978), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n900), .B1(new_n979), .B2(new_n980), .ZN(G367));
  NAND2_X1  g0781(.A1(new_n612), .A2(new_n697), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n722), .B2(new_n723), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n613), .B1(new_n983), .B2(new_n709), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n698), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n592), .A2(new_n612), .A3(new_n697), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n983), .A2(new_n986), .ZN(new_n987));
  AND3_X1   g0787(.A1(new_n987), .A2(KEYINPUT42), .A3(new_n714), .ZN(new_n988));
  AOI21_X1  g0788(.A(KEYINPUT42), .B1(new_n987), .B2(new_n714), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n985), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n698), .B1(new_n650), .B2(new_n654), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n991), .A2(new_n651), .A3(new_n673), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n726), .B2(new_n991), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT43), .Z(new_n994));
  NAND2_X1  g0794(.A1(new_n990), .A2(new_n994), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT107), .Z(new_n996));
  NOR2_X1   g0796(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n985), .B(new_n997), .C1(new_n988), .C2(new_n989), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT106), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n996), .A2(new_n999), .A3(KEYINPUT108), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(KEYINPUT108), .B1(new_n996), .B2(new_n999), .ZN(new_n1002));
  AND2_X1   g0802(.A1(new_n983), .A2(new_n986), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n1001), .A2(new_n1002), .B1(new_n711), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1002), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n711), .A2(new_n1003), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1005), .A2(new_n1006), .A3(new_n1000), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n987), .A2(new_n715), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1008), .B(KEYINPUT45), .Z(new_n1009));
  NOR2_X1   g0809(.A1(new_n987), .A2(new_n715), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT44), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(new_n711), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n704), .A2(KEYINPUT109), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n714), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n712), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1015), .B1(new_n710), .B2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1014), .B(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n767), .B1(new_n1013), .B2(new_n1018), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n770), .B(KEYINPUT41), .Z(new_n1020));
  OAI21_X1  g0820(.A(new_n779), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1004), .A2(new_n1007), .A3(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n769), .A2(new_n265), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n237), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n212), .A2(new_n456), .ZN(new_n1025));
  NOR3_X1   g0825(.A1(new_n1025), .A2(new_n793), .A3(new_n794), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n856), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G303), .A2(new_n870), .B1(new_n814), .B2(G283), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n536), .B2(new_n816), .C1(new_n551), .C2(new_n862), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(G311), .B2(new_n834), .ZN(new_n1030));
  INV_X1    g0830(.A(G317), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n272), .B1(new_n801), .B2(new_n1031), .C1(new_n824), .C2(new_n488), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1033), .A2(KEYINPUT110), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(KEYINPUT110), .ZN(new_n1035));
  OAI21_X1  g0835(.A(KEYINPUT46), .B1(new_n822), .B2(new_n477), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n623), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1037), .A2(KEYINPUT46), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1036), .B1(new_n1038), .B2(new_n822), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1030), .A2(new_n1034), .A3(new_n1035), .A4(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n834), .A2(G143), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n817), .A2(G68), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1041), .B(new_n1042), .C1(new_n425), .C2(new_n811), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT111), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n265), .B1(new_n801), .B2(new_n878), .C1(new_n822), .C2(new_n202), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(G77), .B2(new_n825), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n862), .A2(new_n291), .B1(new_n216), .B2(new_n813), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT112), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1045), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1040), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT47), .Z(new_n1053));
  OAI221_X1 g0853(.A(new_n1027), .B1(new_n842), .B2(new_n993), .C1(new_n1053), .C2(new_n798), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1022), .A2(new_n1054), .ZN(G387));
  AOI21_X1  g0855(.A(new_n265), .B1(new_n832), .B2(G326), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n1037), .B2(new_n824), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n822), .A2(new_n551), .B1(new_n861), .B2(new_n816), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(G317), .A2(new_n870), .B1(new_n814), .B2(G303), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n830), .B2(new_n862), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(G322), .B2(new_n834), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1058), .B1(new_n1061), .B2(KEYINPUT48), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT115), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(KEYINPUT48), .B2(new_n1061), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n1064), .A2(KEYINPUT49), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(KEYINPUT49), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1057), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n641), .A2(new_n817), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n823), .A2(G77), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1068), .B(new_n1069), .C1(new_n488), .C2(new_n824), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n265), .B1(new_n813), .B2(new_n203), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n811), .A2(new_n216), .B1(new_n801), .B2(new_n425), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n862), .A2(new_n424), .B1(new_n291), .B2(new_n805), .ZN(new_n1073));
  NOR4_X1   g0873(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .A4(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n794), .B1(new_n1067), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n772), .ZN(new_n1076));
  AOI211_X1 g0876(.A(G45), .B(new_n1076), .C1(G68), .C2(G77), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT113), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  OR3_X1    g0879(.A1(new_n424), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1080));
  OAI21_X1  g0880(.A(KEYINPUT50), .B1(new_n424), .B2(G50), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n1023), .B1(new_n314), .B2(new_n234), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n785), .A2(new_n1076), .B1(new_n536), .B2(new_n769), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1086), .A2(KEYINPUT114), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1087), .A2(new_n796), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1086), .A2(KEYINPUT114), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n856), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1075), .B(new_n1090), .C1(new_n710), .C2(new_n842), .ZN(new_n1091));
  OR2_X1    g0891(.A1(new_n1091), .A2(KEYINPUT116), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(KEYINPUT116), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1092), .A2(new_n1093), .B1(new_n780), .B2(new_n1018), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1018), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n1095), .A2(new_n767), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n770), .B1(new_n1095), .B2(new_n767), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1094), .B1(new_n1096), .B2(new_n1097), .ZN(G393));
  NOR2_X1   g0898(.A1(new_n1095), .A2(new_n767), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n771), .B1(new_n1099), .B2(new_n1013), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n1013), .B2(new_n1099), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1023), .A2(new_n244), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1102), .B(new_n795), .C1(new_n488), .C2(new_n212), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n868), .B1(new_n203), .B2(new_n822), .ZN(new_n1104));
  INV_X1    g0904(.A(G143), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n265), .B1(new_n801), .B2(new_n1105), .C1(new_n424), .C2(new_n813), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n862), .A2(new_n216), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n816), .A2(new_n358), .ZN(new_n1108));
  NOR4_X1   g0908(.A1(new_n1104), .A2(new_n1106), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n805), .A2(new_n425), .B1(new_n811), .B2(new_n291), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT51), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n805), .A2(new_n1031), .B1(new_n811), .B2(new_n830), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT52), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n862), .A2(new_n499), .B1(new_n816), .B2(new_n1037), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n272), .B1(new_n801), .B2(new_n828), .C1(new_n551), .C2(new_n813), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n822), .A2(new_n861), .B1(new_n824), .B2(new_n536), .ZN(new_n1116));
  NOR3_X1   g0916(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1109), .A2(new_n1111), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n784), .B(new_n1103), .C1(new_n1118), .C2(new_n798), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(new_n1003), .B2(new_n793), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(new_n1013), .B2(new_n780), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1101), .A2(new_n1121), .ZN(G390));
  NAND2_X1  g0922(.A1(new_n969), .A2(new_n970), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n971), .B1(new_n961), .B2(new_n962), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n765), .A2(G330), .A3(new_n850), .A4(new_n962), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n962), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n724), .A2(new_n729), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n847), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n468), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1129), .A2(new_n698), .A3(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1128), .B1(new_n1132), .B2(new_n846), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n949), .A2(new_n955), .B1(new_n931), .B2(new_n697), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1126), .B(new_n1127), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(G330), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(new_n924), .B2(new_n929), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1124), .B1(new_n969), .B2(new_n970), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n935), .B(new_n1137), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1135), .A2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1141), .A2(new_n779), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1123), .A2(new_n791), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n857), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n784), .B1(new_n249), .B2(new_n1144), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n813), .A2(new_n488), .B1(new_n801), .B2(new_n551), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n265), .B(new_n1146), .C1(G116), .C2(new_n870), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n805), .A2(new_n861), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n1108), .B(new_n1148), .C1(G107), .C2(new_n807), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n823), .A2(G87), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1147), .A2(new_n1149), .A3(new_n1150), .A4(new_n882), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n862), .A2(new_n878), .B1(new_n816), .B2(new_n291), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(G128), .B2(new_n859), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n825), .A2(G50), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(KEYINPUT54), .B(G143), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n272), .B1(new_n814), .B2(new_n1156), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(G132), .A2(new_n870), .B1(new_n832), .B2(G125), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1153), .A2(new_n1154), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n823), .A2(G150), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT53), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1151), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1145), .B1(new_n1162), .B2(new_n794), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1142), .B1(new_n1143), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n475), .A2(new_n1137), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n976), .A2(new_n666), .A3(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n765), .A2(G330), .A3(new_n850), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1128), .A2(new_n1167), .B1(new_n1137), .B2(new_n935), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n961), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1127), .A2(new_n1132), .A3(new_n846), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n962), .B1(new_n1137), .B2(new_n850), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n1168), .A2(new_n1169), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT117), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n1166), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1173), .B1(new_n1166), .B2(new_n1172), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n1141), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1135), .B(new_n1140), .C1(new_n1174), .C2(new_n1175), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1177), .A2(new_n770), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1164), .A2(new_n1179), .ZN(G378));
  OAI21_X1  g0980(.A(KEYINPUT122), .B1(new_n973), .B2(new_n974), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n974), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT122), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1182), .A2(new_n1183), .A3(new_n972), .A4(new_n967), .ZN(new_n1184));
  AND2_X1   g0984(.A1(new_n1181), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n952), .A2(new_n954), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(new_n917), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n947), .B1(new_n1187), .B2(new_n919), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n943), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1136), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n441), .A2(new_n447), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n430), .A2(new_n901), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1191), .B(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1194));
  XOR2_X1   g0994(.A(new_n1193), .B(new_n1194), .Z(new_n1195));
  INV_X1    g0995(.A(KEYINPUT120), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n948), .A2(new_n1190), .A3(new_n1195), .A4(new_n1196), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n918), .A2(new_n919), .B1(new_n943), .B2(new_n944), .ZN(new_n1198));
  AOI21_X1  g0998(.A(KEYINPUT40), .B1(new_n1198), .B2(new_n936), .ZN(new_n1199));
  OAI21_X1  g0999(.A(G330), .B1(new_n956), .B2(new_n943), .ZN(new_n1200));
  OAI21_X1  g1000(.A(KEYINPUT120), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n948), .A2(new_n1190), .A3(new_n1196), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1195), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1185), .A2(KEYINPUT121), .A3(new_n1197), .A4(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1204), .A2(KEYINPUT121), .A3(new_n1197), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1181), .A2(new_n1184), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1178), .A2(new_n1166), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1205), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT57), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(KEYINPUT123), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT123), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1210), .A2(new_n1214), .A3(new_n1211), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1204), .A2(new_n1197), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n975), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1204), .A2(new_n975), .A3(new_n1197), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1211), .B1(new_n1178), .B2(new_n1166), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n771), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1213), .A2(new_n1215), .A3(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1205), .A2(new_n1208), .A3(new_n780), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n781), .B1(G50), .B2(new_n1144), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n825), .A2(G58), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n641), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1227), .B1(new_n1228), .B2(new_n813), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1042), .B1(new_n477), .B2(new_n805), .C1(new_n862), .C2(new_n488), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n832), .A2(G283), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n265), .A2(G41), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n870), .A2(G107), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1069), .A2(new_n1231), .A3(new_n1232), .A4(new_n1233), .ZN(new_n1234));
  NOR3_X1   g1034(.A1(new_n1229), .A2(new_n1230), .A3(new_n1234), .ZN(new_n1235));
  XOR2_X1   g1035(.A(new_n1235), .B(KEYINPUT58), .Z(new_n1236));
  INV_X1    g1036(.A(G128), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n811), .A2(new_n1237), .B1(new_n813), .B2(new_n878), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(G125), .B2(new_n859), .ZN(new_n1239));
  OR3_X1    g1039(.A1(new_n822), .A2(KEYINPUT118), .A3(new_n1155), .ZN(new_n1240));
  OAI21_X1  g1040(.A(KEYINPUT118), .B1(new_n822), .B2(new_n1155), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(G132), .A2(new_n807), .B1(new_n817), .B2(G150), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1239), .A2(new_n1240), .A3(new_n1241), .A4(new_n1242), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1243), .A2(KEYINPUT59), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(KEYINPUT59), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n825), .A2(G159), .ZN(new_n1246));
  AOI211_X1 g1046(.A(G33), .B(G41), .C1(new_n832), .C2(G124), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n1236), .B1(new_n1244), .B2(new_n1248), .C1(new_n1232), .C2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT119), .ZN(new_n1251));
  OR2_X1    g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n798), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1226), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1254), .B1(new_n1203), .B2(new_n792), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1225), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1224), .A2(new_n1257), .ZN(G375));
  OR2_X1    g1058(.A1(new_n1166), .A2(new_n1172), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1176), .A2(new_n1259), .ZN(new_n1260));
  OR2_X1    g1060(.A1(new_n1260), .A2(new_n1020), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1128), .A2(new_n791), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n784), .B1(G68), .B2(new_n1144), .ZN(new_n1263));
  OAI221_X1 g1063(.A(new_n1068), .B1(new_n358), .B2(new_n824), .C1(new_n488), .C2(new_n822), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n859), .A2(G294), .B1(new_n807), .B2(new_n623), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(G107), .A2(new_n814), .B1(new_n832), .B2(G303), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n265), .B1(new_n870), .B2(G283), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1265), .A2(new_n1266), .A3(new_n1267), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n859), .A2(G132), .B1(new_n807), .B2(new_n1156), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n216), .B2(new_n816), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(G150), .A2(new_n814), .B1(new_n832), .B2(G128), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n272), .B1(new_n870), .B2(G137), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n823), .A2(G159), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1271), .A2(new_n1272), .A3(new_n1227), .A4(new_n1273), .ZN(new_n1274));
  OAI22_X1  g1074(.A1(new_n1264), .A2(new_n1268), .B1(new_n1270), .B2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1263), .B1(new_n1275), .B2(new_n794), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(new_n1172), .A2(new_n780), .B1(new_n1262), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1261), .A2(new_n1277), .ZN(G381));
  INV_X1    g1078(.A(KEYINPUT124), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(G378), .A2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1164), .A2(new_n1179), .A3(KEYINPUT124), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(G375), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(G387), .ZN(new_n1284));
  INV_X1    g1084(.A(G381), .ZN(new_n1285));
  NOR4_X1   g1085(.A1(G390), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1283), .A2(new_n1284), .A3(new_n1285), .A4(new_n1286), .ZN(G407));
  NAND2_X1  g1087(.A1(new_n696), .A2(G213), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1283), .A2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(G407), .A2(G213), .A3(new_n1290), .ZN(G409));
  XNOR2_X1  g1091(.A(G393), .B(new_n844), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1022), .A2(new_n1054), .A3(G390), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(G390), .B1(new_n1022), .B2(new_n1054), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1293), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1296), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1298), .A2(new_n1292), .A3(new_n1294), .ZN(new_n1299));
  AND2_X1   g1099(.A1(new_n1297), .A2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1277), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1260), .A2(KEYINPUT60), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT60), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n771), .B1(new_n1259), .B2(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1302), .B1(new_n1303), .B2(new_n1305), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(new_n1306), .B(G384), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1289), .A2(G2897), .ZN(new_n1308));
  XOR2_X1   g1108(.A(new_n1308), .B(KEYINPUT126), .Z(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  XNOR2_X1  g1110(.A(new_n1307), .B(new_n1310), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1210), .A2(new_n1020), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1255), .B1(new_n1220), .B2(new_n779), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1314), .A2(new_n1282), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1214), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1222), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n770), .B1(new_n1317), .B2(new_n1220), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1316), .A2(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1256), .B1(new_n1319), .B2(new_n1215), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1315), .B1(new_n1320), .B2(G378), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1311), .B1(new_n1321), .B2(new_n1289), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT61), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1224), .A2(G378), .A3(new_n1257), .ZN(new_n1324));
  OR2_X1    g1124(.A1(new_n1314), .A2(new_n1282), .ZN(new_n1325));
  AOI211_X1 g1125(.A(new_n1289), .B(new_n1307), .C1(new_n1324), .C2(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(KEYINPUT125), .B1(KEYINPUT127), .B2(KEYINPUT62), .ZN(new_n1327));
  OAI211_X1 g1127(.A(new_n1322), .B(new_n1323), .C1(new_n1326), .C2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT125), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1307), .ZN(new_n1331));
  NAND4_X1  g1131(.A1(new_n1329), .A2(new_n1330), .A3(new_n1288), .A4(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(KEYINPUT62), .B1(new_n1332), .B2(KEYINPUT127), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1301), .B1(new_n1328), .B2(new_n1333), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1289), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1335));
  XNOR2_X1  g1135(.A(new_n1307), .B(new_n1309), .ZN(new_n1336));
  OAI211_X1 g1136(.A(new_n1300), .B(new_n1323), .C1(new_n1335), .C2(new_n1336), .ZN(new_n1337));
  AND4_X1   g1137(.A1(KEYINPUT63), .A2(new_n1329), .A3(new_n1288), .A4(new_n1331), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1329), .A2(new_n1288), .A3(new_n1331), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1340), .A2(KEYINPUT125), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT63), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1341), .A2(new_n1342), .A3(new_n1332), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1339), .A2(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1334), .A2(new_n1344), .ZN(G405));
  NAND3_X1  g1145(.A1(G375), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1346), .A2(new_n1324), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1347), .A2(new_n1331), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1346), .A2(new_n1324), .A3(new_n1307), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1350));
  XNOR2_X1  g1150(.A(new_n1350), .B(new_n1301), .ZN(G402));
endmodule


