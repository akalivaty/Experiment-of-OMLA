//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 1 0 0 1 0 0 0 0 0 1 1 1 0 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1325,
    new_n1326, new_n1328, new_n1329, new_n1330, new_n1331, new_n1332,
    new_n1333, new_n1335, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1402, new_n1403, new_n1404, new_n1405, new_n1406, new_n1407,
    new_n1408, new_n1409;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(KEYINPUT64), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT64), .ZN(new_n212));
  NAND3_X1  g0012(.A1(new_n212), .A2(G1), .A3(G13), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(new_n201), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G50), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n209), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n222));
  INV_X1    g0022(.A(G77), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  INV_X1    g0024(.A(G107), .ZN(new_n225));
  INV_X1    g0025(.A(G264), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n206), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(KEYINPUT1), .ZN(new_n232));
  OR2_X1    g0032(.A1(new_n231), .A2(KEYINPUT1), .ZN(new_n233));
  NAND3_X1  g0033(.A1(new_n221), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(KEYINPUT65), .Z(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n244), .B(new_n245), .Z(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  OAI21_X1  g0051(.A(KEYINPUT79), .B1(new_n251), .B2(KEYINPUT3), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT79), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT3), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n253), .A2(new_n254), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n252), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G223), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n260), .B1(G226), .B2(new_n259), .ZN(new_n261));
  INV_X1    g0061(.A(G87), .ZN(new_n262));
  OAI22_X1  g0062(.A1(new_n257), .A2(new_n261), .B1(new_n251), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G41), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n214), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G274), .ZN(new_n268));
  INV_X1    g0068(.A(new_n210), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n268), .B1(new_n269), .B2(new_n264), .ZN(new_n270));
  OR2_X1    g0070(.A1(KEYINPUT66), .A2(G41), .ZN(new_n271));
  INV_X1    g0071(.A(G45), .ZN(new_n272));
  NAND2_X1  g0072(.A1(KEYINPUT66), .A2(G41), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G1), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n270), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G232), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n264), .A2(G1), .A3(G13), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n275), .B1(G41), .B2(G45), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n276), .B1(new_n277), .B2(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n267), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G169), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G179), .ZN(new_n285));
  NOR3_X1   g0085(.A1(new_n267), .A2(new_n285), .A3(new_n281), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT80), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT7), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n257), .A2(new_n289), .A3(new_n216), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G68), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n289), .B1(new_n257), .B2(new_n216), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n288), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  AND3_X1   g0093(.A1(new_n252), .A2(new_n255), .A3(new_n256), .ZN(new_n294));
  OAI21_X1  g0094(.A(KEYINPUT7), .B1(new_n294), .B2(G20), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n295), .A2(KEYINPUT80), .A3(G68), .A4(new_n290), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G58), .ZN(new_n298));
  INV_X1    g0098(.A(G68), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OR2_X1    g0100(.A1(new_n300), .A2(new_n201), .ZN(new_n301));
  NOR2_X1   g0101(.A1(G20), .A2(G33), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n301), .A2(G20), .B1(G159), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n297), .A2(KEYINPUT16), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT16), .ZN(new_n305));
  INV_X1    g0105(.A(new_n303), .ZN(new_n306));
  XNOR2_X1  g0106(.A(KEYINPUT3), .B(G33), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n289), .B1(new_n307), .B2(G20), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n254), .A2(G33), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n256), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n310), .A2(KEYINPUT7), .A3(new_n216), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n299), .B1(new_n308), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n305), .B1(new_n306), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n211), .A2(new_n213), .A3(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n304), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n298), .A2(KEYINPUT8), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT8), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G58), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n317), .A2(new_n319), .A3(KEYINPUT69), .ZN(new_n320));
  OR3_X1    g0120(.A1(new_n318), .A2(KEYINPUT69), .A3(G58), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n216), .A2(G1), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n275), .A2(G13), .A3(G20), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n211), .A2(new_n213), .A3(new_n325), .A4(new_n314), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n325), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n324), .A2(new_n327), .B1(new_n328), .B2(new_n322), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n287), .B1(new_n316), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT18), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n329), .ZN(new_n333));
  AND3_X1   g0133(.A1(new_n211), .A2(new_n213), .A3(new_n314), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n306), .B1(new_n293), .B2(new_n296), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n334), .B1(new_n335), .B2(KEYINPUT16), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n333), .B1(new_n336), .B2(new_n313), .ZN(new_n337));
  OAI21_X1  g0137(.A(KEYINPUT18), .B1(new_n337), .B2(new_n287), .ZN(new_n338));
  AND2_X1   g0138(.A1(new_n332), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G190), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n282), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(G200), .B2(new_n282), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n316), .A2(new_n329), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT17), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n316), .A2(KEYINPUT17), .A3(new_n329), .A4(new_n342), .ZN(new_n346));
  AND3_X1   g0146(.A1(new_n345), .A2(KEYINPUT81), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(KEYINPUT81), .B1(new_n345), .B2(new_n346), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n339), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT14), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT13), .ZN(new_n351));
  NAND2_X1  g0151(.A1(G33), .A2(G97), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n310), .A2(G1698), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n353), .B1(new_n354), .B2(G226), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n256), .A2(new_n309), .A3(G232), .A4(G1698), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT74), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n307), .A2(KEYINPUT74), .A3(G232), .A4(G1698), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n266), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT75), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n276), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n270), .A2(new_n274), .A3(KEYINPUT75), .A4(new_n275), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n278), .A2(G238), .A3(new_n279), .ZN(new_n366));
  AND3_X1   g0166(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n351), .B1(new_n362), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n265), .B1(new_n355), .B2(new_n360), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n370));
  NOR3_X1   g0170(.A1(new_n369), .A2(new_n370), .A3(KEYINPUT13), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n350), .B(G169), .C1(new_n368), .C2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT78), .ZN(new_n373));
  OAI21_X1  g0173(.A(G169), .B1(new_n368), .B2(new_n371), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT14), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n362), .A2(new_n367), .A3(new_n351), .ZN(new_n376));
  OAI21_X1  g0176(.A(KEYINPUT13), .B1(new_n369), .B2(new_n370), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n283), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT78), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n378), .A2(new_n379), .A3(new_n350), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n376), .A2(G179), .A3(new_n377), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n373), .A2(new_n375), .A3(new_n380), .A4(new_n381), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n302), .A2(G50), .B1(G20), .B2(new_n299), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n251), .A2(G20), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n383), .B1(new_n385), .B2(new_n223), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n315), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n387), .B(KEYINPUT11), .ZN(new_n388));
  OR2_X1    g0188(.A1(new_n388), .A2(KEYINPUT77), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(KEYINPUT77), .ZN(new_n390));
  NOR3_X1   g0190(.A1(new_n326), .A2(new_n299), .A3(new_n323), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT12), .B1(new_n325), .B2(G68), .ZN(new_n392));
  OR3_X1    g0192(.A1(new_n325), .A2(KEYINPUT12), .A3(G68), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n389), .A2(new_n390), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n382), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n320), .A2(new_n321), .A3(new_n384), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n302), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n334), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n323), .A2(new_n202), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  OAI22_X1  g0201(.A1(new_n401), .A2(new_n326), .B1(G50), .B2(new_n325), .ZN(new_n402));
  OR2_X1    g0202(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT68), .B1(new_n310), .B2(new_n259), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT68), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n307), .A2(new_n405), .A3(G1698), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n258), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n307), .A2(new_n259), .ZN(new_n408));
  INV_X1    g0208(.A(G222), .ZN(new_n409));
  OAI22_X1  g0209(.A1(new_n408), .A2(new_n409), .B1(new_n223), .B2(new_n307), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n266), .B1(new_n407), .B2(new_n410), .ZN(new_n411));
  XNOR2_X1  g0211(.A(KEYINPUT67), .B(G226), .ZN(new_n412));
  OR2_X1    g0212(.A1(new_n280), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n276), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n403), .B1(new_n417), .B2(G169), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT70), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n416), .B2(G179), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n417), .A2(KEYINPUT70), .A3(new_n285), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n418), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n402), .ZN(new_n423));
  AND2_X1   g0223(.A1(new_n397), .A2(new_n398), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n423), .B(KEYINPUT9), .C1(new_n424), .C2(new_n334), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT9), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(new_n399), .B2(new_n402), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n411), .A2(G190), .A3(new_n415), .ZN(new_n429));
  INV_X1    g0229(.A(G200), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n430), .B1(new_n411), .B2(new_n415), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n428), .B(new_n429), .C1(new_n431), .C2(KEYINPUT73), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(KEYINPUT73), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(KEYINPUT10), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n428), .A2(new_n429), .ZN(new_n436));
  OR2_X1    g0236(.A1(new_n431), .A2(KEYINPUT73), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT10), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n436), .A2(new_n437), .A3(new_n438), .A4(new_n433), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n422), .B1(new_n435), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n376), .A2(G190), .A3(new_n377), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT76), .ZN(new_n442));
  XNOR2_X1  g0242(.A(new_n441), .B(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n430), .B1(new_n376), .B2(new_n377), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n395), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n278), .A2(G244), .A3(new_n279), .ZN(new_n447));
  OAI22_X1  g0247(.A1(new_n408), .A2(new_n277), .B1(new_n225), .B2(new_n307), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n404), .A2(new_n406), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n448), .B1(new_n449), .B2(G238), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n276), .B(new_n447), .C1(new_n450), .C2(new_n265), .ZN(new_n451));
  OR2_X1    g0251(.A1(new_n451), .A2(G179), .ZN(new_n452));
  NOR3_X1   g0252(.A1(new_n326), .A2(new_n223), .A3(new_n323), .ZN(new_n453));
  XNOR2_X1  g0253(.A(new_n453), .B(KEYINPUT72), .ZN(new_n454));
  XNOR2_X1  g0254(.A(KEYINPUT8), .B(G58), .ZN(new_n455));
  INV_X1    g0255(.A(new_n302), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n457), .B1(G20), .B2(G77), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n262), .A2(KEYINPUT15), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT15), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G87), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT71), .ZN(new_n463));
  XNOR2_X1  g0263(.A(KEYINPUT15), .B(G87), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT71), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n463), .A2(new_n466), .A3(new_n384), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n334), .B1(new_n458), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n325), .A2(G77), .ZN(new_n469));
  NOR3_X1   g0269(.A1(new_n454), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n451), .A2(new_n283), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n452), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n451), .A2(G200), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n474), .B(new_n470), .C1(new_n340), .C2(new_n451), .ZN(new_n475));
  AND2_X1   g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n396), .A2(new_n440), .A3(new_n446), .A4(new_n476), .ZN(new_n477));
  NOR3_X1   g0277(.A1(new_n349), .A2(new_n477), .A3(KEYINPUT82), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT82), .ZN(new_n479));
  AND4_X1   g0279(.A1(new_n396), .A2(new_n440), .A3(new_n446), .A4(new_n476), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n332), .A2(new_n338), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT81), .ZN(new_n482));
  AOI21_X1  g0282(.A(KEYINPUT17), .B1(new_n337), .B2(new_n342), .ZN(new_n483));
  INV_X1    g0283(.A(new_n346), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n345), .A2(KEYINPUT81), .A3(new_n346), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n481), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n479), .B1(new_n480), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n478), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n251), .A2(G1), .ZN(new_n491));
  OAI21_X1  g0291(.A(G116), .B1(new_n326), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(G116), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n325), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(G33), .A2(G283), .ZN(new_n496));
  INV_X1    g0296(.A(G97), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n496), .B(new_n216), .C1(G33), .C2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT20), .ZN(new_n499));
  AOI22_X1  g0299(.A1(KEYINPUT89), .A2(new_n499), .B1(new_n493), .B2(G20), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n315), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT89), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT20), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(KEYINPUT20), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n315), .A2(new_n498), .A3(new_n500), .A4(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n495), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT88), .ZN(new_n508));
  AOI21_X1  g0308(.A(KEYINPUT5), .B1(new_n271), .B2(new_n273), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT5), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n275), .B(G45), .C1(new_n510), .C2(G41), .ZN(new_n511));
  OAI211_X1 g0311(.A(G270), .B(new_n278), .C1(new_n509), .C2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n273), .ZN(new_n513));
  NOR2_X1   g0313(.A1(KEYINPUT66), .A2(G41), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n510), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n511), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n515), .A2(new_n270), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n508), .B1(new_n512), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(G257), .A2(G1698), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n520), .B1(new_n226), .B2(G1698), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n294), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n310), .A2(G303), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n266), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n512), .A2(new_n517), .A3(new_n508), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n519), .A2(new_n525), .A3(G190), .A4(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n526), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n265), .B1(new_n522), .B2(new_n523), .ZN(new_n529));
  NOR3_X1   g0329(.A1(new_n528), .A2(new_n518), .A3(new_n529), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n507), .B(new_n527), .C1(new_n530), .C2(new_n430), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT21), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n506), .A2(G169), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n532), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n530), .A2(G179), .A3(new_n506), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n519), .A2(new_n525), .A3(new_n526), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n536), .A2(KEYINPUT21), .A3(G169), .A4(new_n506), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n531), .A2(new_n534), .A3(new_n535), .A4(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT22), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n216), .A2(G87), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n539), .B1(new_n310), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G116), .ZN(new_n542));
  OR3_X1    g0342(.A1(new_n542), .A2(KEYINPUT90), .A3(G20), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT23), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n216), .B2(G107), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n225), .A2(KEYINPUT23), .A3(G20), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n216), .A2(G33), .A3(G116), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(KEYINPUT90), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n541), .A2(new_n543), .A3(new_n547), .A4(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n252), .A2(new_n255), .A3(new_n216), .A4(new_n256), .ZN(new_n551));
  NAND2_X1  g0351(.A1(KEYINPUT22), .A2(G87), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(KEYINPUT24), .B1(new_n550), .B2(new_n553), .ZN(new_n554));
  OR2_X1    g0354(.A1(new_n551), .A2(new_n552), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT24), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n543), .A2(new_n547), .A3(new_n549), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n555), .A2(new_n556), .A3(new_n541), .A4(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n315), .ZN(new_n560));
  INV_X1    g0360(.A(G250), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n259), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(G257), .B2(new_n259), .ZN(new_n563));
  XNOR2_X1  g0363(.A(KEYINPUT91), .B(G294), .ZN(new_n564));
  OAI22_X1  g0364(.A1(new_n257), .A2(new_n563), .B1(new_n251), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n266), .ZN(new_n566));
  OAI211_X1 g0366(.A(G264), .B(new_n278), .C1(new_n509), .C2(new_n511), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n568), .A2(G190), .A3(new_n517), .ZN(new_n569));
  INV_X1    g0369(.A(new_n491), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n334), .A2(KEYINPUT83), .A3(new_n325), .A4(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT83), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n572), .B1(new_n326), .B2(new_n491), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n571), .A2(new_n573), .A3(G107), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n325), .A2(G107), .ZN(new_n575));
  XNOR2_X1  g0375(.A(new_n575), .B(KEYINPUT25), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n566), .A2(new_n567), .A3(new_n517), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(G200), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n560), .A2(new_n569), .A3(new_n578), .A4(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n283), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n566), .A2(new_n567), .A3(new_n285), .A4(new_n517), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n334), .B1(new_n554), .B2(new_n558), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n582), .B(new_n583), .C1(new_n584), .C2(new_n577), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n538), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n463), .A2(new_n466), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n328), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT19), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n216), .B1(new_n352), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(G97), .A2(G107), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n262), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n216), .A2(G33), .A3(G97), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n591), .A2(new_n593), .B1(new_n590), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n299), .B2(new_n551), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n589), .B1(new_n597), .B2(new_n334), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n571), .A2(new_n573), .A3(G87), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT87), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n571), .A2(new_n573), .A3(KEYINPUT87), .A4(G87), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n598), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT85), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n224), .A2(G1698), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(G238), .B2(G1698), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n542), .B1(new_n257), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n266), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n561), .B1(new_n272), .B2(G1), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n275), .A2(new_n268), .A3(G45), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n278), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n604), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n611), .ZN(new_n613));
  AOI211_X1 g0413(.A(KEYINPUT85), .B(new_n613), .C1(new_n607), .C2(new_n266), .ZN(new_n614));
  OAI21_X1  g0414(.A(G200), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(G238), .A2(G1698), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(new_n224), .B2(G1698), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n617), .A2(new_n256), .A3(new_n252), .A4(new_n255), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n265), .B1(new_n618), .B2(new_n542), .ZN(new_n619));
  OAI21_X1  g0419(.A(KEYINPUT85), .B1(new_n619), .B2(new_n613), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n608), .A2(new_n604), .A3(new_n611), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n620), .A2(G190), .A3(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n603), .A2(new_n615), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n620), .A2(new_n285), .A3(new_n621), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT86), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n588), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n463), .A2(new_n466), .A3(KEYINPUT86), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n626), .A2(new_n573), .A3(new_n571), .A4(new_n627), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n596), .A2(new_n315), .B1(new_n328), .B2(new_n588), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n612), .A2(new_n614), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n624), .B(new_n630), .C1(new_n631), .C2(G169), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n623), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n325), .A2(G97), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n307), .A2(new_n289), .A3(G20), .ZN(new_n635));
  AOI21_X1  g0435(.A(KEYINPUT7), .B1(new_n310), .B2(new_n216), .ZN(new_n636));
  OAI21_X1  g0436(.A(G107), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT6), .ZN(new_n638));
  AND2_X1   g0438(.A1(G97), .A2(G107), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n638), .B1(new_n639), .B2(new_n592), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n225), .A2(KEYINPUT6), .A3(G97), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n642), .A2(G20), .B1(G77), .B2(new_n302), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n637), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n634), .B1(new_n644), .B2(new_n315), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n256), .A2(new_n309), .A3(G250), .A4(G1698), .ZN(new_n646));
  AND2_X1   g0446(.A1(KEYINPUT4), .A2(G244), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n256), .A2(new_n309), .A3(new_n647), .A4(new_n259), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n646), .A2(new_n648), .A3(new_n496), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n224), .A2(G1698), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n252), .A2(new_n255), .A3(new_n256), .A4(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT4), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n265), .B1(new_n649), .B2(new_n653), .ZN(new_n654));
  OAI211_X1 g0454(.A(G257), .B(new_n278), .C1(new_n509), .C2(new_n511), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n517), .ZN(new_n656));
  OAI21_X1  g0456(.A(G200), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n571), .A2(new_n573), .A3(G97), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n651), .A2(new_n652), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n646), .A2(new_n648), .A3(new_n496), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n266), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n655), .A2(new_n517), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(new_n662), .A3(G190), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n645), .A2(new_n657), .A3(new_n658), .A4(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(KEYINPUT84), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n642), .A2(G20), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n302), .A2(G77), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n225), .B1(new_n308), .B2(new_n311), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n315), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n634), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(new_n658), .A3(new_n672), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n654), .A2(new_n285), .A3(new_n656), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n283), .B1(new_n661), .B2(new_n662), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(KEYINPUT84), .B1(new_n676), .B2(new_n664), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n666), .A2(new_n677), .ZN(new_n678));
  AND4_X1   g0478(.A1(new_n490), .A2(new_n587), .A3(new_n633), .A4(new_n678), .ZN(G372));
  INV_X1    g0479(.A(new_n446), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n396), .B1(new_n680), .B2(new_n473), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n485), .A2(new_n486), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n339), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n435), .A2(new_n439), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n422), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n608), .A2(new_n611), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n283), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n624), .A2(new_n630), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT84), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n654), .A2(new_n340), .A3(new_n656), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n430), .B1(new_n661), .B2(new_n662), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n673), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(G169), .B1(new_n654), .B2(new_n656), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n661), .A2(new_n662), .A3(G179), .ZN(new_n695));
  AOI22_X1  g0495(.A1(new_n658), .A2(new_n645), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n690), .B1(new_n693), .B2(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n585), .A2(new_n534), .A3(new_n535), .A4(new_n537), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n697), .A2(new_n698), .A3(new_n581), .A4(new_n665), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n601), .A2(new_n602), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n687), .A2(G200), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n622), .A2(new_n700), .A3(new_n629), .A4(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT92), .ZN(new_n703));
  AND3_X1   g0503(.A1(new_n702), .A2(new_n703), .A3(new_n689), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n703), .B1(new_n702), .B2(new_n689), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n689), .B1(new_n699), .B2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n623), .A2(new_n632), .A3(new_n696), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT26), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n702), .A2(new_n689), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT92), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n702), .A2(new_n703), .A3(new_n689), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(KEYINPUT93), .B1(new_n674), .B2(new_n675), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT93), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n694), .A2(new_n695), .A3(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n715), .A2(new_n673), .A3(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(KEYINPUT26), .B1(new_n714), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n710), .B1(new_n720), .B2(KEYINPUT94), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT94), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n718), .B1(new_n712), .B2(new_n713), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n722), .B1(new_n723), .B2(KEYINPUT26), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n707), .B1(new_n721), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n686), .B1(new_n489), .B2(new_n725), .ZN(G369));
  NAND3_X1  g0526(.A1(new_n275), .A2(new_n216), .A3(G13), .ZN(new_n727));
  OR2_X1    g0527(.A1(new_n727), .A2(KEYINPUT27), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(KEYINPUT27), .ZN(new_n729));
  AND3_X1   g0529(.A1(new_n728), .A2(G213), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(G343), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n506), .A2(new_n732), .ZN(new_n733));
  XOR2_X1   g0533(.A(new_n733), .B(KEYINPUT95), .Z(new_n734));
  NAND3_X1  g0534(.A1(new_n534), .A2(new_n537), .A3(new_n535), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(new_n538), .B2(new_n734), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n737), .A2(G330), .ZN(new_n738));
  INV_X1    g0538(.A(new_n586), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n732), .B1(new_n584), .B2(new_n577), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n741), .B1(new_n585), .B2(new_n731), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n735), .A2(new_n731), .ZN(new_n744));
  INV_X1    g0544(.A(new_n585), .ZN(new_n745));
  AOI22_X1  g0545(.A1(new_n744), .A2(new_n739), .B1(new_n745), .B2(new_n731), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n743), .A2(new_n746), .ZN(G399));
  NOR2_X1   g0547(.A1(new_n513), .A2(new_n514), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n207), .ZN(new_n750));
  OR3_X1    g0550(.A1(new_n749), .A2(KEYINPUT96), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(KEYINPUT96), .B1(new_n749), .B2(new_n750), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n593), .A2(G116), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n753), .A2(G1), .A3(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(new_n219), .B2(new_n753), .ZN(new_n756));
  XNOR2_X1  g0556(.A(new_n756), .B(KEYINPUT28), .ZN(new_n757));
  INV_X1    g0557(.A(G330), .ZN(new_n758));
  AND3_X1   g0558(.A1(new_n568), .A2(new_n661), .A3(new_n662), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n759), .A2(G179), .A3(new_n530), .A4(new_n631), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT30), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n760), .A2(new_n761), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n661), .A2(new_n662), .ZN(new_n765));
  AOI21_X1  g0565(.A(G179), .B1(new_n608), .B2(new_n611), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n536), .A2(new_n579), .A3(new_n765), .A4(new_n766), .ZN(new_n767));
  AND2_X1   g0567(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n763), .B1(new_n768), .B2(KEYINPUT97), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n764), .A2(new_n767), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT97), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OAI211_X1 g0572(.A(KEYINPUT31), .B(new_n732), .C1(new_n769), .C2(new_n772), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n587), .A2(new_n678), .A3(new_n633), .A4(new_n731), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(KEYINPUT31), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n768), .A2(new_n763), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(new_n732), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n758), .B1(new_n773), .B2(new_n778), .ZN(new_n779));
  XOR2_X1   g0579(.A(KEYINPUT98), .B(KEYINPUT29), .Z(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(new_n725), .B2(new_n732), .ZN(new_n782));
  INV_X1    g0582(.A(new_n689), .ZN(new_n783));
  AND4_X1   g0583(.A1(new_n581), .A2(new_n697), .A3(new_n698), .A4(new_n665), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n783), .B1(new_n784), .B2(new_n714), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n708), .A2(new_n709), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n719), .B1(new_n704), .B2(new_n705), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n786), .B1(new_n787), .B2(new_n709), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n732), .B1(new_n785), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(KEYINPUT29), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n779), .B1(new_n782), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n757), .B1(new_n791), .B2(G1), .ZN(G364));
  INV_X1    g0592(.A(new_n753), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n216), .A2(G13), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n275), .B1(new_n794), .B2(G45), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n738), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(G330), .B2(new_n737), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n307), .A2(new_n207), .ZN(new_n800));
  INV_X1    g0600(.A(G355), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n800), .A2(new_n801), .B1(G116), .B2(new_n207), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n294), .A2(new_n750), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(new_n272), .B2(new_n220), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n246), .A2(new_n272), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n802), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n215), .B1(G20), .B2(new_n283), .ZN(new_n808));
  NOR2_X1   g0608(.A1(G13), .A2(G33), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(G20), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT99), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n797), .B1(new_n807), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(G190), .A2(G200), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n815), .A2(G20), .A3(new_n285), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n307), .B1(new_n817), .B2(G329), .ZN(new_n818));
  INV_X1    g0618(.A(G311), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n216), .A2(new_n285), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n815), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n818), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n820), .A2(G190), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n823), .A2(G200), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(G322), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n823), .A2(new_n430), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n822), .B(new_n827), .C1(G326), .C2(new_n828), .ZN(new_n829));
  NOR4_X1   g0629(.A1(new_n216), .A2(new_n340), .A3(new_n430), .A4(G179), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G303), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n285), .A2(new_n430), .A3(G190), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(G20), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n831), .A2(new_n832), .B1(new_n564), .B2(new_n835), .ZN(new_n836));
  NOR4_X1   g0636(.A1(new_n216), .A2(new_n430), .A3(G179), .A4(G190), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n836), .B1(G283), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n820), .A2(new_n340), .A3(G200), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n839), .A2(KEYINPUT102), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n839), .A2(KEYINPUT102), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XOR2_X1   g0642(.A(KEYINPUT33), .B(G317), .Z(new_n843));
  OAI211_X1 g0643(.A(new_n829), .B(new_n838), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n828), .ZN(new_n845));
  INV_X1    g0645(.A(new_n837), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n845), .A2(new_n202), .B1(new_n225), .B2(new_n846), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n825), .A2(new_n298), .B1(new_n497), .B2(new_n835), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n842), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(G68), .ZN(new_n851));
  XOR2_X1   g0651(.A(KEYINPUT100), .B(G159), .Z(new_n852));
  NOR2_X1   g0652(.A1(new_n852), .A2(new_n816), .ZN(new_n853));
  XNOR2_X1  g0653(.A(KEYINPUT101), .B(KEYINPUT32), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n853), .B(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n307), .B1(new_n821), .B2(new_n223), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(G87), .B2(new_n830), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n849), .A2(new_n851), .A3(new_n855), .A4(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n844), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n814), .B1(new_n859), .B2(new_n808), .ZN(new_n860));
  INV_X1    g0660(.A(new_n811), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n860), .B1(new_n737), .B2(new_n861), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n799), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(G396));
  INV_X1    g0664(.A(KEYINPUT103), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n473), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n452), .A2(new_n471), .A3(KEYINPUT103), .A4(new_n472), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n471), .A2(new_n732), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n866), .A2(new_n475), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n473), .A2(new_n731), .ZN(new_n870));
  AND2_X1   g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n725), .B2(new_n732), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n872), .B(KEYINPUT104), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n866), .A2(new_n475), .A3(new_n867), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n731), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n787), .A2(KEYINPUT94), .A3(new_n709), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n724), .B(new_n876), .C1(new_n709), .C2(new_n708), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n875), .B1(new_n877), .B2(new_n785), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n779), .B1(new_n873), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n880), .A2(new_n797), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n873), .A2(new_n779), .A3(new_n879), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n797), .ZN(new_n884));
  INV_X1    g0684(.A(new_n808), .ZN(new_n885));
  INV_X1    g0685(.A(new_n852), .ZN(new_n886));
  INV_X1    g0686(.A(new_n821), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n828), .A2(G137), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(G143), .ZN(new_n889));
  INV_X1    g0689(.A(G150), .ZN(new_n890));
  OAI221_X1 g0690(.A(new_n888), .B1(new_n889), .B2(new_n825), .C1(new_n842), .C2(new_n890), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n891), .B(KEYINPUT34), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n257), .B1(G132), .B2(new_n817), .ZN(new_n893));
  OAI22_X1  g0693(.A1(new_n831), .A2(new_n202), .B1(new_n846), .B2(new_n299), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n894), .B1(G58), .B2(new_n834), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n892), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(G294), .ZN(new_n897));
  OAI22_X1  g0697(.A1(new_n897), .A2(new_n825), .B1(new_n845), .B2(new_n832), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n846), .A2(new_n262), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n850), .A2(G283), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n310), .B1(new_n816), .B2(new_n819), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n902), .B1(G116), .B2(new_n887), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n830), .A2(G107), .B1(new_n834), .B2(G97), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n900), .A2(new_n901), .A3(new_n903), .A4(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n885), .B1(new_n896), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n808), .A2(new_n809), .ZN(new_n907));
  AOI211_X1 g0707(.A(new_n884), .B(new_n906), .C1(new_n223), .C2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n869), .A2(new_n870), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n908), .B1(new_n909), .B2(new_n810), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n883), .A2(new_n910), .ZN(G384));
  OR2_X1    g0711(.A1(new_n642), .A2(KEYINPUT35), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n642), .A2(KEYINPUT35), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n912), .A2(G116), .A3(new_n217), .A4(new_n913), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n914), .B(KEYINPUT36), .Z(new_n915));
  OR3_X1    g0715(.A1(new_n219), .A2(new_n223), .A3(new_n300), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n202), .A2(G68), .ZN(new_n917));
  AOI211_X1 g0717(.A(new_n275), .B(G13), .C1(new_n916), .C2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT106), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n297), .A2(new_n303), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT105), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n335), .A2(KEYINPUT105), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n923), .A2(new_n305), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n333), .B1(new_n925), .B2(new_n336), .ZN(new_n926));
  INV_X1    g0726(.A(new_n730), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n920), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n316), .A2(new_n329), .A3(new_n342), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n305), .B1(new_n335), .B2(KEYINPUT105), .ZN(new_n930));
  AOI211_X1 g0730(.A(new_n922), .B(new_n306), .C1(new_n293), .C2(new_n296), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n336), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n329), .ZN(new_n933));
  INV_X1    g0733(.A(new_n287), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n929), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n933), .A2(KEYINPUT106), .A3(new_n730), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n928), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(KEYINPUT37), .ZN(new_n938));
  INV_X1    g0738(.A(new_n330), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n343), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n927), .B1(new_n316), .B2(new_n329), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n941), .A2(KEYINPUT37), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n938), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n928), .A2(new_n936), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n349), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n945), .A2(KEYINPUT38), .A3(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT38), .ZN(new_n949));
  INV_X1    g0749(.A(new_n941), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n939), .A2(new_n950), .A3(new_n343), .ZN(new_n951));
  OAI21_X1  g0751(.A(KEYINPUT37), .B1(new_n941), .B2(KEYINPUT107), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n951), .B(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n483), .A2(new_n484), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n950), .B1(new_n339), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n949), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n948), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n395), .A2(new_n732), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n396), .A2(new_n446), .A3(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n958), .B1(new_n396), .B2(new_n446), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n909), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n732), .A2(KEYINPUT31), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(new_n768), .B2(new_n763), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(new_n775), .B2(new_n777), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n957), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(KEYINPUT40), .ZN(new_n968));
  NOR2_X1   g0768(.A1(KEYINPUT109), .A2(KEYINPUT40), .ZN(new_n969));
  NOR3_X1   g0769(.A1(new_n962), .A2(new_n965), .A3(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n964), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n778), .A2(new_n971), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n395), .B(new_n732), .C1(new_n680), .C2(new_n382), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n871), .B1(new_n973), .B2(new_n959), .ZN(new_n974));
  AOI21_X1  g0774(.A(KEYINPUT109), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n970), .A2(new_n975), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n682), .A2(new_n339), .B1(new_n928), .B2(new_n936), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n943), .B1(new_n937), .B2(KEYINPUT37), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n949), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n948), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n976), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n968), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(new_n490), .B2(new_n972), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n967), .A2(KEYINPUT40), .B1(new_n976), .B2(new_n980), .ZN(new_n984));
  NOR3_X1   g0784(.A1(new_n984), .A2(new_n489), .A3(new_n965), .ZN(new_n985));
  NOR3_X1   g0785(.A1(new_n983), .A2(new_n985), .A3(new_n758), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n973), .A2(new_n959), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n866), .A2(new_n867), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n988), .A2(new_n732), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n987), .B1(new_n878), .B2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n991), .A2(new_n980), .B1(new_n481), .B2(new_n927), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT39), .ZN(new_n993));
  NOR3_X1   g0793(.A1(new_n977), .A2(new_n978), .A3(new_n949), .ZN(new_n994));
  AND2_X1   g0794(.A1(new_n951), .A2(new_n952), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n951), .A2(new_n952), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n955), .ZN(new_n998));
  AOI21_X1  g0798(.A(KEYINPUT38), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n993), .B1(new_n994), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n396), .A2(new_n732), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n948), .A2(new_n979), .A3(KEYINPUT39), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n992), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n686), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT108), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n790), .B1(new_n478), .B2(new_n488), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n877), .A2(new_n785), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n780), .B1(new_n1008), .B2(new_n731), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1006), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(KEYINPUT82), .B1(new_n349), .B2(new_n477), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n480), .A2(new_n487), .A3(new_n479), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n1011), .A2(new_n1012), .B1(KEYINPUT29), .B2(new_n789), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1013), .A2(new_n782), .A3(KEYINPUT108), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1005), .B1(new_n1010), .B2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1004), .B(new_n1015), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n986), .A2(new_n1016), .B1(new_n275), .B2(new_n794), .ZN(new_n1017));
  AND2_X1   g0817(.A1(new_n986), .A2(new_n1016), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n919), .B1(new_n1017), .B2(new_n1018), .ZN(G367));
  XOR2_X1   g0819(.A(KEYINPUT111), .B(KEYINPUT44), .Z(new_n1020));
  NAND2_X1  g0820(.A1(new_n673), .A2(new_n732), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n678), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n719), .A2(new_n732), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n746), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1020), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1020), .ZN(new_n1028));
  NOR3_X1   g0828(.A1(new_n1027), .A2(new_n746), .A3(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT45), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1027), .A2(KEYINPUT45), .A3(new_n746), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1030), .A2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n743), .A2(KEYINPUT112), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1036), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1038), .A2(new_n1030), .A3(new_n1034), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n744), .A2(new_n739), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n742), .B2(new_n744), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(new_n738), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1040), .A2(KEYINPUT113), .A3(new_n791), .A4(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT113), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n791), .A2(new_n1043), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1045), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1044), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n791), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT114), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n753), .B(KEYINPUT41), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1050), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n791), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n1044), .B2(new_n1048), .ZN(new_n1056));
  OAI21_X1  g0856(.A(KEYINPUT114), .B1(new_n1056), .B2(new_n1052), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1054), .A2(new_n795), .A3(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1024), .A2(new_n1041), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT42), .Z(new_n1060));
  NAND2_X1  g0860(.A1(new_n1027), .A2(new_n745), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n732), .B1(new_n1061), .B2(new_n676), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT43), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n714), .B1(new_n603), .B2(new_n731), .ZN(new_n1064));
  NOR3_X1   g0864(.A1(new_n689), .A2(new_n603), .A3(new_n731), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT110), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n1060), .A2(new_n1062), .B1(new_n1063), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(new_n1063), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1068), .B(new_n1069), .Z(new_n1070));
  NOR2_X1   g0870(.A1(new_n743), .A2(new_n1024), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1070), .B(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1058), .A2(new_n1072), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n1067), .A2(new_n811), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n812), .B1(new_n207), .B2(new_n588), .C1(new_n242), .C2(new_n804), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n889), .A2(new_n845), .B1(new_n825), .B2(new_n890), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(G58), .B2(new_n830), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n850), .A2(new_n886), .ZN(new_n1078));
  INV_X1    g0878(.A(G137), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n307), .B1(new_n816), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(G50), .B2(new_n887), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n837), .A2(G77), .B1(new_n834), .B2(G68), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1077), .A2(new_n1078), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(G317), .ZN(new_n1084));
  INV_X1    g0884(.A(G283), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n257), .B1(new_n1084), .B2(new_n816), .C1(new_n1085), .C2(new_n821), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n564), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1086), .B1(new_n850), .B2(new_n1087), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n824), .A2(G303), .B1(G107), .B2(new_n834), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n846), .A2(new_n497), .ZN(new_n1090));
  XOR2_X1   g0890(.A(KEYINPUT115), .B(G311), .Z(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1090), .B1(new_n828), .B2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1088), .A2(new_n1089), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n830), .A2(G116), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT46), .Z(new_n1096));
  OAI21_X1  g0896(.A(new_n1083), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT47), .Z(new_n1098));
  OAI211_X1 g0898(.A(new_n797), .B(new_n1075), .C1(new_n1098), .C2(new_n885), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1074), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1073), .A2(new_n1101), .ZN(G387));
  NAND2_X1  g0902(.A1(new_n1043), .A2(new_n796), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n828), .A2(G322), .B1(new_n887), .B2(G303), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n1104), .B1(new_n1084), .B2(new_n825), .C1(new_n842), .C2(new_n1091), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT48), .ZN(new_n1106));
  OR2_X1    g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n830), .A2(new_n1087), .B1(new_n834), .B2(G283), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT117), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1107), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT49), .ZN(new_n1112));
  OR2_X1    g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n846), .A2(new_n493), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n294), .B(new_n1115), .C1(G326), .C2(new_n817), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1113), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(G159), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n202), .A2(new_n825), .B1(new_n845), .B2(new_n1118), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n1090), .B(new_n1119), .C1(G77), .C2(new_n830), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n626), .A2(new_n627), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n834), .ZN(new_n1122));
  OR2_X1    g0922(.A1(new_n842), .A2(new_n322), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n821), .A2(new_n299), .B1(new_n816), .B2(new_n890), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1124), .A2(new_n257), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1120), .A2(new_n1122), .A3(new_n1123), .A4(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1117), .A2(new_n1126), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n1127), .A2(KEYINPUT118), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1127), .A2(KEYINPUT118), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n1128), .A2(new_n1129), .A3(new_n885), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n455), .A2(G50), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT50), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n272), .B1(new_n299), .B2(new_n223), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n754), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT116), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1133), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1132), .B(new_n1136), .C1(new_n1135), .C2(new_n1134), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1137), .B(new_n803), .C1(new_n239), .C2(new_n272), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n1138), .B1(G107), .B2(new_n207), .C1(new_n754), .C2(new_n800), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n813), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n884), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1141), .B1(new_n742), .B2(new_n861), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1046), .A2(new_n793), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n791), .A2(new_n1043), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1103), .B1(new_n1130), .B2(new_n1142), .C1(new_n1143), .C2(new_n1144), .ZN(G393));
  XOR2_X1   g0945(.A(new_n1035), .B(new_n743), .Z(new_n1146));
  AOI21_X1  g0946(.A(new_n753), .B1(new_n1146), .B2(new_n1046), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1049), .A2(new_n1147), .ZN(new_n1148));
  OR2_X1    g0948(.A1(new_n1146), .A2(new_n795), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n812), .B1(new_n497), .B2(new_n207), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n804), .A2(new_n249), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n797), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(G311), .A2(new_n824), .B1(new_n828), .B2(G317), .ZN(new_n1153));
  XOR2_X1   g0953(.A(new_n1153), .B(KEYINPUT52), .Z(new_n1154));
  OAI221_X1 g0954(.A(new_n310), .B1(new_n816), .B2(new_n826), .C1(new_n821), .C2(new_n897), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(new_n850), .B2(G303), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n831), .A2(new_n1085), .B1(new_n846), .B2(new_n225), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(G116), .B2(new_n834), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1154), .A2(new_n1156), .A3(new_n1158), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(G150), .A2(new_n828), .B1(new_n824), .B2(G159), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT51), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n835), .A2(new_n223), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1162), .B(new_n899), .C1(G68), .C2(new_n830), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n821), .A2(new_n455), .B1(new_n816), .B2(new_n889), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1164), .A2(new_n257), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1163), .B(new_n1165), .C1(new_n202), .C2(new_n842), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1159), .B1(new_n1161), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1152), .B1(new_n1167), .B2(new_n808), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n1027), .B2(new_n861), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n1148), .A2(new_n1149), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(G390));
  INV_X1    g0971(.A(KEYINPUT119), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n965), .A2(new_n758), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n974), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1001), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n1000), .A2(new_n1002), .B1(new_n1176), .B2(new_n990), .ZN(new_n1177));
  AND2_X1   g0977(.A1(new_n708), .A2(new_n709), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n723), .B2(KEYINPUT26), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n731), .B(new_n874), .C1(new_n1179), .C2(new_n707), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n989), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  AOI221_X4 g0982(.A(new_n1001), .B1(new_n1182), .B2(new_n987), .C1(new_n948), .C2(new_n956), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1172), .B(new_n1175), .C1(new_n1177), .C2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n990), .A2(new_n1176), .ZN(new_n1185));
  AND3_X1   g0985(.A1(new_n948), .A2(new_n979), .A3(KEYINPUT39), .ZN(new_n1186));
  AOI21_X1  g0986(.A(KEYINPUT39), .B1(new_n948), .B2(new_n956), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1185), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n987), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1182), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n957), .B(new_n1176), .C1(new_n1189), .C2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n779), .A2(new_n909), .A3(new_n987), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1188), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1184), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1188), .A2(new_n1191), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1172), .B1(new_n1195), .B2(new_n1175), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n796), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(new_n809), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n842), .A2(new_n225), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n310), .B1(new_n816), .B2(new_n897), .C1(new_n821), .C2(new_n497), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n831), .A2(new_n262), .B1(new_n846), .B2(new_n299), .ZN(new_n1203));
  NOR3_X1   g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1162), .B1(G116), .B2(new_n824), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1204), .B(new_n1205), .C1(new_n1085), .C2(new_n845), .ZN(new_n1206));
  INV_X1    g1006(.A(G125), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(KEYINPUT54), .B(G143), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n307), .B1(new_n816), .B2(new_n1207), .C1(new_n821), .C2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n850), .B2(G137), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n830), .A2(G150), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1211), .B(KEYINPUT53), .Z(new_n1212));
  AOI22_X1  g1012(.A1(new_n824), .A2(G132), .B1(G159), .B2(new_n834), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n828), .A2(G128), .B1(G50), .B2(new_n837), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1210), .A2(new_n1212), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n885), .B1(new_n1206), .B2(new_n1215), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n884), .B(new_n1216), .C1(new_n322), .C2(new_n907), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1200), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n490), .A2(new_n1173), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1013), .A2(new_n782), .A3(KEYINPUT108), .ZN(new_n1220));
  AOI21_X1  g1020(.A(KEYINPUT108), .B1(new_n1013), .B2(new_n782), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n686), .B(new_n1219), .C1(new_n1220), .C2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT120), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1015), .A2(KEYINPUT120), .A3(new_n1219), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n779), .A2(new_n909), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1174), .B1(new_n1227), .B2(new_n987), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n878), .A2(new_n989), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1228), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1173), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1189), .B1(new_n1232), .B2(new_n871), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1233), .A2(new_n1190), .A3(new_n1192), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1231), .A2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1224), .A2(new_n1225), .A3(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n1194), .B2(new_n1196), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n793), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1183), .B1(new_n1199), .B2(new_n1185), .ZN(new_n1239));
  OAI21_X1  g1039(.A(KEYINPUT119), .B1(new_n1239), .B2(new_n1174), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1240), .A2(new_n1193), .A3(new_n1184), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1241), .A2(new_n1236), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1198), .B(new_n1218), .C1(new_n1238), .C2(new_n1242), .ZN(G378));
  NAND2_X1  g1043(.A1(new_n403), .A2(new_n730), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(new_n440), .B(new_n1244), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1245), .B(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(new_n982), .B2(G330), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n984), .A2(new_n758), .A3(new_n1247), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1004), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1247), .B1(new_n984), .B2(new_n758), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1004), .ZN(new_n1253));
  AND2_X1   g1053(.A1(new_n976), .A2(new_n980), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT40), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(new_n957), .B2(new_n966), .ZN(new_n1256));
  OAI211_X1 g1056(.A(G330), .B(new_n1248), .C1(new_n1254), .C2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1252), .A2(new_n1253), .A3(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1251), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1247), .A2(new_n809), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n907), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n797), .B1(G50), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n257), .A2(new_n748), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n835), .A2(new_n299), .B1(new_n1085), .B2(new_n816), .ZN(new_n1264));
  AOI211_X1 g1064(.A(new_n1263), .B(new_n1264), .C1(new_n850), .C2(G97), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1121), .A2(new_n887), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n828), .A2(G116), .B1(G77), .B2(new_n830), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n824), .A2(G107), .B1(G58), .B2(new_n837), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1265), .A2(new_n1266), .A3(new_n1267), .A4(new_n1268), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(new_n1269), .B(KEYINPUT121), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT58), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1263), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1208), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n830), .A2(new_n1275), .B1(new_n834), .B2(G150), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n845), .B2(new_n1207), .ZN(new_n1277));
  INV_X1    g1077(.A(G128), .ZN(new_n1278));
  OAI22_X1  g1078(.A1(new_n825), .A2(new_n1278), .B1(new_n821), .B2(new_n1079), .ZN(new_n1279));
  AOI211_X1 g1079(.A(new_n1277), .B(new_n1279), .C1(G132), .C2(new_n850), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(new_n1280), .B(KEYINPUT59), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1282), .A2(KEYINPUT122), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(KEYINPUT122), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n886), .A2(new_n837), .ZN(new_n1285));
  AOI211_X1 g1085(.A(G33), .B(G41), .C1(new_n817), .C2(G124), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1284), .A2(new_n1285), .A3(new_n1286), .ZN(new_n1287));
  OAI221_X1 g1087(.A(new_n1274), .B1(new_n1271), .B2(new_n1270), .C1(new_n1283), .C2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1262), .B1(new_n1288), .B2(new_n808), .ZN(new_n1289));
  AOI22_X1  g1089(.A1(new_n1259), .A2(new_n796), .B1(new_n1260), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1291), .B1(new_n1197), .B2(new_n1235), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1252), .A2(new_n1253), .A3(new_n1257), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1253), .B1(new_n1252), .B2(new_n1257), .ZN(new_n1294));
  OAI21_X1  g1094(.A(KEYINPUT57), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n793), .B1(new_n1292), .B2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1291), .ZN(new_n1297));
  AND2_X1   g1097(.A1(new_n1231), .A2(new_n1234), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1297), .B1(new_n1241), .B2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(KEYINPUT57), .B1(new_n1299), .B2(new_n1259), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1290), .B1(new_n1296), .B2(new_n1300), .ZN(G375));
  OAI21_X1  g1101(.A(new_n797), .B1(G68), .B2(new_n1261), .ZN(new_n1302));
  OAI22_X1  g1102(.A1(new_n825), .A2(new_n1079), .B1(new_n202), .B2(new_n835), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1303), .B1(G132), .B2(new_n828), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n850), .A2(new_n1275), .ZN(new_n1305));
  OAI22_X1  g1105(.A1(new_n821), .A2(new_n890), .B1(new_n816), .B2(new_n1278), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1306), .A2(new_n257), .ZN(new_n1307));
  AOI22_X1  g1107(.A1(new_n830), .A2(G159), .B1(new_n837), .B2(G58), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1304), .A2(new_n1305), .A3(new_n1307), .A4(new_n1308), .ZN(new_n1309));
  OAI22_X1  g1109(.A1(new_n845), .A2(new_n897), .B1(new_n821), .B2(new_n225), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1310), .B1(new_n850), .B2(G116), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(new_n1311), .B(KEYINPUT124), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n310), .B1(new_n816), .B2(new_n832), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1313), .B1(G77), .B2(new_n837), .ZN(new_n1314));
  AOI22_X1  g1114(.A1(new_n824), .A2(G283), .B1(G97), .B2(new_n830), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1122), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1309), .B1(new_n1312), .B2(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1302), .B1(new_n1317), .B2(new_n808), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1318), .B1(new_n987), .B2(new_n810), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1319), .B1(new_n1298), .B2(new_n795), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT125), .ZN(new_n1321));
  XNOR2_X1  g1121(.A(new_n1320), .B(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT123), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1291), .A2(new_n1298), .ZN(new_n1324));
  AND3_X1   g1124(.A1(new_n1324), .A2(new_n1053), .A3(new_n1236), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1322), .B1(new_n1323), .B2(new_n1325), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1326), .B1(new_n1323), .B2(new_n1325), .ZN(G381));
  OAI21_X1  g1127(.A(new_n1218), .B1(new_n1241), .B2(new_n795), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1242), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n753), .B1(new_n1241), .B2(new_n1236), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1328), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1331));
  NOR3_X1   g1131(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1331), .A2(new_n1170), .A3(new_n1332), .ZN(new_n1333));
  OR4_X1    g1133(.A1(G387), .A2(G381), .A3(G375), .A4(new_n1333), .ZN(G407));
  OR2_X1    g1134(.A1(G378), .A2(G343), .ZN(new_n1335));
  OAI211_X1 g1135(.A(G407), .B(G213), .C1(G375), .C2(new_n1335), .ZN(G409));
  OAI211_X1 g1136(.A(G378), .B(new_n1290), .C1(new_n1296), .C2(new_n1300), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1299), .A2(new_n1053), .A3(new_n1259), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1338), .A2(new_n1290), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1339), .A2(new_n1331), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1337), .A2(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1322), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1235), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n753), .B1(new_n1343), .B2(KEYINPUT60), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1343), .B1(KEYINPUT60), .B2(new_n1236), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1344), .B1(new_n1345), .B2(KEYINPUT126), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1236), .A2(KEYINPUT60), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1347), .A2(KEYINPUT126), .A3(new_n1324), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1348), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1342), .B1(new_n1346), .B2(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(G384), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1347), .A2(new_n1324), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT126), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1353), .A2(new_n1354), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1355), .A2(new_n1348), .A3(new_n1344), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1356), .A2(G384), .A3(new_n1342), .ZN(new_n1357));
  INV_X1    g1157(.A(G213), .ZN(new_n1358));
  NOR2_X1   g1158(.A1(new_n1358), .A2(G343), .ZN(new_n1359));
  INV_X1    g1159(.A(new_n1359), .ZN(new_n1360));
  NAND4_X1  g1160(.A1(new_n1341), .A2(new_n1352), .A3(new_n1357), .A4(new_n1360), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1361), .A2(KEYINPUT62), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1341), .A2(new_n1360), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1359), .A2(G2897), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1352), .A2(new_n1357), .A3(new_n1364), .ZN(new_n1365));
  INV_X1    g1165(.A(new_n1364), .ZN(new_n1366));
  NOR2_X1   g1166(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1367));
  AOI21_X1  g1167(.A(KEYINPUT120), .B1(new_n1015), .B2(new_n1219), .ZN(new_n1368));
  OAI211_X1 g1168(.A(KEYINPUT60), .B(new_n1298), .C1(new_n1367), .C2(new_n1368), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1369), .A2(new_n793), .ZN(new_n1370));
  AOI21_X1  g1170(.A(new_n1370), .B1(new_n1353), .B2(new_n1354), .ZN(new_n1371));
  AOI211_X1 g1171(.A(new_n1351), .B(new_n1322), .C1(new_n1371), .C2(new_n1348), .ZN(new_n1372));
  AOI21_X1  g1172(.A(G384), .B1(new_n1356), .B2(new_n1342), .ZN(new_n1373));
  OAI21_X1  g1173(.A(new_n1366), .B1(new_n1372), .B2(new_n1373), .ZN(new_n1374));
  NAND3_X1  g1174(.A1(new_n1363), .A2(new_n1365), .A3(new_n1374), .ZN(new_n1375));
  INV_X1    g1175(.A(KEYINPUT61), .ZN(new_n1376));
  AOI21_X1  g1176(.A(new_n1359), .B1(new_n1337), .B2(new_n1340), .ZN(new_n1377));
  NOR2_X1   g1177(.A1(new_n1372), .A2(new_n1373), .ZN(new_n1378));
  INV_X1    g1178(.A(KEYINPUT62), .ZN(new_n1379));
  NAND3_X1  g1179(.A1(new_n1377), .A2(new_n1378), .A3(new_n1379), .ZN(new_n1380));
  NAND4_X1  g1180(.A1(new_n1362), .A2(new_n1375), .A3(new_n1376), .A4(new_n1380), .ZN(new_n1381));
  NAND2_X1  g1181(.A1(G387), .A2(new_n1170), .ZN(new_n1382));
  XNOR2_X1  g1182(.A(G393), .B(new_n863), .ZN(new_n1383));
  NAND3_X1  g1183(.A1(new_n1073), .A2(G390), .A3(new_n1101), .ZN(new_n1384));
  NAND3_X1  g1184(.A1(new_n1382), .A2(new_n1383), .A3(new_n1384), .ZN(new_n1385));
  INV_X1    g1185(.A(new_n1383), .ZN(new_n1386));
  AOI21_X1  g1186(.A(G390), .B1(new_n1073), .B2(new_n1101), .ZN(new_n1387));
  AOI211_X1 g1187(.A(new_n1100), .B(new_n1170), .C1(new_n1058), .C2(new_n1072), .ZN(new_n1388));
  OAI21_X1  g1188(.A(new_n1386), .B1(new_n1387), .B2(new_n1388), .ZN(new_n1389));
  AND2_X1   g1189(.A1(new_n1385), .A2(new_n1389), .ZN(new_n1390));
  INV_X1    g1190(.A(new_n1390), .ZN(new_n1391));
  NAND2_X1  g1191(.A1(new_n1381), .A2(new_n1391), .ZN(new_n1392));
  NAND2_X1  g1192(.A1(new_n1352), .A2(new_n1357), .ZN(new_n1393));
  AOI22_X1  g1193(.A1(new_n1393), .A2(new_n1366), .B1(new_n1341), .B2(new_n1360), .ZN(new_n1394));
  AOI21_X1  g1194(.A(KEYINPUT61), .B1(new_n1394), .B2(new_n1365), .ZN(new_n1395));
  NAND3_X1  g1195(.A1(new_n1377), .A2(new_n1378), .A3(KEYINPUT63), .ZN(new_n1396));
  AND2_X1   g1196(.A1(new_n1396), .A2(new_n1390), .ZN(new_n1397));
  INV_X1    g1197(.A(KEYINPUT63), .ZN(new_n1398));
  NAND2_X1  g1198(.A1(new_n1361), .A2(new_n1398), .ZN(new_n1399));
  NAND3_X1  g1199(.A1(new_n1395), .A2(new_n1397), .A3(new_n1399), .ZN(new_n1400));
  NAND2_X1  g1200(.A1(new_n1392), .A2(new_n1400), .ZN(G405));
  NAND2_X1  g1201(.A1(G375), .A2(new_n1331), .ZN(new_n1402));
  NAND2_X1  g1202(.A1(new_n1402), .A2(new_n1337), .ZN(new_n1403));
  NAND2_X1  g1203(.A1(new_n1403), .A2(new_n1378), .ZN(new_n1404));
  INV_X1    g1204(.A(new_n1404), .ZN(new_n1405));
  NOR2_X1   g1205(.A1(new_n1403), .A2(new_n1378), .ZN(new_n1406));
  OAI21_X1  g1206(.A(new_n1391), .B1(new_n1405), .B2(new_n1406), .ZN(new_n1407));
  INV_X1    g1207(.A(new_n1406), .ZN(new_n1408));
  NAND3_X1  g1208(.A1(new_n1408), .A2(new_n1390), .A3(new_n1404), .ZN(new_n1409));
  NAND2_X1  g1209(.A1(new_n1407), .A2(new_n1409), .ZN(G402));
endmodule


