//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 0 1 1 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 1 1 0 0 0 1 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 1 0 1 0 0 0 0 1 0 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1309, new_n1310, new_n1312, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1373, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378, new_n1379;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT64), .Z(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G68), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n217));
  INV_X1    g0017(.A(G77), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  INV_X1    g0019(.A(G264), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n206), .C2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n210), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  OR2_X1    g0022(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  OAI21_X1  g0023(.A(G50), .B1(G58), .B2(G68), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT65), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  OR2_X1    g0029(.A1(new_n225), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n210), .A2(G13), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n231), .B(G250), .C1(G257), .C2(G264), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT0), .ZN(new_n233));
  NAND3_X1  g0033(.A1(new_n223), .A2(new_n230), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G50), .B(G68), .Z(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G1), .A3(G13), .ZN(new_n252));
  INV_X1    g0052(.A(G1), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n253), .B1(G41), .B2(G45), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n252), .A2(G232), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT81), .ZN(new_n256));
  INV_X1    g0056(.A(G41), .ZN(new_n257));
  INV_X1    g0057(.A(G45), .ZN(new_n258));
  AOI21_X1  g0058(.A(G1), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(new_n252), .A3(G274), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT81), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n252), .A2(new_n254), .A3(new_n261), .A4(G232), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n256), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  AND4_X1   g0063(.A1(KEYINPUT67), .A2(new_n251), .A3(G1), .A4(G13), .ZN(new_n264));
  AND2_X1   g0064(.A1(G1), .A2(G13), .ZN(new_n265));
  AOI21_X1  g0065(.A(KEYINPUT67), .B1(new_n265), .B2(new_n251), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT78), .ZN(new_n268));
  INV_X1    g0068(.A(G33), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n268), .B1(new_n269), .B2(KEYINPUT3), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(KEYINPUT3), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n272), .A2(KEYINPUT78), .A3(G33), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n270), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G226), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G1698), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n276), .B1(G223), .B2(G1698), .ZN(new_n277));
  OAI22_X1  g0077(.A1(new_n274), .A2(new_n277), .B1(new_n269), .B2(new_n214), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n263), .A2(KEYINPUT82), .B1(new_n267), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT82), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n256), .A2(new_n280), .A3(new_n260), .A4(new_n262), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(G179), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n263), .A2(KEYINPUT82), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n278), .A2(new_n267), .ZN(new_n284));
  AND3_X1   g0084(.A1(new_n283), .A2(new_n281), .A3(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G169), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n282), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G58), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n288), .A2(new_n212), .ZN(new_n289));
  OAI21_X1  g0089(.A(G20), .B1(new_n289), .B2(new_n201), .ZN(new_n290));
  NOR2_X1   g0090(.A1(G20), .A2(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G159), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT79), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT7), .ZN(new_n296));
  AOI21_X1  g0096(.A(G20), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(KEYINPUT79), .A2(KEYINPUT7), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n274), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G68), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n298), .B1(new_n274), .B2(new_n297), .ZN(new_n301));
  OAI211_X1 g0101(.A(KEYINPUT16), .B(new_n294), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT69), .ZN(new_n304));
  AND3_X1   g0104(.A1(new_n303), .A2(new_n304), .A3(new_n226), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n304), .B1(new_n303), .B2(new_n226), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT16), .ZN(new_n308));
  XNOR2_X1  g0108(.A(KEYINPUT3), .B(G33), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n296), .B1(new_n309), .B2(G20), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n272), .A2(G33), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n271), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n312), .A2(KEYINPUT7), .A3(new_n227), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n212), .B1(new_n310), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n308), .B1(new_n314), .B2(new_n293), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n302), .A2(new_n307), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT8), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(new_n288), .B2(KEYINPUT70), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT70), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n319), .A2(KEYINPUT8), .A3(G58), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n253), .A2(G13), .A3(G20), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n322), .B1(new_n305), .B2(new_n306), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n253), .A2(G20), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n318), .A2(new_n320), .A3(new_n326), .ZN(new_n327));
  OAI211_X1 g0127(.A(KEYINPUT80), .B(new_n324), .C1(new_n325), .C2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n303), .A2(new_n226), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT69), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n303), .A2(new_n304), .A3(new_n226), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n327), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n333), .A2(new_n334), .A3(new_n322), .ZN(new_n335));
  AOI21_X1  g0135(.A(KEYINPUT80), .B1(new_n335), .B2(new_n324), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n329), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n316), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n287), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT18), .ZN(new_n340));
  INV_X1    g0140(.A(G190), .ZN(new_n341));
  AND4_X1   g0141(.A1(new_n341), .A2(new_n283), .A3(new_n281), .A4(new_n284), .ZN(new_n342));
  AOI21_X1  g0142(.A(G200), .B1(new_n279), .B2(new_n281), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n337), .B(new_n316), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT17), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT18), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n287), .A2(new_n338), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n279), .A2(new_n341), .A3(new_n281), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(new_n285), .B2(G200), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n350), .A2(KEYINPUT17), .A3(new_n337), .A4(new_n316), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n340), .A2(new_n346), .A3(new_n348), .A4(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n260), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n252), .A2(new_n254), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n354), .B1(G226), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n309), .A2(G1698), .ZN(new_n358));
  INV_X1    g0158(.A(G223), .ZN(new_n359));
  OAI22_X1  g0159(.A1(new_n358), .A2(new_n359), .B1(new_n218), .B2(new_n309), .ZN(new_n360));
  INV_X1    g0160(.A(G1698), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n309), .A2(G222), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT66), .ZN(new_n363));
  OR2_X1    g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n363), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n360), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT67), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n252), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n265), .A2(KEYINPUT67), .A3(new_n251), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n357), .B1(new_n366), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(KEYINPUT68), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT68), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n373), .B(new_n357), .C1(new_n366), .C2(new_n370), .ZN(new_n374));
  AND3_X1   g0174(.A1(new_n372), .A2(new_n286), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(G179), .B1(new_n372), .B2(new_n374), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n326), .A2(G50), .ZN(new_n377));
  XNOR2_X1  g0177(.A(new_n377), .B(KEYINPUT71), .ZN(new_n378));
  OR2_X1    g0178(.A1(new_n378), .A2(new_n325), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n291), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n227), .A2(G33), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n380), .B1(new_n321), .B2(new_n381), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n382), .A2(new_n307), .B1(new_n202), .B2(new_n323), .ZN(new_n383));
  AND2_X1   g0183(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  NOR3_X1   g0184(.A1(new_n375), .A2(new_n376), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n372), .A2(G200), .A3(new_n374), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n379), .A2(new_n383), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n387), .B(KEYINPUT9), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n341), .B1(new_n372), .B2(new_n374), .ZN(new_n390));
  OAI21_X1  g0190(.A(KEYINPUT10), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n390), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT10), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n392), .A2(new_n393), .A3(new_n386), .A4(new_n388), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n385), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n260), .B1(new_n219), .B2(new_n355), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n309), .A2(G232), .A3(new_n361), .ZN(new_n397));
  OAI221_X1 g0197(.A(new_n397), .B1(new_n206), .B2(new_n309), .C1(new_n358), .C2(new_n213), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n396), .B1(new_n398), .B2(new_n267), .ZN(new_n399));
  INV_X1    g0199(.A(G200), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT72), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n398), .A2(new_n267), .ZN(new_n402));
  INV_X1    g0202(.A(new_n396), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n401), .B1(new_n341), .B2(new_n404), .ZN(new_n405));
  XNOR2_X1  g0205(.A(KEYINPUT8), .B(G58), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n407), .A2(new_n291), .B1(G20), .B2(G77), .ZN(new_n408));
  XNOR2_X1  g0208(.A(KEYINPUT15), .B(G87), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n408), .B1(new_n381), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n307), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n333), .A2(G77), .A3(new_n322), .A4(new_n326), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n323), .A2(new_n218), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT73), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n411), .A2(KEYINPUT73), .A3(new_n412), .A4(new_n413), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n399), .A2(KEYINPUT72), .A3(G190), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n405), .A2(new_n416), .A3(new_n417), .A4(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n404), .A2(new_n286), .ZN(new_n420));
  INV_X1    g0220(.A(G179), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n399), .A2(new_n421), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n416), .A2(new_n417), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n419), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT74), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT74), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n419), .A2(new_n425), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(G33), .A2(G97), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n275), .A2(new_n361), .ZN(new_n432));
  INV_X1    g0232(.A(G232), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(G1698), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n431), .B1(new_n312), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n267), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n252), .A2(G238), .A3(new_n254), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n260), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT13), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n437), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n441), .B1(new_n437), .B2(new_n440), .ZN(new_n443));
  OAI21_X1  g0243(.A(G169), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT14), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n437), .A2(new_n440), .A3(new_n441), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n439), .B1(new_n267), .B2(new_n436), .ZN(new_n447));
  OAI21_X1  g0247(.A(KEYINPUT13), .B1(new_n447), .B2(KEYINPUT75), .ZN(new_n448));
  INV_X1    g0248(.A(new_n431), .ZN(new_n449));
  NOR2_X1   g0249(.A1(G226), .A2(G1698), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n450), .B1(new_n433), .B2(G1698), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n449), .B1(new_n451), .B2(new_n309), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n260), .B(new_n438), .C1(new_n452), .C2(new_n370), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT75), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI211_X1 g0255(.A(G179), .B(new_n446), .C1(new_n448), .C2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT14), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n457), .B(G169), .C1(new_n442), .C2(new_n443), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n445), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n212), .B1(new_n253), .B2(G20), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n333), .A2(new_n322), .A3(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n253), .A2(new_n212), .A3(G13), .A4(G20), .ZN(new_n462));
  XNOR2_X1  g0262(.A(new_n462), .B(KEYINPUT12), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n461), .A2(KEYINPUT76), .A3(new_n463), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n291), .A2(G50), .B1(G20), .B2(new_n212), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n465), .B1(new_n218), .B2(new_n381), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n307), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT11), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n307), .A2(new_n466), .A3(KEYINPUT11), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n464), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT76), .B1(new_n461), .B2(new_n463), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n459), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT77), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n453), .A2(KEYINPUT13), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n400), .B1(new_n477), .B2(new_n446), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n441), .B1(new_n453), .B2(new_n454), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n447), .A2(KEYINPUT75), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n442), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n478), .B1(new_n481), .B2(G190), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n476), .B1(new_n482), .B2(new_n473), .ZN(new_n483));
  OAI211_X1 g0283(.A(G190), .B(new_n446), .C1(new_n448), .C2(new_n455), .ZN(new_n484));
  OAI21_X1  g0284(.A(G200), .B1(new_n442), .B2(new_n443), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n484), .A2(new_n473), .A3(new_n476), .A4(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n475), .B1(new_n483), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  AND4_X1   g0289(.A1(new_n353), .A2(new_n395), .A3(new_n430), .A4(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n271), .A2(new_n311), .A3(G250), .A4(G1698), .ZN(new_n492));
  AND2_X1   g0292(.A1(KEYINPUT4), .A2(G244), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n271), .A2(new_n311), .A3(new_n493), .A4(new_n361), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G33), .A2(G283), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n492), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n219), .A2(G1698), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n270), .A2(new_n273), .A3(new_n497), .A4(new_n271), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n370), .B1(new_n496), .B2(new_n500), .ZN(new_n501));
  XNOR2_X1  g0301(.A(KEYINPUT5), .B(G41), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n258), .A2(G1), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n502), .A2(new_n503), .B1(new_n265), .B2(new_n251), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G257), .ZN(new_n505));
  INV_X1    g0305(.A(G274), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n506), .B1(new_n265), .B2(new_n251), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n507), .A2(new_n502), .A3(new_n503), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT84), .ZN(new_n510));
  NOR3_X1   g0310(.A1(new_n501), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n498), .A2(new_n499), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n492), .A2(new_n494), .A3(new_n495), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n267), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n252), .A2(G274), .ZN(new_n515));
  NAND2_X1  g0315(.A1(KEYINPUT5), .A2(G41), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(KEYINPUT5), .A2(G41), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n503), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n520), .B1(G257), .B2(new_n504), .ZN(new_n521));
  AOI21_X1  g0321(.A(KEYINPUT84), .B1(new_n514), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n286), .B1(new_n511), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n514), .A2(new_n521), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n524), .A2(G179), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n291), .A2(G77), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT6), .ZN(new_n528));
  NOR3_X1   g0328(.A1(new_n528), .A2(new_n205), .A3(G107), .ZN(new_n529));
  XNOR2_X1  g0329(.A(G97), .B(G107), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n529), .B1(new_n530), .B2(new_n528), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n527), .B1(new_n531), .B2(new_n227), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n206), .B1(new_n310), .B2(new_n313), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n307), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n253), .A2(G33), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n322), .B(new_n535), .C1(new_n305), .C2(new_n306), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(G97), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n322), .A2(G97), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n534), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n523), .A2(new_n526), .A3(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT83), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n510), .B1(new_n501), .B2(new_n509), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n514), .A2(KEYINPUT84), .A3(new_n521), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(G190), .A3(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n534), .A2(KEYINPUT83), .A3(new_n538), .A4(new_n540), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n524), .A2(G200), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n544), .A2(new_n547), .A3(new_n548), .A4(new_n549), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n270), .A2(new_n271), .A3(new_n273), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT22), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n552), .A2(new_n214), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n551), .A2(new_n227), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n227), .A2(G87), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n552), .B1(new_n312), .B2(new_n555), .ZN(new_n556));
  OR2_X1    g0356(.A1(KEYINPUT86), .A2(G116), .ZN(new_n557));
  NAND2_X1  g0357(.A1(KEYINPUT86), .A2(G116), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n269), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT23), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n227), .B2(G107), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n559), .A2(new_n227), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n554), .A2(new_n556), .A3(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT24), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n333), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n554), .A2(new_n563), .A3(KEYINPUT24), .A4(new_n556), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n536), .A2(new_n206), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT25), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(KEYINPUT90), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT90), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT25), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT91), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n322), .A2(G107), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT91), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n570), .A2(new_n572), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n574), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  XNOR2_X1  g0378(.A(KEYINPUT90), .B(KEYINPUT25), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n579), .B(new_n576), .C1(G107), .C2(new_n322), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(KEYINPUT92), .B1(new_n568), .B2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n333), .A2(G107), .A3(new_n322), .A4(new_n535), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT92), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n583), .A2(new_n584), .A3(new_n580), .A4(new_n578), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n566), .A2(new_n567), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n215), .A2(new_n361), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(G257), .B2(new_n361), .ZN(new_n588));
  INV_X1    g0388(.A(G294), .ZN(new_n589));
  OAI22_X1  g0389(.A1(new_n274), .A2(new_n588), .B1(new_n269), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n590), .A2(new_n267), .B1(G264), .B2(new_n504), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n591), .A2(new_n341), .A3(new_n508), .ZN(new_n592));
  AOI21_X1  g0392(.A(G200), .B1(new_n591), .B2(new_n508), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT93), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AOI211_X1 g0395(.A(KEYINPUT93), .B(G200), .C1(new_n591), .C2(new_n508), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n586), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(G169), .B1(new_n591), .B2(new_n508), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n591), .A2(new_n508), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n598), .B1(new_n600), .B2(new_n421), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n582), .A2(new_n585), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n564), .A2(new_n565), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n603), .A2(new_n307), .A3(new_n567), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n542), .A2(new_n550), .A3(new_n597), .A4(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n519), .A2(G270), .A3(new_n252), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n608), .A2(new_n508), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n220), .A2(G1698), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(G257), .B2(G1698), .ZN(new_n611));
  INV_X1    g0411(.A(G303), .ZN(new_n612));
  OAI22_X1  g0412(.A1(new_n274), .A2(new_n611), .B1(new_n612), .B2(new_n309), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n267), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n286), .B1(new_n609), .B2(new_n614), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n495), .B(new_n227), .C1(G33), .C2(new_n205), .ZN(new_n616));
  XNOR2_X1  g0416(.A(KEYINPUT86), .B(G116), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n330), .B(new_n616), .C1(new_n617), .C2(new_n227), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT20), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n616), .A2(new_n330), .ZN(new_n621));
  INV_X1    g0421(.A(new_n558), .ZN(new_n622));
  NOR2_X1   g0422(.A1(KEYINPUT86), .A2(G116), .ZN(new_n623));
  NOR3_X1   g0423(.A1(new_n622), .A2(new_n623), .A3(new_n227), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n619), .B1(new_n621), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(KEYINPUT89), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT89), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n618), .A2(new_n627), .A3(new_n619), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n620), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(G116), .ZN(new_n630));
  OAI22_X1  g0430(.A1(new_n536), .A2(new_n630), .B1(new_n322), .B2(new_n617), .ZN(new_n631));
  OAI211_X1 g0431(.A(KEYINPUT21), .B(new_n615), .C1(new_n629), .C2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n608), .A2(new_n508), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n633), .B1(new_n267), .B2(new_n613), .ZN(new_n634));
  OAI211_X1 g0434(.A(G179), .B(new_n634), .C1(new_n629), .C2(new_n631), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n618), .A2(new_n627), .A3(new_n619), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n627), .B1(new_n618), .B2(new_n619), .ZN(new_n638));
  OAI22_X1  g0438(.A1(new_n637), .A2(new_n638), .B1(new_n619), .B2(new_n618), .ZN(new_n639));
  INV_X1    g0439(.A(new_n631), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(KEYINPUT21), .B1(new_n641), .B2(new_n615), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n636), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n503), .A2(new_n215), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n252), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT85), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n646), .B1(new_n507), .B2(new_n503), .ZN(new_n647));
  AND4_X1   g0447(.A1(new_n646), .A2(new_n252), .A3(G274), .A4(new_n503), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(G238), .A2(G1698), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n650), .B1(new_n219), .B2(G1698), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n651), .A2(new_n271), .A3(new_n270), .A4(new_n273), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n617), .A2(G33), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n370), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n649), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n421), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT19), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n227), .B1(new_n431), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(G87), .B2(new_n207), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n227), .A2(G33), .A3(G97), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n660), .A2(KEYINPUT87), .A3(new_n657), .ZN(new_n661));
  AOI21_X1  g0461(.A(KEYINPUT87), .B1(new_n660), .B2(new_n657), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n659), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n274), .A2(G20), .A3(new_n212), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n307), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n409), .A2(new_n323), .ZN(new_n666));
  OAI211_X1 g0466(.A(new_n665), .B(new_n666), .C1(new_n409), .C2(new_n536), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n656), .B(new_n667), .C1(G169), .C2(new_n655), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n537), .A2(G87), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n665), .A2(new_n669), .A3(new_n666), .ZN(new_n670));
  INV_X1    g0470(.A(new_n503), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT85), .B1(new_n515), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n507), .A2(new_n646), .A3(new_n503), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n672), .A2(new_n673), .B1(new_n252), .B2(new_n644), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n219), .A2(G1698), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(G238), .B2(G1698), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n653), .B1(new_n274), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n267), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n400), .B1(new_n674), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(KEYINPUT88), .B1(new_n670), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n551), .A2(new_n227), .A3(G68), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n660), .A2(new_n657), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT87), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n660), .A2(KEYINPUT87), .A3(new_n657), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n681), .A2(new_n686), .A3(new_n659), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n687), .A2(new_n307), .B1(new_n323), .B2(new_n409), .ZN(new_n688));
  OAI21_X1  g0488(.A(G200), .B1(new_n649), .B2(new_n654), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT88), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n688), .A2(new_n689), .A3(new_n690), .A4(new_n669), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n655), .A2(G190), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n680), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n609), .A2(new_n614), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(G200), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n609), .A2(new_n614), .A3(G190), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n695), .A2(new_n639), .A3(new_n640), .A4(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n643), .A2(new_n668), .A3(new_n693), .A4(new_n697), .ZN(new_n698));
  NOR3_X1   g0498(.A1(new_n491), .A2(new_n607), .A3(new_n698), .ZN(G372));
  NAND2_X1  g0499(.A1(new_n391), .A2(new_n394), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n346), .A2(new_n351), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n484), .A2(new_n473), .A3(new_n485), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(KEYINPUT77), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n486), .ZN(new_n704));
  INV_X1    g0504(.A(new_n425), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n701), .B1(new_n706), .B2(new_n475), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n340), .A2(new_n348), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n700), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n385), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n668), .B(KEYINPUT94), .ZN(new_n713));
  INV_X1    g0513(.A(new_n670), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n714), .A2(new_n689), .A3(new_n692), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n668), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n716), .A2(new_n542), .A3(new_n550), .A4(new_n597), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n615), .B1(new_n629), .B2(new_n631), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT21), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AND4_X1   g0520(.A1(new_n606), .A2(new_n720), .A3(new_n635), .A4(new_n632), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n713), .B1(new_n717), .B2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT26), .ZN(new_n723));
  AOI21_X1  g0523(.A(G169), .B1(new_n545), .B2(new_n546), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n525), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n544), .A2(new_n548), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n668), .A2(new_n715), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n723), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n542), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n730), .A2(KEYINPUT26), .A3(new_n668), .A4(new_n693), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n490), .B1(new_n722), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n712), .A2(new_n733), .ZN(G369));
  NAND3_X1  g0534(.A1(new_n253), .A2(new_n227), .A3(G13), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n735), .A2(KEYINPUT27), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(KEYINPUT27), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n736), .A2(G213), .A3(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G343), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n641), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n643), .A2(new_n697), .A3(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n742), .B1(new_n643), .B2(new_n741), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G330), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n597), .A2(new_n606), .ZN(new_n746));
  INV_X1    g0546(.A(new_n740), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n586), .A2(new_n747), .ZN(new_n748));
  OAI22_X1  g0548(.A1(new_n746), .A2(new_n748), .B1(new_n606), .B2(new_n747), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n643), .A2(new_n740), .ZN(new_n751));
  INV_X1    g0551(.A(new_n746), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n601), .A2(new_n605), .A3(new_n747), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT95), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n753), .A2(KEYINPUT95), .A3(new_n754), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n750), .A2(new_n759), .ZN(G399));
  INV_X1    g0560(.A(new_n231), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G41), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n763), .A2(G1), .A3(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n765), .B1(new_n224), .B2(new_n763), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT28), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n747), .B1(new_n732), .B2(new_n722), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT29), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n693), .A2(new_n668), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n723), .B1(new_n771), .B2(new_n542), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n716), .A2(KEYINPUT26), .A3(new_n725), .A4(new_n726), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  OAI211_X1 g0575(.A(KEYINPUT29), .B(new_n747), .C1(new_n775), .C2(new_n722), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n770), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT30), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n545), .A2(new_n546), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n655), .A2(new_n634), .A3(G179), .A4(new_n591), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n591), .A2(new_n678), .A3(new_n674), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n609), .A2(new_n614), .A3(G179), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n784), .A2(KEYINPUT30), .A3(new_n545), .A4(new_n546), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n655), .A2(new_n634), .A3(G179), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n786), .A2(new_n524), .A3(new_n599), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n781), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(new_n740), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT31), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT96), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n720), .A2(new_n635), .A3(new_n632), .A4(new_n697), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n771), .A2(new_n794), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n542), .A2(new_n550), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n795), .A2(new_n796), .A3(new_n752), .A4(new_n747), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n788), .A2(KEYINPUT31), .A3(new_n740), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n792), .B1(new_n791), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(G330), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  AND2_X1   g0601(.A1(new_n777), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n767), .B1(new_n802), .B2(G1), .ZN(G364));
  INV_X1    g0603(.A(G13), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(G20), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n253), .B1(new_n805), .B2(G45), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n762), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(G13), .A2(G33), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(G20), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  OR2_X1    g0613(.A1(new_n743), .A2(new_n813), .ZN(new_n814));
  NOR4_X1   g0614(.A1(new_n227), .A2(new_n421), .A3(new_n341), .A4(G200), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(G322), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n312), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n227), .A2(G179), .ZN(new_n819));
  NOR2_X1   g0619(.A1(G190), .A2(G200), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n818), .B1(G329), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n227), .A2(new_n421), .ZN(new_n824));
  AND3_X1   g0624(.A1(new_n824), .A2(KEYINPUT98), .A3(new_n820), .ZN(new_n825));
  AOI21_X1  g0625(.A(KEYINPUT98), .B1(new_n824), .B2(new_n820), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(G311), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n824), .A2(G200), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n830), .A2(new_n341), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n819), .A2(G190), .A3(G200), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n831), .A2(G326), .B1(new_n833), .B2(G303), .ZN(new_n834));
  NOR3_X1   g0634(.A1(new_n341), .A2(G179), .A3(G200), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(new_n227), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n819), .A2(new_n341), .A3(G200), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n837), .A2(G294), .B1(new_n839), .B2(G283), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n823), .A2(new_n829), .A3(new_n834), .A4(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n824), .A2(new_n341), .A3(G200), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n842), .A2(KEYINPUT100), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n842), .A2(KEYINPUT100), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XOR2_X1   g0645(.A(KEYINPUT33), .B(G317), .Z(new_n846));
  NOR2_X1   g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n828), .A2(G77), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT32), .ZN(new_n849));
  INV_X1    g0649(.A(G159), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n821), .A2(new_n850), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n849), .A2(new_n851), .B1(new_n839), .B2(G107), .ZN(new_n852));
  AOI22_X1  g0652(.A1(G97), .A2(new_n837), .B1(new_n831), .B2(G50), .ZN(new_n853));
  INV_X1    g0653(.A(new_n851), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n854), .A2(KEYINPUT32), .B1(G58), .B2(new_n815), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n848), .A2(new_n852), .A3(new_n853), .A4(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n832), .A2(new_n214), .ZN(new_n857));
  OR3_X1    g0657(.A1(new_n857), .A2(KEYINPUT99), .A3(new_n312), .ZN(new_n858));
  OAI21_X1  g0658(.A(KEYINPUT99), .B1(new_n857), .B2(new_n312), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n858), .B(new_n859), .C1(new_n845), .C2(new_n212), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n841), .A2(new_n847), .B1(new_n856), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n226), .B1(G20), .B2(new_n286), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n812), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n761), .A2(new_n312), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n864), .B(KEYINPUT97), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n865), .A2(G355), .B1(new_n630), .B2(new_n761), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n249), .A2(new_n258), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n551), .A2(new_n761), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(G45), .B2(new_n225), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n866), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n861), .A2(new_n862), .B1(new_n863), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n809), .B1(new_n814), .B2(new_n871), .ZN(new_n872));
  OR2_X1    g0672(.A1(new_n743), .A2(G330), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n808), .B1(new_n873), .B2(new_n744), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n875), .B(KEYINPUT101), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(G396));
  NOR2_X1   g0677(.A1(new_n425), .A2(new_n740), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n424), .A2(new_n740), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n419), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n878), .B1(new_n880), .B2(new_n425), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n768), .B(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n808), .B1(new_n882), .B2(new_n801), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n801), .B2(new_n882), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n881), .A2(new_n811), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n828), .A2(new_n617), .B1(G303), .B2(new_n831), .ZN(new_n886));
  INV_X1    g0686(.A(G283), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n886), .B1(new_n887), .B2(new_n845), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n888), .B(KEYINPUT102), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n312), .B1(new_n832), .B2(new_n206), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n890), .B(KEYINPUT103), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n822), .A2(G311), .B1(new_n815), .B2(G294), .ZN(new_n892));
  OAI221_X1 g0692(.A(new_n892), .B1(new_n214), .B2(new_n838), .C1(new_n205), .C2(new_n836), .ZN(new_n893));
  NOR3_X1   g0693(.A1(new_n889), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  OAI22_X1  g0694(.A1(new_n836), .A2(new_n288), .B1(new_n838), .B2(new_n212), .ZN(new_n895));
  INV_X1    g0695(.A(G132), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n551), .B1(new_n896), .B2(new_n821), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n895), .B(new_n897), .C1(G50), .C2(new_n833), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n831), .A2(G137), .B1(G143), .B2(new_n815), .ZN(new_n899));
  INV_X1    g0699(.A(G150), .ZN(new_n900));
  OAI221_X1 g0700(.A(new_n899), .B1(new_n850), .B2(new_n827), .C1(new_n845), .C2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT34), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n898), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n903), .B1(new_n902), .B2(new_n901), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n862), .B1(new_n894), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n862), .A2(new_n810), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n905), .B1(G77), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n808), .B1(new_n885), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n884), .A2(new_n909), .ZN(new_n910));
  XOR2_X1   g0710(.A(new_n910), .B(KEYINPUT104), .Z(G384));
  NOR2_X1   g0711(.A1(new_n805), .A2(new_n253), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n302), .A2(new_n307), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n274), .A2(new_n297), .ZN(new_n914));
  INV_X1    g0714(.A(new_n298), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n916), .A2(G68), .A3(new_n299), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT16), .B1(new_n917), .B2(new_n294), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n337), .B1(new_n913), .B2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n738), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n352), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n338), .A2(new_n920), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT37), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n339), .A2(new_n344), .A3(new_n924), .A4(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n287), .A2(new_n919), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n927), .A2(new_n921), .A3(new_n344), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n926), .B1(new_n928), .B2(new_n925), .ZN(new_n929));
  AND3_X1   g0729(.A1(new_n923), .A2(new_n929), .A3(KEYINPUT38), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT38), .B1(new_n923), .B2(new_n929), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT39), .ZN(new_n932));
  OR3_X1    g0732(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n923), .A2(new_n929), .A3(KEYINPUT38), .ZN(new_n934));
  INV_X1    g0734(.A(new_n924), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n339), .A2(new_n344), .A3(new_n924), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(KEYINPUT37), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n352), .A2(new_n935), .B1(new_n937), .B2(new_n926), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n934), .B1(KEYINPUT38), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n932), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n933), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n475), .A2(new_n740), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n878), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n880), .A2(new_n425), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n944), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n944), .B1(new_n768), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n473), .A2(new_n747), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n488), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n948), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n704), .A2(new_n475), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n947), .B(new_n952), .C1(new_n930), .C2(new_n931), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n708), .A2(new_n738), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n943), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n770), .A2(new_n490), .A3(new_n776), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(KEYINPUT106), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT106), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n770), .A2(new_n958), .A3(new_n490), .A4(new_n776), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n712), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n955), .B(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(G330), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT107), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n352), .A2(new_n935), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n937), .A2(new_n926), .ZN(new_n966));
  AOI21_X1  g0766(.A(KEYINPUT38), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n930), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n797), .A2(new_n791), .A3(new_n799), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n969), .A2(new_n952), .A3(KEYINPUT40), .A4(new_n881), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n964), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n791), .A2(new_n799), .ZN(new_n972));
  NOR3_X1   g0772(.A1(new_n698), .A2(new_n607), .A3(new_n740), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI221_X4 g0774(.A(new_n948), .B1(new_n459), .B2(new_n474), .C1(new_n703), .C2(new_n486), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n950), .B1(new_n704), .B2(new_n475), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n881), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n978), .A2(KEYINPUT107), .A3(KEYINPUT40), .A4(new_n939), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT40), .ZN(new_n980));
  INV_X1    g0780(.A(new_n977), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n981), .B(new_n969), .C1(new_n930), .C2(new_n931), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n971), .A2(new_n979), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n491), .A2(new_n974), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n963), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n983), .B2(new_n984), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n912), .B1(new_n962), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n962), .B2(new_n986), .ZN(new_n988));
  INV_X1    g0788(.A(new_n531), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n630), .B(new_n229), .C1(new_n989), .C2(KEYINPUT35), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(KEYINPUT35), .B2(new_n989), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT36), .ZN(new_n992));
  NOR3_X1   g0792(.A1(new_n289), .A2(new_n224), .A3(new_n218), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT105), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n993), .A2(new_n994), .B1(new_n202), .B2(G68), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n994), .B2(new_n993), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n996), .A2(G1), .A3(new_n804), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n988), .A2(new_n992), .A3(new_n997), .ZN(G367));
  INV_X1    g0798(.A(new_n868), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n863), .B1(new_n231), .B2(new_n409), .C1(new_n999), .C2(new_n242), .ZN(new_n1000));
  AND2_X1   g0800(.A1(new_n1000), .A2(new_n808), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n670), .A2(new_n740), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n716), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n713), .B2(new_n1002), .ZN(new_n1004));
  INV_X1    g0804(.A(G137), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n309), .B1(new_n821), .B2(new_n1005), .C1(new_n816), .C2(new_n900), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(new_n828), .B2(G50), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n836), .A2(new_n212), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n288), .A2(new_n832), .B1(new_n838), .B2(new_n218), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n1008), .B(new_n1009), .C1(G143), .C2(new_n831), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1007), .B(new_n1010), .C1(new_n850), .C2(new_n845), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT46), .ZN(new_n1012));
  NOR3_X1   g0812(.A1(new_n832), .A2(new_n1012), .A3(new_n630), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(G107), .B2(new_n837), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n831), .A2(G311), .B1(new_n839), .B2(G97), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1014), .B(new_n1015), .C1(new_n589), .C2(new_n845), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n828), .A2(G283), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n617), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1012), .B1(new_n1018), .B2(new_n832), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n822), .A2(G317), .B1(new_n815), .B2(G303), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1017), .A2(new_n274), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1011), .B1(new_n1016), .B2(new_n1021), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT47), .Z(new_n1023));
  INV_X1    g0823(.A(new_n862), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1001), .B1(new_n1004), .B2(new_n813), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n747), .B1(new_n544), .B2(new_n548), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n724), .B2(new_n525), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n796), .B2(new_n1026), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n542), .B1(new_n1028), .B2(new_n606), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT108), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1031), .A2(new_n747), .A3(new_n1032), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1028), .A2(new_n753), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(KEYINPUT42), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT109), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1033), .A2(KEYINPUT109), .A3(new_n1035), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT110), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1034), .A2(KEYINPUT42), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1040), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1041), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n1045), .A2(new_n1046), .B1(KEYINPUT43), .B2(new_n1004), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1046), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1004), .B(KEYINPUT43), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1048), .A2(new_n1044), .A3(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n750), .A2(new_n1028), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1051), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1047), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n762), .B(KEYINPUT41), .Z(new_n1054));
  INV_X1    g0854(.A(new_n759), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1055), .A2(new_n1028), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT45), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n757), .A2(new_n758), .A3(new_n1028), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT44), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1060), .A2(KEYINPUT112), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(KEYINPUT112), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT111), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1055), .A2(KEYINPUT111), .A3(KEYINPUT44), .A4(new_n1028), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1061), .A2(new_n1062), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n750), .B1(new_n1057), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n753), .B1(new_n749), .B2(new_n751), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n744), .B(new_n1069), .Z(new_n1070));
  NAND3_X1  g0870(.A1(new_n1057), .A2(new_n1066), .A3(new_n750), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1068), .A2(new_n802), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1054), .B1(new_n1072), .B2(new_n802), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1053), .B1(new_n1073), .B2(new_n807), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1052), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1025), .B1(new_n1074), .B2(new_n1075), .ZN(G387));
  AOI22_X1  g0876(.A1(new_n831), .A2(G322), .B1(G317), .B2(new_n815), .ZN(new_n1077));
  INV_X1    g0877(.A(G311), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1077), .B1(new_n612), .B2(new_n827), .C1(new_n845), .C2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT48), .ZN(new_n1080));
  OR2_X1    g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n837), .A2(G283), .B1(new_n833), .B2(G294), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT49), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1018), .A2(new_n838), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n551), .B(new_n1088), .C1(G326), .C2(new_n822), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1086), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n836), .A2(new_n409), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n831), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n1092), .A2(new_n850), .B1(new_n832), .B2(new_n218), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n1091), .B(new_n1093), .C1(G97), .C2(new_n839), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n816), .A2(new_n202), .B1(new_n821), .B2(new_n900), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n274), .B(new_n1095), .C1(new_n828), .C2(G68), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1094), .B(new_n1096), .C1(new_n321), .C2(new_n845), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1024), .B1(new_n1090), .B2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n868), .B1(new_n239), .B2(new_n258), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n865), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1099), .B1(new_n764), .B2(new_n1100), .ZN(new_n1101));
  OR3_X1    g0901(.A1(new_n406), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1102));
  OAI21_X1  g0902(.A(KEYINPUT50), .B1(new_n406), .B2(G50), .ZN(new_n1103));
  AOI21_X1  g0903(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1102), .A2(new_n764), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n1101), .A2(new_n1105), .B1(new_n206), .B2(new_n761), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n863), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n808), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1098), .A2(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT113), .ZN(new_n1110));
  OR2_X1    g0910(.A1(new_n749), .A2(new_n813), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n1110), .A2(new_n1111), .B1(new_n807), .B2(new_n1070), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n802), .A2(new_n1070), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n762), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n802), .A2(new_n1070), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1112), .B1(new_n1114), .B2(new_n1115), .ZN(G393));
  INV_X1    g0916(.A(new_n1071), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1113), .B1(new_n1117), .B2(new_n1067), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1072), .A2(new_n1118), .A3(new_n762), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n246), .A2(new_n868), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n863), .B1(new_n205), .B2(new_n231), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n831), .A2(G317), .B1(G311), .B2(new_n815), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT52), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n845), .A2(new_n612), .B1(new_n1018), .B2(new_n836), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT116), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n1123), .B(new_n1126), .C1(G294), .C2(new_n828), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n312), .B1(new_n821), .B2(new_n817), .C1(new_n206), .C2(new_n838), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(G283), .B2(new_n833), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT115), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(new_n1125), .B2(new_n1124), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n836), .A2(new_n218), .B1(new_n838), .B2(new_n214), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n274), .B1(new_n822), .B2(G143), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n827), .B2(new_n406), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n1132), .B(new_n1134), .C1(G68), .C2(new_n833), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n1092), .A2(new_n900), .B1(new_n850), .B2(new_n816), .ZN(new_n1136));
  XOR2_X1   g0936(.A(KEYINPUT114), .B(KEYINPUT51), .Z(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  AND2_X1   g0939(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n845), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n1139), .B(new_n1140), .C1(G50), .C2(new_n1141), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n1127), .A2(new_n1131), .B1(new_n1135), .B2(new_n1142), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n808), .B1(new_n1120), .B2(new_n1121), .C1(new_n1143), .C2(new_n1024), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(new_n812), .B2(new_n1028), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1117), .A2(new_n1067), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1145), .B1(new_n1146), .B2(new_n807), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1119), .A2(new_n1147), .ZN(G390));
  OAI21_X1  g0948(.A(new_n309), .B1(new_n816), .B2(new_n896), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(G125), .B2(new_n822), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n832), .A2(new_n900), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT53), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(KEYINPUT54), .B(G143), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1150), .B(new_n1152), .C1(new_n827), .C2(new_n1153), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n831), .A2(G128), .B1(new_n839), .B2(G50), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n1155), .B1(new_n850), .B2(new_n836), .C1(new_n845), .C2(new_n1005), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n845), .A2(new_n206), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n828), .A2(G97), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n857), .B1(G68), .B2(new_n839), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(G77), .A2(new_n837), .B1(new_n831), .B2(G283), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n312), .B1(new_n821), .B2(new_n589), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(G116), .B2(new_n815), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .A4(new_n1162), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n1154), .A2(new_n1156), .B1(new_n1157), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n862), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n809), .B1(new_n321), .B2(new_n906), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1165), .B(new_n1166), .C1(new_n941), .C2(new_n811), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n974), .A2(new_n963), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1168), .A2(KEYINPUT118), .A3(new_n981), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT118), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n969), .A2(G330), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1170), .B1(new_n1171), .B2(new_n977), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1173));
  XOR2_X1   g0973(.A(new_n942), .B(KEYINPUT117), .Z(new_n1174));
  NOR2_X1   g0974(.A1(new_n968), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n713), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n717), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n721), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1176), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n740), .B1(new_n1179), .B2(new_n774), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n878), .B1(new_n1180), .B2(new_n945), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n952), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1175), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n947), .A2(new_n952), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n942), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n1185), .A2(new_n1186), .B1(new_n933), .B2(new_n940), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1173), .B1(new_n1184), .B2(new_n1187), .ZN(new_n1188));
  OAI211_X1 g0988(.A(G330), .B(new_n881), .C1(new_n798), .C2(new_n800), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1189), .A2(new_n1182), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n942), .B1(new_n947), .B2(new_n952), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1183), .B(new_n1190), .C1(new_n941), .C2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1188), .A2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1167), .B1(new_n1193), .B2(new_n806), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1189), .A2(new_n1182), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1169), .A2(new_n1195), .A3(new_n1172), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(new_n947), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1182), .B1(new_n1171), .B2(new_n946), .ZN(new_n1198));
  AND2_X1   g0998(.A1(new_n1198), .A2(new_n1181), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(new_n1190), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n491), .A2(new_n1171), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n711), .B(new_n1202), .C1(new_n957), .C2(new_n959), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1201), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n763), .B1(new_n1193), .B2(new_n1204), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1188), .A2(new_n1201), .A3(new_n1203), .A4(new_n1192), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1194), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(G378));
  NAND2_X1  g1008(.A1(new_n971), .A2(new_n979), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n963), .B1(new_n982), .B2(new_n980), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT121), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1209), .A2(new_n1210), .A3(KEYINPUT121), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n387), .A2(new_n920), .ZN(new_n1215));
  XOR2_X1   g1015(.A(new_n1215), .B(KEYINPUT55), .Z(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  AND2_X1   g1017(.A1(new_n395), .A2(new_n1217), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n395), .A2(new_n1217), .ZN(new_n1219));
  XOR2_X1   g1019(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  OR3_X1    g1021(.A1(new_n1218), .A2(new_n1219), .A3(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1221), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1213), .A2(new_n1214), .A3(new_n1225), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1209), .A2(new_n1210), .A3(KEYINPUT121), .A4(new_n1224), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n955), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n955), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1226), .A2(new_n1227), .A3(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1229), .A2(new_n807), .A3(new_n1231), .ZN(new_n1232));
  OR2_X1    g1032(.A1(new_n827), .A2(new_n409), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1008), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n551), .A2(G41), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n822), .A2(G283), .B1(new_n815), .B2(G107), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .A4(new_n1236), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n845), .A2(new_n205), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n838), .A2(new_n288), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n1092), .A2(new_n630), .B1(new_n832), .B2(new_n218), .ZN(new_n1240));
  NOR4_X1   g1040(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .A4(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(KEYINPUT58), .ZN(new_n1242));
  AOI211_X1 g1042(.A(G50), .B(new_n1235), .C1(new_n269), .C2(new_n257), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n1243), .B(KEYINPUT119), .ZN(new_n1244));
  AND2_X1   g1044(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n836), .A2(new_n900), .B1(new_n832), .B2(new_n1153), .ZN(new_n1246));
  INV_X1    g1046(.A(G128), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n816), .A2(new_n1247), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1246), .B(new_n1248), .C1(G125), .C2(new_n831), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n1249), .B1(new_n896), .B2(new_n845), .C1(new_n1005), .C2(new_n827), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(KEYINPUT59), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n839), .A2(G159), .ZN(new_n1252));
  AOI211_X1 g1052(.A(G33), .B(G41), .C1(new_n822), .C2(G124), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1251), .A2(new_n1252), .A3(new_n1253), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1250), .A2(KEYINPUT59), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n1245), .B1(KEYINPUT58), .B2(new_n1241), .C1(new_n1254), .C2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n862), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n809), .B1(new_n202), .B2(new_n906), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1257), .B(new_n1258), .C1(new_n1225), .C2(new_n811), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1232), .A2(new_n1259), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1226), .A2(new_n1230), .A3(new_n1227), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1230), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT57), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(new_n1206), .B2(new_n1203), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n763), .B1(new_n1263), .B2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1206), .A2(new_n1203), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1229), .A2(new_n1231), .A3(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1264), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1260), .B1(new_n1266), .B2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1271), .A2(KEYINPUT122), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT122), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1270), .A2(new_n1273), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1272), .A2(new_n1274), .ZN(G375));
  NAND2_X1  g1075(.A1(new_n1201), .A2(new_n807), .ZN(new_n1276));
  OAI22_X1  g1076(.A1(new_n1092), .A2(new_n896), .B1(new_n1005), .B2(new_n816), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1153), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1277), .B1(new_n1141), .B2(new_n1278), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1279), .A2(KEYINPUT124), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1279), .A2(KEYINPUT124), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1239), .B1(G50), .B2(new_n837), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1282), .B1(new_n850), .B2(new_n832), .ZN(new_n1283));
  OAI221_X1 g1083(.A(new_n551), .B1(new_n1247), .B2(new_n821), .C1(new_n827), .C2(new_n900), .ZN(new_n1284));
  NOR4_X1   g1084(.A1(new_n1280), .A2(new_n1281), .A3(new_n1283), .A4(new_n1284), .ZN(new_n1285));
  OAI221_X1 g1085(.A(new_n312), .B1(new_n821), .B2(new_n612), .C1(new_n816), .C2(new_n887), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1286), .B1(new_n828), .B2(G107), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1091), .B1(G77), .B2(new_n839), .ZN(new_n1288));
  AOI22_X1  g1088(.A1(new_n831), .A2(G294), .B1(new_n833), .B2(G97), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1287), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1290), .B1(new_n617), .B2(new_n1141), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n862), .B1(new_n1285), .B2(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n809), .B1(new_n212), .B2(new_n906), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1292), .B(new_n1293), .C1(new_n952), .C2(new_n811), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1276), .A2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(KEYINPUT125), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT125), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1276), .A2(new_n1297), .A3(new_n1294), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1296), .A2(new_n1298), .ZN(new_n1299));
  AOI22_X1  g1099(.A1(new_n947), .A2(new_n1196), .B1(new_n1199), .B2(new_n1190), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1202), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n960), .A2(new_n712), .A3(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1300), .A2(new_n1302), .ZN(new_n1303));
  XOR2_X1   g1103(.A(new_n1054), .B(KEYINPUT123), .Z(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1204), .A2(new_n1303), .A3(new_n1305), .ZN(new_n1306));
  AND2_X1   g1106(.A1(new_n1299), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(G381));
  NOR4_X1   g1108(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1309), .A2(new_n1207), .A3(new_n1307), .ZN(new_n1310));
  OR3_X1    g1110(.A1(G375), .A2(G387), .A3(new_n1310), .ZN(G407));
  OAI21_X1  g1111(.A(new_n1207), .B1(new_n1272), .B2(new_n1274), .ZN(new_n1312));
  OAI211_X1 g1112(.A(G407), .B(G213), .C1(G343), .C2(new_n1312), .ZN(G409));
  INV_X1    g1113(.A(new_n1259), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1314), .B1(new_n1263), .B2(new_n807), .ZN(new_n1315));
  AOI21_X1  g1115(.A(KEYINPUT57), .B1(new_n1263), .B2(new_n1267), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1265), .A2(new_n1229), .A3(new_n1231), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(new_n762), .ZN(new_n1318));
  OAI211_X1 g1118(.A(G378), .B(new_n1315), .C1(new_n1316), .C2(new_n1318), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1268), .A2(new_n1304), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1207), .B1(new_n1320), .B2(new_n1260), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1319), .A2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(G384), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1300), .A2(new_n1302), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT60), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1303), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1300), .A2(new_n1302), .A3(KEYINPUT60), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1326), .A2(KEYINPUT126), .A3(new_n762), .A4(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1328), .A2(new_n1299), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1204), .A2(KEYINPUT60), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n763), .B1(new_n1330), .B2(new_n1303), .ZN(new_n1331));
  AOI21_X1  g1131(.A(KEYINPUT126), .B1(new_n1331), .B2(new_n1327), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1323), .B1(new_n1329), .B2(new_n1332), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1326), .A2(new_n762), .A3(new_n1327), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT126), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  NAND4_X1  g1136(.A1(new_n1336), .A2(G384), .A3(new_n1299), .A4(new_n1328), .ZN(new_n1337));
  AND2_X1   g1137(.A1(new_n1333), .A2(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(G213), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1339), .A2(G343), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1340), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1322), .A2(new_n1338), .A3(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(KEYINPUT62), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1333), .A2(new_n1337), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1344), .A2(G2897), .A3(new_n1340), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1340), .A2(G2897), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1333), .A2(new_n1337), .A3(new_n1346), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1263), .A2(new_n1267), .A3(new_n1305), .ZN(new_n1348));
  AOI21_X1  g1148(.A(G378), .B1(new_n1315), .B2(new_n1348), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1349), .B1(G378), .B2(new_n1270), .ZN(new_n1350));
  OAI211_X1 g1150(.A(new_n1345), .B(new_n1347), .C1(new_n1350), .C2(new_n1340), .ZN(new_n1351));
  XNOR2_X1  g1151(.A(KEYINPUT127), .B(KEYINPUT61), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT62), .ZN(new_n1353));
  NAND4_X1  g1153(.A1(new_n1322), .A2(new_n1338), .A3(new_n1353), .A4(new_n1341), .ZN(new_n1354));
  NAND4_X1  g1154(.A1(new_n1343), .A2(new_n1351), .A3(new_n1352), .A4(new_n1354), .ZN(new_n1355));
  XNOR2_X1  g1155(.A(G393), .B(new_n876), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(G390), .A2(new_n1356), .ZN(new_n1357));
  INV_X1    g1157(.A(new_n1356), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1358), .A2(new_n1119), .A3(new_n1147), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1357), .A2(new_n1359), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(G387), .A2(new_n1360), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1075), .ZN(new_n1362));
  OAI211_X1 g1162(.A(new_n1362), .B(new_n1053), .C1(new_n807), .C2(new_n1073), .ZN(new_n1363));
  NAND4_X1  g1163(.A1(new_n1363), .A2(new_n1025), .A3(new_n1357), .A4(new_n1359), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1361), .A2(new_n1364), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1355), .A2(new_n1365), .ZN(new_n1366));
  NOR2_X1   g1166(.A1(new_n1365), .A2(KEYINPUT61), .ZN(new_n1367));
  INV_X1    g1167(.A(KEYINPUT63), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1342), .A2(new_n1368), .ZN(new_n1369));
  NAND4_X1  g1169(.A1(new_n1322), .A2(new_n1338), .A3(KEYINPUT63), .A4(new_n1341), .ZN(new_n1370));
  NAND4_X1  g1170(.A1(new_n1367), .A2(new_n1369), .A3(new_n1351), .A4(new_n1370), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1366), .A2(new_n1371), .ZN(G405));
  NAND2_X1  g1172(.A1(new_n1271), .A2(G378), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1312), .A2(new_n1373), .ZN(new_n1374));
  NOR2_X1   g1174(.A1(G387), .A2(new_n1360), .ZN(new_n1375));
  AOI22_X1  g1175(.A1(new_n1363), .A2(new_n1025), .B1(new_n1357), .B2(new_n1359), .ZN(new_n1376));
  OAI21_X1  g1176(.A(new_n1344), .B1(new_n1375), .B2(new_n1376), .ZN(new_n1377));
  NAND3_X1  g1177(.A1(new_n1361), .A2(new_n1364), .A3(new_n1338), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1377), .A2(new_n1378), .ZN(new_n1379));
  XNOR2_X1  g1179(.A(new_n1374), .B(new_n1379), .ZN(G402));
endmodule


