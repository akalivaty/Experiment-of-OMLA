

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580;

  XNOR2_X1 U323 ( .A(n450), .B(KEYINPUT38), .ZN(n495) );
  XOR2_X1 U324 ( .A(n471), .B(KEYINPUT28), .Z(n518) );
  XOR2_X1 U325 ( .A(n440), .B(n439), .Z(n291) );
  XOR2_X1 U326 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n292) );
  NOR2_X1 U327 ( .A1(n465), .A2(n464), .ZN(n466) );
  XNOR2_X1 U328 ( .A(n441), .B(n291), .ZN(n442) );
  INV_X1 U329 ( .A(G169GAT), .ZN(n305) );
  XNOR2_X1 U330 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U331 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U332 ( .A(n308), .B(n307), .ZN(n360) );
  XOR2_X1 U333 ( .A(KEYINPUT79), .B(n547), .Z(n559) );
  INV_X1 U334 ( .A(G43GAT), .ZN(n451) );
  XNOR2_X1 U335 ( .A(G183GAT), .B(KEYINPUT122), .ZN(n474) );
  XNOR2_X1 U336 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U337 ( .A(n475), .B(n474), .ZN(G1350GAT) );
  XNOR2_X1 U338 ( .A(n454), .B(n453), .ZN(G1330GAT) );
  XOR2_X1 U339 ( .A(KEYINPUT83), .B(KEYINPUT87), .Z(n298) );
  XNOR2_X1 U340 ( .A(G134GAT), .B(G43GAT), .ZN(n293) );
  XNOR2_X1 U341 ( .A(n293), .B(G190GAT), .ZN(n430) );
  XOR2_X1 U342 ( .A(KEYINPUT20), .B(KEYINPUT86), .Z(n295) );
  XNOR2_X1 U343 ( .A(G99GAT), .B(KEYINPUT85), .ZN(n294) );
  XNOR2_X1 U344 ( .A(n295), .B(n294), .ZN(n296) );
  XNOR2_X1 U345 ( .A(n430), .B(n296), .ZN(n297) );
  XNOR2_X1 U346 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U347 ( .A(G127GAT), .B(G15GAT), .Z(n422) );
  XOR2_X1 U348 ( .A(G120GAT), .B(G71GAT), .Z(n333) );
  XOR2_X1 U349 ( .A(n422), .B(n333), .Z(n300) );
  NAND2_X1 U350 ( .A1(G227GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U351 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U352 ( .A(n302), .B(n301), .Z(n310) );
  XOR2_X1 U353 ( .A(KEYINPUT0), .B(G113GAT), .Z(n388) );
  XOR2_X1 U354 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n304) );
  XNOR2_X1 U355 ( .A(KEYINPUT18), .B(KEYINPUT84), .ZN(n303) );
  XNOR2_X1 U356 ( .A(n304), .B(n303), .ZN(n308) );
  XNOR2_X1 U357 ( .A(G183GAT), .B(G176GAT), .ZN(n306) );
  XNOR2_X1 U358 ( .A(n388), .B(n360), .ZN(n309) );
  XNOR2_X2 U359 ( .A(n310), .B(n309), .ZN(n524) );
  XNOR2_X1 U360 ( .A(G29GAT), .B(KEYINPUT70), .ZN(n311) );
  XNOR2_X1 U361 ( .A(n292), .B(n311), .ZN(n434) );
  XOR2_X1 U362 ( .A(n434), .B(KEYINPUT69), .Z(n313) );
  NAND2_X1 U363 ( .A1(G229GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U364 ( .A(n313), .B(n312), .ZN(n328) );
  XOR2_X1 U365 ( .A(G197GAT), .B(G8GAT), .Z(n315) );
  XNOR2_X1 U366 ( .A(G141GAT), .B(G22GAT), .ZN(n314) );
  XNOR2_X1 U367 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U368 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n317) );
  XNOR2_X1 U369 ( .A(KEYINPUT68), .B(KEYINPUT30), .ZN(n316) );
  XNOR2_X1 U370 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U371 ( .A(n319), .B(n318), .ZN(n326) );
  XOR2_X1 U372 ( .A(G15GAT), .B(G50GAT), .Z(n321) );
  XNOR2_X1 U373 ( .A(G36GAT), .B(G43GAT), .ZN(n320) );
  XNOR2_X1 U374 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U375 ( .A(n322), .B(G169GAT), .Z(n324) );
  XOR2_X1 U376 ( .A(G1GAT), .B(KEYINPUT71), .Z(n419) );
  XNOR2_X1 U377 ( .A(G113GAT), .B(n419), .ZN(n323) );
  XNOR2_X1 U378 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U379 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U380 ( .A(n328), .B(n327), .ZN(n497) );
  XOR2_X1 U381 ( .A(G92GAT), .B(G99GAT), .Z(n330) );
  XNOR2_X1 U382 ( .A(G85GAT), .B(G106GAT), .ZN(n329) );
  XNOR2_X1 U383 ( .A(n330), .B(n329), .ZN(n437) );
  XOR2_X1 U384 ( .A(n437), .B(KEYINPUT72), .Z(n332) );
  NAND2_X1 U385 ( .A1(G230GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U386 ( .A(n332), .B(n331), .ZN(n334) );
  XOR2_X1 U387 ( .A(n334), .B(n333), .Z(n337) );
  XNOR2_X1 U388 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n335) );
  XNOR2_X1 U389 ( .A(n335), .B(G64GAT), .ZN(n414) );
  XOR2_X1 U390 ( .A(G148GAT), .B(G78GAT), .Z(n367) );
  XNOR2_X1 U391 ( .A(n414), .B(n367), .ZN(n336) );
  XNOR2_X1 U392 ( .A(n337), .B(n336), .ZN(n345) );
  XOR2_X1 U393 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n339) );
  XNOR2_X1 U394 ( .A(G176GAT), .B(G204GAT), .ZN(n338) );
  XNOR2_X1 U395 ( .A(n339), .B(n338), .ZN(n343) );
  XOR2_X1 U396 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n341) );
  XNOR2_X1 U397 ( .A(KEYINPUT75), .B(KEYINPUT31), .ZN(n340) );
  XNOR2_X1 U398 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U399 ( .A(n343), .B(n342), .Z(n344) );
  XNOR2_X1 U400 ( .A(n345), .B(n344), .ZN(n570) );
  NOR2_X1 U401 ( .A1(n497), .A2(n570), .ZN(n481) );
  XOR2_X1 U402 ( .A(KEYINPUT105), .B(KEYINPUT37), .Z(n449) );
  XOR2_X1 U403 ( .A(KEYINPUT80), .B(G8GAT), .Z(n420) );
  XOR2_X1 U404 ( .A(n420), .B(G190GAT), .Z(n348) );
  XNOR2_X1 U405 ( .A(G218GAT), .B(G36GAT), .ZN(n346) );
  XNOR2_X1 U406 ( .A(n346), .B(KEYINPUT78), .ZN(n438) );
  XNOR2_X1 U407 ( .A(n438), .B(G92GAT), .ZN(n347) );
  XNOR2_X1 U408 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U409 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n350) );
  NAND2_X1 U410 ( .A1(G226GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U411 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U412 ( .A(n352), .B(n351), .Z(n358) );
  XNOR2_X1 U413 ( .A(G204GAT), .B(KEYINPUT91), .ZN(n353) );
  XNOR2_X1 U414 ( .A(n353), .B(G197GAT), .ZN(n354) );
  XOR2_X1 U415 ( .A(n354), .B(KEYINPUT21), .Z(n356) );
  XNOR2_X1 U416 ( .A(G211GAT), .B(KEYINPUT90), .ZN(n355) );
  XNOR2_X1 U417 ( .A(n356), .B(n355), .ZN(n372) );
  XNOR2_X1 U418 ( .A(G64GAT), .B(n372), .ZN(n357) );
  XNOR2_X1 U419 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U420 ( .A(n360), .B(n359), .ZN(n514) );
  XNOR2_X1 U421 ( .A(KEYINPUT27), .B(n514), .ZN(n404) );
  XOR2_X1 U422 ( .A(KEYINPUT94), .B(KEYINPUT26), .Z(n376) );
  XOR2_X1 U423 ( .A(KEYINPUT23), .B(KEYINPUT89), .Z(n366) );
  XNOR2_X1 U424 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n361) );
  XNOR2_X1 U425 ( .A(n361), .B(KEYINPUT2), .ZN(n392) );
  XOR2_X1 U426 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n363) );
  XNOR2_X1 U427 ( .A(G218GAT), .B(G106GAT), .ZN(n362) );
  XNOR2_X1 U428 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n392), .B(n364), .ZN(n365) );
  XNOR2_X1 U430 ( .A(n366), .B(n365), .ZN(n371) );
  XOR2_X1 U431 ( .A(G155GAT), .B(G22GAT), .Z(n421) );
  XOR2_X1 U432 ( .A(n421), .B(n367), .Z(n369) );
  NAND2_X1 U433 ( .A1(G228GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U434 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U435 ( .A(n371), .B(n370), .Z(n374) );
  XOR2_X1 U436 ( .A(G162GAT), .B(G50GAT), .Z(n431) );
  XNOR2_X1 U437 ( .A(n431), .B(n372), .ZN(n373) );
  XNOR2_X1 U438 ( .A(n374), .B(n373), .ZN(n471) );
  NAND2_X1 U439 ( .A1(n524), .A2(n471), .ZN(n375) );
  XOR2_X1 U440 ( .A(n376), .B(n375), .Z(n565) );
  NOR2_X1 U441 ( .A1(n404), .A2(n565), .ZN(n377) );
  XOR2_X1 U442 ( .A(KEYINPUT95), .B(n377), .Z(n383) );
  OR2_X1 U443 ( .A1(n524), .A2(n514), .ZN(n379) );
  INV_X1 U444 ( .A(n471), .ZN(n378) );
  NAND2_X1 U445 ( .A1(n379), .A2(n378), .ZN(n380) );
  XNOR2_X1 U446 ( .A(n380), .B(KEYINPUT25), .ZN(n381) );
  XNOR2_X1 U447 ( .A(KEYINPUT96), .B(n381), .ZN(n382) );
  NOR2_X1 U448 ( .A1(n383), .A2(n382), .ZN(n384) );
  XNOR2_X1 U449 ( .A(n384), .B(KEYINPUT97), .ZN(n403) );
  XOR2_X1 U450 ( .A(G162GAT), .B(G134GAT), .Z(n386) );
  XNOR2_X1 U451 ( .A(G29GAT), .B(G85GAT), .ZN(n385) );
  XNOR2_X1 U452 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U453 ( .A(n388), .B(n387), .Z(n390) );
  NAND2_X1 U454 ( .A1(G225GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U455 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U456 ( .A(n391), .B(KEYINPUT6), .Z(n394) );
  XNOR2_X1 U457 ( .A(n392), .B(KEYINPUT4), .ZN(n393) );
  XNOR2_X1 U458 ( .A(n394), .B(n393), .ZN(n402) );
  XOR2_X1 U459 ( .A(G148GAT), .B(G155GAT), .Z(n396) );
  XNOR2_X1 U460 ( .A(G127GAT), .B(G120GAT), .ZN(n395) );
  XNOR2_X1 U461 ( .A(n396), .B(n395), .ZN(n400) );
  XOR2_X1 U462 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n398) );
  XNOR2_X1 U463 ( .A(G1GAT), .B(G57GAT), .ZN(n397) );
  XNOR2_X1 U464 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U465 ( .A(n400), .B(n399), .Z(n401) );
  XNOR2_X1 U466 ( .A(n402), .B(n401), .ZN(n512) );
  NAND2_X1 U467 ( .A1(n403), .A2(n512), .ZN(n408) );
  NOR2_X1 U468 ( .A1(n404), .A2(n512), .ZN(n523) );
  INV_X1 U469 ( .A(n518), .ZN(n527) );
  XOR2_X1 U470 ( .A(n524), .B(KEYINPUT88), .Z(n405) );
  NOR2_X1 U471 ( .A1(n527), .A2(n405), .ZN(n406) );
  NAND2_X1 U472 ( .A1(n523), .A2(n406), .ZN(n407) );
  NAND2_X1 U473 ( .A1(n408), .A2(n407), .ZN(n409) );
  XNOR2_X1 U474 ( .A(n409), .B(KEYINPUT98), .ZN(n478) );
  XOR2_X1 U475 ( .A(G78GAT), .B(G211GAT), .Z(n411) );
  XNOR2_X1 U476 ( .A(G71GAT), .B(G183GAT), .ZN(n410) );
  XNOR2_X1 U477 ( .A(n411), .B(n410), .ZN(n428) );
  XOR2_X1 U478 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n413) );
  XNOR2_X1 U479 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n412) );
  XNOR2_X1 U480 ( .A(n413), .B(n412), .ZN(n418) );
  XOR2_X1 U481 ( .A(KEYINPUT12), .B(n414), .Z(n416) );
  NAND2_X1 U482 ( .A1(G231GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U483 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U484 ( .A(n418), .B(n417), .ZN(n426) );
  XOR2_X1 U485 ( .A(n420), .B(n419), .Z(n424) );
  XNOR2_X1 U486 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U487 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U488 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U489 ( .A(n428), .B(n427), .ZN(n476) );
  NAND2_X1 U490 ( .A1(n478), .A2(n476), .ZN(n429) );
  XOR2_X1 U491 ( .A(KEYINPUT104), .B(n429), .Z(n447) );
  XOR2_X1 U492 ( .A(KEYINPUT36), .B(KEYINPUT103), .Z(n446) );
  XOR2_X1 U493 ( .A(n431), .B(n430), .Z(n433) );
  XNOR2_X1 U494 ( .A(KEYINPUT77), .B(KEYINPUT65), .ZN(n432) );
  XNOR2_X1 U495 ( .A(n433), .B(n432), .ZN(n445) );
  XOR2_X1 U496 ( .A(KEYINPUT9), .B(n434), .Z(n436) );
  NAND2_X1 U497 ( .A1(G232GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U498 ( .A(n436), .B(n435), .ZN(n443) );
  XNOR2_X1 U499 ( .A(n438), .B(n437), .ZN(n441) );
  XOR2_X1 U500 ( .A(KEYINPUT11), .B(KEYINPUT76), .Z(n440) );
  XNOR2_X1 U501 ( .A(KEYINPUT66), .B(KEYINPUT10), .ZN(n439) );
  XOR2_X1 U502 ( .A(n445), .B(n444), .Z(n547) );
  XNOR2_X1 U503 ( .A(n446), .B(n559), .ZN(n578) );
  NAND2_X1 U504 ( .A1(n447), .A2(n578), .ZN(n448) );
  XNOR2_X1 U505 ( .A(n449), .B(n448), .ZN(n510) );
  NAND2_X1 U506 ( .A1(n481), .A2(n510), .ZN(n450) );
  NOR2_X1 U507 ( .A1(n524), .A2(n495), .ZN(n454) );
  XNOR2_X1 U508 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n452) );
  INV_X1 U509 ( .A(n514), .ZN(n467) );
  XNOR2_X1 U510 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n455) );
  XNOR2_X1 U511 ( .A(n455), .B(n570), .ZN(n530) );
  NOR2_X1 U512 ( .A1(n497), .A2(n530), .ZN(n456) );
  XNOR2_X1 U513 ( .A(n456), .B(KEYINPUT46), .ZN(n457) );
  NOR2_X1 U514 ( .A1(n547), .A2(n457), .ZN(n458) );
  NAND2_X1 U515 ( .A1(n476), .A2(n458), .ZN(n459) );
  XNOR2_X1 U516 ( .A(n459), .B(KEYINPUT47), .ZN(n460) );
  XNOR2_X1 U517 ( .A(n460), .B(KEYINPUT112), .ZN(n465) );
  INV_X1 U518 ( .A(n476), .ZN(n574) );
  NAND2_X1 U519 ( .A1(n574), .A2(n578), .ZN(n461) );
  XOR2_X1 U520 ( .A(KEYINPUT45), .B(n461), .Z(n462) );
  NAND2_X1 U521 ( .A1(n462), .A2(n497), .ZN(n463) );
  NOR2_X1 U522 ( .A1(n570), .A2(n463), .ZN(n464) );
  XOR2_X1 U523 ( .A(n466), .B(KEYINPUT48), .Z(n522) );
  NAND2_X1 U524 ( .A1(n467), .A2(n522), .ZN(n469) );
  XNOR2_X1 U525 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n468) );
  XNOR2_X1 U526 ( .A(n469), .B(n468), .ZN(n470) );
  NAND2_X1 U527 ( .A1(n470), .A2(n512), .ZN(n564) );
  NOR2_X1 U528 ( .A1(n471), .A2(n564), .ZN(n472) );
  XNOR2_X1 U529 ( .A(n472), .B(KEYINPUT55), .ZN(n473) );
  NOR2_X1 U530 ( .A1(n524), .A2(n473), .ZN(n551) );
  NAND2_X1 U531 ( .A1(n551), .A2(n574), .ZN(n475) );
  XNOR2_X1 U532 ( .A(KEYINPUT102), .B(KEYINPUT34), .ZN(n486) );
  OR2_X1 U533 ( .A1(n476), .A2(n559), .ZN(n477) );
  XOR2_X1 U534 ( .A(KEYINPUT16), .B(n477), .Z(n479) );
  NAND2_X1 U535 ( .A1(n479), .A2(n478), .ZN(n480) );
  XNOR2_X1 U536 ( .A(n480), .B(KEYINPUT99), .ZN(n498) );
  NAND2_X1 U537 ( .A1(n498), .A2(n481), .ZN(n482) );
  XNOR2_X1 U538 ( .A(n482), .B(KEYINPUT100), .ZN(n490) );
  NOR2_X1 U539 ( .A1(n490), .A2(n512), .ZN(n484) );
  XNOR2_X1 U540 ( .A(G1GAT), .B(KEYINPUT101), .ZN(n483) );
  XNOR2_X1 U541 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U542 ( .A(n486), .B(n485), .ZN(G1324GAT) );
  NOR2_X1 U543 ( .A1(n490), .A2(n514), .ZN(n487) );
  XOR2_X1 U544 ( .A(G8GAT), .B(n487), .Z(G1325GAT) );
  XNOR2_X1 U545 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n489) );
  NOR2_X1 U546 ( .A1(n524), .A2(n490), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n489), .B(n488), .ZN(G1326GAT) );
  NOR2_X1 U548 ( .A1(n518), .A2(n490), .ZN(n491) );
  XOR2_X1 U549 ( .A(G22GAT), .B(n491), .Z(G1327GAT) );
  NOR2_X1 U550 ( .A1(n495), .A2(n512), .ZN(n492) );
  XNOR2_X1 U551 ( .A(G29GAT), .B(n492), .ZN(n493) );
  XNOR2_X1 U552 ( .A(n493), .B(KEYINPUT39), .ZN(G1328GAT) );
  NOR2_X1 U553 ( .A1(n495), .A2(n514), .ZN(n494) );
  XOR2_X1 U554 ( .A(G36GAT), .B(n494), .Z(G1329GAT) );
  NOR2_X1 U555 ( .A1(n518), .A2(n495), .ZN(n496) );
  XOR2_X1 U556 ( .A(G50GAT), .B(n496), .Z(G1331GAT) );
  INV_X1 U557 ( .A(n497), .ZN(n566) );
  NOR2_X1 U558 ( .A1(n566), .A2(n530), .ZN(n509) );
  NAND2_X1 U559 ( .A1(n498), .A2(n509), .ZN(n499) );
  XOR2_X1 U560 ( .A(KEYINPUT107), .B(n499), .Z(n505) );
  NOR2_X1 U561 ( .A1(n512), .A2(n505), .ZN(n500) );
  XOR2_X1 U562 ( .A(G57GAT), .B(n500), .Z(n501) );
  XNOR2_X1 U563 ( .A(KEYINPUT42), .B(n501), .ZN(G1332GAT) );
  NOR2_X1 U564 ( .A1(n514), .A2(n505), .ZN(n502) );
  XOR2_X1 U565 ( .A(G64GAT), .B(n502), .Z(G1333GAT) );
  NOR2_X1 U566 ( .A1(n524), .A2(n505), .ZN(n503) );
  XOR2_X1 U567 ( .A(KEYINPUT108), .B(n503), .Z(n504) );
  XNOR2_X1 U568 ( .A(G71GAT), .B(n504), .ZN(G1334GAT) );
  NOR2_X1 U569 ( .A1(n518), .A2(n505), .ZN(n507) );
  XNOR2_X1 U570 ( .A(KEYINPUT109), .B(KEYINPUT43), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U572 ( .A(G78GAT), .B(n508), .Z(G1335GAT) );
  NAND2_X1 U573 ( .A1(n510), .A2(n509), .ZN(n511) );
  XNOR2_X1 U574 ( .A(KEYINPUT110), .B(n511), .ZN(n517) );
  NOR2_X1 U575 ( .A1(n517), .A2(n512), .ZN(n513) );
  XOR2_X1 U576 ( .A(G85GAT), .B(n513), .Z(G1336GAT) );
  NOR2_X1 U577 ( .A1(n517), .A2(n514), .ZN(n515) );
  XOR2_X1 U578 ( .A(G92GAT), .B(n515), .Z(G1337GAT) );
  NOR2_X1 U579 ( .A1(n524), .A2(n517), .ZN(n516) );
  XOR2_X1 U580 ( .A(G99GAT), .B(n516), .Z(G1338GAT) );
  XNOR2_X1 U581 ( .A(KEYINPUT111), .B(KEYINPUT44), .ZN(n520) );
  NOR2_X1 U582 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U583 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U584 ( .A(G106GAT), .B(n521), .ZN(G1339GAT) );
  XNOR2_X1 U585 ( .A(G113GAT), .B(KEYINPUT114), .ZN(n529) );
  NAND2_X1 U586 ( .A1(n523), .A2(n522), .ZN(n539) );
  NOR2_X1 U587 ( .A1(n524), .A2(n539), .ZN(n525) );
  XNOR2_X1 U588 ( .A(n525), .B(KEYINPUT113), .ZN(n526) );
  NOR2_X1 U589 ( .A1(n527), .A2(n526), .ZN(n536) );
  NAND2_X1 U590 ( .A1(n566), .A2(n536), .ZN(n528) );
  XNOR2_X1 U591 ( .A(n529), .B(n528), .ZN(G1340GAT) );
  XOR2_X1 U592 ( .A(G120GAT), .B(KEYINPUT49), .Z(n532) );
  INV_X1 U593 ( .A(n530), .ZN(n556) );
  NAND2_X1 U594 ( .A1(n536), .A2(n556), .ZN(n531) );
  XNOR2_X1 U595 ( .A(n532), .B(n531), .ZN(G1341GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n534) );
  NAND2_X1 U597 ( .A1(n536), .A2(n574), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U599 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U600 ( .A(G134GAT), .B(KEYINPUT51), .Z(n538) );
  NAND2_X1 U601 ( .A1(n536), .A2(n559), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n538), .B(n537), .ZN(G1343GAT) );
  NOR2_X1 U603 ( .A1(n539), .A2(n565), .ZN(n540) );
  XNOR2_X1 U604 ( .A(n540), .B(KEYINPUT116), .ZN(n548) );
  NAND2_X1 U605 ( .A1(n566), .A2(n548), .ZN(n541) );
  XNOR2_X1 U606 ( .A(G141GAT), .B(n541), .ZN(G1344GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n543) );
  NAND2_X1 U608 ( .A1(n556), .A2(n548), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(n544), .ZN(G1345GAT) );
  XOR2_X1 U611 ( .A(G155GAT), .B(KEYINPUT117), .Z(n546) );
  NAND2_X1 U612 ( .A1(n574), .A2(n548), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(G1346GAT) );
  NAND2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n549), .B(KEYINPUT118), .ZN(n550) );
  XNOR2_X1 U616 ( .A(G162GAT), .B(n550), .ZN(G1347GAT) );
  NAND2_X1 U617 ( .A1(n566), .A2(n551), .ZN(n552) );
  XNOR2_X1 U618 ( .A(G169GAT), .B(n552), .ZN(G1348GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n554) );
  XNOR2_X1 U620 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U622 ( .A(KEYINPUT120), .B(n555), .Z(n558) );
  NAND2_X1 U623 ( .A1(n551), .A2(n556), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1349GAT) );
  AND2_X1 U625 ( .A1(n559), .A2(n551), .ZN(n563) );
  XNOR2_X1 U626 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n560), .B(KEYINPUT123), .ZN(n561) );
  XNOR2_X1 U628 ( .A(KEYINPUT124), .B(n561), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1351GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n568) );
  NOR2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n577) );
  NAND2_X1 U632 ( .A1(n577), .A2(n566), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n572) );
  NAND2_X1 U636 ( .A1(n577), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XOR2_X1 U638 ( .A(G204GAT), .B(n573), .Z(G1353GAT) );
  NAND2_X1 U639 ( .A1(n577), .A2(n574), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(KEYINPUT126), .ZN(n576) );
  XNOR2_X1 U641 ( .A(G211GAT), .B(n576), .ZN(G1354GAT) );
  NAND2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U643 ( .A(n579), .B(KEYINPUT62), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(n580), .ZN(G1355GAT) );
endmodule

