

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600;

  NOR2_X2 U324 ( .A1(n545), .A2(n544), .ZN(n555) );
  XOR2_X1 U325 ( .A(n310), .B(n309), .Z(n542) );
  XNOR2_X1 U326 ( .A(KEYINPUT89), .B(n379), .ZN(n578) );
  XNOR2_X1 U327 ( .A(n345), .B(n435), .ZN(n346) );
  XNOR2_X1 U328 ( .A(n347), .B(n346), .ZN(n348) );
  INV_X1 U329 ( .A(KEYINPUT86), .ZN(n311) );
  XNOR2_X1 U330 ( .A(n311), .B(KEYINPUT21), .ZN(n312) );
  INV_X1 U331 ( .A(KEYINPUT31), .ZN(n455) );
  XNOR2_X1 U332 ( .A(n313), .B(n312), .ZN(n315) );
  XNOR2_X1 U333 ( .A(n456), .B(n455), .ZN(n457) );
  NAND2_X1 U334 ( .A1(n368), .A2(n367), .ZN(n540) );
  XNOR2_X1 U335 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U336 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U337 ( .A(n463), .B(KEYINPUT40), .ZN(n464) );
  XNOR2_X1 U338 ( .A(n491), .B(n490), .ZN(G1351GAT) );
  XNOR2_X1 U339 ( .A(n465), .B(n464), .ZN(G1330GAT) );
  XOR2_X1 U340 ( .A(G127GAT), .B(KEYINPUT0), .Z(n293) );
  XNOR2_X1 U341 ( .A(G113GAT), .B(KEYINPUT82), .ZN(n292) );
  XNOR2_X1 U342 ( .A(n293), .B(n292), .ZN(n334) );
  XOR2_X1 U343 ( .A(n334), .B(G120GAT), .Z(n295) );
  NAND2_X1 U344 ( .A1(G227GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U345 ( .A(n295), .B(n294), .ZN(n310) );
  XOR2_X1 U346 ( .A(G134GAT), .B(G99GAT), .Z(n297) );
  XNOR2_X1 U347 ( .A(G43GAT), .B(G190GAT), .ZN(n296) );
  XNOR2_X1 U348 ( .A(n297), .B(n296), .ZN(n300) );
  XOR2_X1 U349 ( .A(G183GAT), .B(KEYINPUT18), .Z(n299) );
  XNOR2_X1 U350 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n298) );
  XNOR2_X1 U351 ( .A(n299), .B(n298), .ZN(n351) );
  XOR2_X1 U352 ( .A(n300), .B(n351), .Z(n308) );
  XOR2_X1 U353 ( .A(G176GAT), .B(KEYINPUT83), .Z(n302) );
  XNOR2_X1 U354 ( .A(G71GAT), .B(KEYINPUT20), .ZN(n301) );
  XNOR2_X1 U355 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U356 ( .A(KEYINPUT65), .B(KEYINPUT84), .Z(n304) );
  XNOR2_X1 U357 ( .A(G169GAT), .B(G15GAT), .ZN(n303) );
  XNOR2_X1 U358 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U359 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U360 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U361 ( .A(G211GAT), .B(KEYINPUT85), .ZN(n313) );
  XNOR2_X1 U362 ( .A(G197GAT), .B(G218GAT), .ZN(n314) );
  XNOR2_X1 U363 ( .A(n315), .B(n314), .ZN(n347) );
  XOR2_X1 U364 ( .A(KEYINPUT24), .B(KEYINPUT87), .Z(n317) );
  XNOR2_X1 U365 ( .A(G50GAT), .B(KEYINPUT22), .ZN(n316) );
  XNOR2_X1 U366 ( .A(n317), .B(n316), .ZN(n320) );
  XOR2_X1 U367 ( .A(G78GAT), .B(G204GAT), .Z(n319) );
  XNOR2_X1 U368 ( .A(G106GAT), .B(KEYINPUT72), .ZN(n318) );
  XNOR2_X1 U369 ( .A(n319), .B(n318), .ZN(n445) );
  XOR2_X1 U370 ( .A(n320), .B(n445), .Z(n325) );
  XOR2_X1 U371 ( .A(KEYINPUT23), .B(G148GAT), .Z(n322) );
  NAND2_X1 U372 ( .A1(G228GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U373 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U374 ( .A(G22GAT), .B(n323), .ZN(n324) );
  XNOR2_X1 U375 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U376 ( .A(n347), .B(n326), .ZN(n330) );
  XOR2_X1 U377 ( .A(KEYINPUT2), .B(G162GAT), .Z(n328) );
  XNOR2_X1 U378 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n327) );
  XNOR2_X1 U379 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U380 ( .A(G141GAT), .B(n329), .Z(n342) );
  XOR2_X1 U381 ( .A(n330), .B(n342), .Z(n484) );
  XOR2_X1 U382 ( .A(KEYINPUT28), .B(n484), .Z(n536) );
  INV_X1 U383 ( .A(n536), .ZN(n545) );
  XNOR2_X1 U384 ( .A(G120GAT), .B(G148GAT), .ZN(n331) );
  XNOR2_X1 U385 ( .A(n331), .B(G57GAT), .ZN(n451) );
  XOR2_X1 U386 ( .A(KEYINPUT88), .B(n451), .Z(n333) );
  XOR2_X1 U387 ( .A(G29GAT), .B(G134GAT), .Z(n388) );
  XNOR2_X1 U388 ( .A(G85GAT), .B(n388), .ZN(n332) );
  XNOR2_X1 U389 ( .A(n333), .B(n332), .ZN(n338) );
  XOR2_X1 U390 ( .A(n334), .B(KEYINPUT6), .Z(n336) );
  NAND2_X1 U391 ( .A1(G225GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U392 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U393 ( .A(n338), .B(n337), .Z(n344) );
  XOR2_X1 U394 ( .A(KEYINPUT4), .B(KEYINPUT1), .Z(n340) );
  XNOR2_X1 U395 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n339) );
  XNOR2_X1 U396 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U397 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U398 ( .A(n344), .B(n343), .ZN(n379) );
  XOR2_X1 U399 ( .A(G36GAT), .B(G190GAT), .Z(n387) );
  XOR2_X1 U400 ( .A(KEYINPUT90), .B(G204GAT), .Z(n345) );
  XOR2_X1 U401 ( .A(G169GAT), .B(G8GAT), .Z(n435) );
  XOR2_X1 U402 ( .A(n387), .B(n348), .Z(n350) );
  NAND2_X1 U403 ( .A1(G226GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U404 ( .A(n350), .B(n349), .ZN(n352) );
  NAND2_X1 U405 ( .A1(n352), .A2(n351), .ZN(n356) );
  INV_X1 U406 ( .A(n351), .ZN(n354) );
  INV_X1 U407 ( .A(n352), .ZN(n353) );
  NAND2_X1 U408 ( .A1(n354), .A2(n353), .ZN(n355) );
  NAND2_X1 U409 ( .A1(n356), .A2(n355), .ZN(n362) );
  INV_X1 U410 ( .A(G92GAT), .ZN(n357) );
  NAND2_X1 U411 ( .A1(G176GAT), .A2(n357), .ZN(n360) );
  INV_X1 U412 ( .A(G176GAT), .ZN(n358) );
  NAND2_X1 U413 ( .A1(n358), .A2(G92GAT), .ZN(n359) );
  NAND2_X1 U414 ( .A1(n360), .A2(n359), .ZN(n361) );
  XOR2_X1 U415 ( .A(G64GAT), .B(n361), .Z(n449) );
  XOR2_X1 U416 ( .A(n362), .B(n449), .Z(n363) );
  INV_X1 U417 ( .A(n363), .ZN(n480) );
  XNOR2_X1 U418 ( .A(KEYINPUT27), .B(n480), .ZN(n372) );
  OR2_X1 U419 ( .A1(n578), .A2(n372), .ZN(n364) );
  NAND2_X1 U420 ( .A1(n364), .A2(KEYINPUT91), .ZN(n368) );
  INV_X1 U421 ( .A(KEYINPUT91), .ZN(n366) );
  NOR2_X1 U422 ( .A1(n578), .A2(n372), .ZN(n365) );
  NAND2_X1 U423 ( .A1(n366), .A2(n365), .ZN(n367) );
  NAND2_X1 U424 ( .A1(n542), .A2(n540), .ZN(n369) );
  NOR2_X1 U425 ( .A1(n545), .A2(n369), .ZN(n370) );
  XNOR2_X1 U426 ( .A(n370), .B(KEYINPUT92), .ZN(n381) );
  NAND2_X1 U427 ( .A1(n484), .A2(n542), .ZN(n371) );
  XNOR2_X1 U428 ( .A(n371), .B(KEYINPUT26), .ZN(n581) );
  NOR2_X1 U429 ( .A1(n581), .A2(n372), .ZN(n377) );
  NOR2_X1 U430 ( .A1(n542), .A2(n480), .ZN(n373) );
  NOR2_X1 U431 ( .A1(n484), .A2(n373), .ZN(n374) );
  XNOR2_X1 U432 ( .A(n374), .B(KEYINPUT93), .ZN(n375) );
  XNOR2_X1 U433 ( .A(n375), .B(KEYINPUT25), .ZN(n376) );
  NOR2_X1 U434 ( .A1(n377), .A2(n376), .ZN(n378) );
  NOR2_X1 U435 ( .A1(n379), .A2(n378), .ZN(n380) );
  NOR2_X1 U436 ( .A1(n381), .A2(n380), .ZN(n497) );
  XOR2_X1 U437 ( .A(KEYINPUT8), .B(KEYINPUT69), .Z(n383) );
  XNOR2_X1 U438 ( .A(G50GAT), .B(G43GAT), .ZN(n382) );
  XNOR2_X1 U439 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U440 ( .A(KEYINPUT7), .B(n384), .ZN(n439) );
  INV_X1 U441 ( .A(n439), .ZN(n402) );
  XOR2_X1 U442 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n386) );
  XNOR2_X1 U443 ( .A(G106GAT), .B(KEYINPUT9), .ZN(n385) );
  XNOR2_X1 U444 ( .A(n386), .B(n385), .ZN(n400) );
  XOR2_X1 U445 ( .A(G92GAT), .B(n387), .Z(n390) );
  XNOR2_X1 U446 ( .A(G162GAT), .B(n388), .ZN(n389) );
  XNOR2_X1 U447 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U448 ( .A(n391), .B(KEYINPUT64), .Z(n398) );
  XOR2_X1 U449 ( .A(G99GAT), .B(G85GAT), .Z(n392) );
  XOR2_X1 U450 ( .A(KEYINPUT73), .B(n392), .Z(n444) );
  INV_X1 U451 ( .A(n444), .ZN(n393) );
  XNOR2_X1 U452 ( .A(n393), .B(KEYINPUT76), .ZN(n395) );
  NAND2_X1 U453 ( .A1(G232GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U454 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U455 ( .A(G218GAT), .B(n396), .ZN(n397) );
  XNOR2_X1 U456 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U457 ( .A(n400), .B(n399), .Z(n401) );
  XOR2_X1 U458 ( .A(n402), .B(n401), .Z(n567) );
  INV_X1 U459 ( .A(n567), .ZN(n469) );
  XOR2_X1 U460 ( .A(KEYINPUT36), .B(KEYINPUT98), .Z(n403) );
  XOR2_X1 U461 ( .A(n469), .B(n403), .Z(n598) );
  XOR2_X1 U462 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n405) );
  XNOR2_X1 U463 ( .A(KEYINPUT80), .B(KEYINPUT81), .ZN(n404) );
  XNOR2_X1 U464 ( .A(n405), .B(n404), .ZN(n417) );
  XOR2_X1 U465 ( .A(G78GAT), .B(G155GAT), .Z(n407) );
  XNOR2_X1 U466 ( .A(G127GAT), .B(G211GAT), .ZN(n406) );
  XNOR2_X1 U467 ( .A(n407), .B(n406), .ZN(n415) );
  XOR2_X1 U468 ( .A(KEYINPUT15), .B(KEYINPUT78), .Z(n409) );
  XNOR2_X1 U469 ( .A(KEYINPUT77), .B(KEYINPUT79), .ZN(n408) );
  XNOR2_X1 U470 ( .A(n409), .B(n408), .ZN(n413) );
  XOR2_X1 U471 ( .A(G64GAT), .B(G57GAT), .Z(n411) );
  XNOR2_X1 U472 ( .A(G8GAT), .B(G183GAT), .ZN(n410) );
  XNOR2_X1 U473 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U474 ( .A(n413), .B(n412), .Z(n414) );
  XNOR2_X1 U475 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U476 ( .A(n417), .B(n416), .ZN(n422) );
  XOR2_X1 U477 ( .A(G71GAT), .B(KEYINPUT13), .Z(n454) );
  XNOR2_X1 U478 ( .A(G22GAT), .B(G15GAT), .ZN(n418) );
  XNOR2_X1 U479 ( .A(n418), .B(G1GAT), .ZN(n434) );
  XOR2_X1 U480 ( .A(n454), .B(n434), .Z(n420) );
  NAND2_X1 U481 ( .A1(G231GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U482 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U483 ( .A(n422), .B(n421), .Z(n591) );
  OR2_X1 U484 ( .A1(n598), .A2(n591), .ZN(n423) );
  OR2_X1 U485 ( .A1(n497), .A2(n423), .ZN(n425) );
  XOR2_X1 U486 ( .A(KEYINPUT99), .B(KEYINPUT37), .Z(n424) );
  XNOR2_X1 U487 ( .A(n425), .B(n424), .ZN(n527) );
  XOR2_X1 U488 ( .A(KEYINPUT70), .B(KEYINPUT29), .Z(n427) );
  XNOR2_X1 U489 ( .A(KEYINPUT66), .B(KEYINPUT71), .ZN(n426) );
  XNOR2_X1 U490 ( .A(n427), .B(n426), .ZN(n443) );
  XOR2_X1 U491 ( .A(G141GAT), .B(G197GAT), .Z(n429) );
  XNOR2_X1 U492 ( .A(G29GAT), .B(G36GAT), .ZN(n428) );
  XNOR2_X1 U493 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U494 ( .A(KEYINPUT67), .B(KEYINPUT30), .Z(n431) );
  XNOR2_X1 U495 ( .A(G113GAT), .B(KEYINPUT68), .ZN(n430) );
  XNOR2_X1 U496 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U497 ( .A(n433), .B(n432), .Z(n441) );
  XOR2_X1 U498 ( .A(n435), .B(n434), .Z(n437) );
  NAND2_X1 U499 ( .A1(G229GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U500 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U501 ( .A(n439), .B(n438), .Z(n440) );
  XNOR2_X1 U502 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U503 ( .A(n443), .B(n442), .ZN(n582) );
  INV_X1 U504 ( .A(n582), .ZN(n475) );
  XOR2_X1 U505 ( .A(n445), .B(n444), .Z(n460) );
  XOR2_X1 U506 ( .A(KEYINPUT33), .B(KEYINPUT75), .Z(n447) );
  NAND2_X1 U507 ( .A1(G230GAT), .A2(G233GAT), .ZN(n446) );
  XNOR2_X1 U508 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U509 ( .A(n448), .B(KEYINPUT32), .Z(n453) );
  INV_X1 U510 ( .A(n449), .ZN(n450) );
  XOR2_X1 U511 ( .A(n451), .B(n450), .Z(n452) );
  XNOR2_X1 U512 ( .A(n453), .B(n452), .ZN(n458) );
  XNOR2_X1 U513 ( .A(n454), .B(KEYINPUT74), .ZN(n456) );
  XNOR2_X1 U514 ( .A(n460), .B(n459), .ZN(n587) );
  NOR2_X1 U515 ( .A1(n475), .A2(n587), .ZN(n499) );
  NAND2_X1 U516 ( .A1(n527), .A2(n499), .ZN(n462) );
  XNOR2_X1 U517 ( .A(KEYINPUT100), .B(KEYINPUT38), .ZN(n461) );
  XNOR2_X1 U518 ( .A(n462), .B(n461), .ZN(n513) );
  NOR2_X1 U519 ( .A1(n542), .A2(n513), .ZN(n465) );
  INV_X1 U520 ( .A(G43GAT), .ZN(n463) );
  XOR2_X1 U521 ( .A(KEYINPUT54), .B(KEYINPUT120), .Z(n482) );
  XOR2_X1 U522 ( .A(KEYINPUT41), .B(n587), .Z(n571) );
  INV_X1 U523 ( .A(n571), .ZN(n515) );
  NOR2_X1 U524 ( .A1(n515), .A2(n475), .ZN(n466) );
  XNOR2_X1 U525 ( .A(n466), .B(KEYINPUT46), .ZN(n467) );
  NOR2_X1 U526 ( .A1(n591), .A2(n467), .ZN(n468) );
  XNOR2_X1 U527 ( .A(n468), .B(KEYINPUT110), .ZN(n470) );
  NAND2_X1 U528 ( .A1(n470), .A2(n469), .ZN(n472) );
  XNOR2_X1 U529 ( .A(KEYINPUT111), .B(KEYINPUT47), .ZN(n471) );
  XNOR2_X1 U530 ( .A(n472), .B(n471), .ZN(n478) );
  INV_X1 U531 ( .A(n591), .ZN(n494) );
  NOR2_X1 U532 ( .A1(n494), .A2(n598), .ZN(n473) );
  XOR2_X1 U533 ( .A(KEYINPUT45), .B(n473), .Z(n474) );
  NOR2_X1 U534 ( .A1(n587), .A2(n474), .ZN(n476) );
  NAND2_X1 U535 ( .A1(n476), .A2(n475), .ZN(n477) );
  NAND2_X1 U536 ( .A1(n478), .A2(n477), .ZN(n479) );
  XNOR2_X1 U537 ( .A(n479), .B(KEYINPUT48), .ZN(n541) );
  NAND2_X1 U538 ( .A1(n541), .A2(n363), .ZN(n481) );
  XNOR2_X1 U539 ( .A(n482), .B(n481), .ZN(n579) );
  INV_X1 U540 ( .A(n578), .ZN(n483) );
  NOR2_X1 U541 ( .A1(n484), .A2(n483), .ZN(n485) );
  AND2_X1 U542 ( .A1(n579), .A2(n485), .ZN(n486) );
  XNOR2_X1 U543 ( .A(n486), .B(KEYINPUT55), .ZN(n487) );
  NOR2_X2 U544 ( .A1(n542), .A2(n487), .ZN(n576) );
  NAND2_X1 U545 ( .A1(n576), .A2(n567), .ZN(n491) );
  XOR2_X1 U546 ( .A(KEYINPUT58), .B(KEYINPUT122), .Z(n489) );
  INV_X1 U547 ( .A(G190GAT), .ZN(n488) );
  XOR2_X1 U548 ( .A(KEYINPUT95), .B(KEYINPUT34), .Z(n493) );
  XNOR2_X1 U549 ( .A(G1GAT), .B(KEYINPUT96), .ZN(n492) );
  XNOR2_X1 U550 ( .A(n493), .B(n492), .ZN(n501) );
  NOR2_X1 U551 ( .A1(n567), .A2(n494), .ZN(n495) );
  XOR2_X1 U552 ( .A(KEYINPUT16), .B(n495), .Z(n496) );
  NOR2_X1 U553 ( .A1(n497), .A2(n496), .ZN(n498) );
  XNOR2_X1 U554 ( .A(KEYINPUT94), .B(n498), .ZN(n516) );
  NAND2_X1 U555 ( .A1(n499), .A2(n516), .ZN(n506) );
  NOR2_X1 U556 ( .A1(n578), .A2(n506), .ZN(n500) );
  XOR2_X1 U557 ( .A(n501), .B(n500), .Z(G1324GAT) );
  NOR2_X1 U558 ( .A1(n480), .A2(n506), .ZN(n503) );
  XNOR2_X1 U559 ( .A(G8GAT), .B(KEYINPUT97), .ZN(n502) );
  XNOR2_X1 U560 ( .A(n503), .B(n502), .ZN(G1325GAT) );
  NOR2_X1 U561 ( .A1(n542), .A2(n506), .ZN(n505) );
  XNOR2_X1 U562 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n504) );
  XNOR2_X1 U563 ( .A(n505), .B(n504), .ZN(G1326GAT) );
  NOR2_X1 U564 ( .A1(n536), .A2(n506), .ZN(n507) );
  XOR2_X1 U565 ( .A(G22GAT), .B(n507), .Z(G1327GAT) );
  NOR2_X1 U566 ( .A1(n578), .A2(n513), .ZN(n509) );
  XNOR2_X1 U567 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n508) );
  XNOR2_X1 U568 ( .A(n509), .B(n508), .ZN(G1328GAT) );
  NOR2_X1 U569 ( .A1(n480), .A2(n513), .ZN(n511) );
  XNOR2_X1 U570 ( .A(KEYINPUT101), .B(KEYINPUT102), .ZN(n510) );
  XNOR2_X1 U571 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U572 ( .A(G36GAT), .B(n512), .ZN(G1329GAT) );
  NOR2_X1 U573 ( .A1(n536), .A2(n513), .ZN(n514) );
  XOR2_X1 U574 ( .A(G50GAT), .B(n514), .Z(G1331GAT) );
  NOR2_X1 U575 ( .A1(n515), .A2(n582), .ZN(n528) );
  NAND2_X1 U576 ( .A1(n528), .A2(n516), .ZN(n523) );
  NOR2_X1 U577 ( .A1(n578), .A2(n523), .ZN(n518) );
  XNOR2_X1 U578 ( .A(KEYINPUT103), .B(KEYINPUT42), .ZN(n517) );
  XNOR2_X1 U579 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U580 ( .A(G57GAT), .B(n519), .ZN(G1332GAT) );
  NOR2_X1 U581 ( .A1(n480), .A2(n523), .ZN(n520) );
  XOR2_X1 U582 ( .A(KEYINPUT104), .B(n520), .Z(n521) );
  XNOR2_X1 U583 ( .A(G64GAT), .B(n521), .ZN(G1333GAT) );
  NOR2_X1 U584 ( .A1(n542), .A2(n523), .ZN(n522) );
  XOR2_X1 U585 ( .A(G71GAT), .B(n522), .Z(G1334GAT) );
  NOR2_X1 U586 ( .A1(n536), .A2(n523), .ZN(n525) );
  XNOR2_X1 U587 ( .A(KEYINPUT105), .B(KEYINPUT43), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U589 ( .A(G78GAT), .B(n526), .Z(G1335GAT) );
  NAND2_X1 U590 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U591 ( .A(n529), .B(KEYINPUT106), .ZN(n537) );
  NOR2_X1 U592 ( .A1(n537), .A2(n578), .ZN(n530) );
  XOR2_X1 U593 ( .A(G85GAT), .B(n530), .Z(G1336GAT) );
  NOR2_X1 U594 ( .A1(n480), .A2(n537), .ZN(n531) );
  XOR2_X1 U595 ( .A(G92GAT), .B(n531), .Z(G1337GAT) );
  XNOR2_X1 U596 ( .A(G99GAT), .B(KEYINPUT107), .ZN(n533) );
  NOR2_X1 U597 ( .A1(n542), .A2(n537), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(G1338GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT108), .B(KEYINPUT44), .Z(n535) );
  XNOR2_X1 U600 ( .A(G106GAT), .B(KEYINPUT109), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n535), .B(n534), .ZN(n539) );
  NOR2_X1 U602 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U603 ( .A(n539), .B(n538), .Z(G1339GAT) );
  XOR2_X1 U604 ( .A(G113GAT), .B(KEYINPUT113), .Z(n547) );
  NAND2_X1 U605 ( .A1(n541), .A2(n540), .ZN(n560) );
  NOR2_X1 U606 ( .A1(n542), .A2(n560), .ZN(n543) );
  XOR2_X1 U607 ( .A(KEYINPUT112), .B(n543), .Z(n544) );
  NAND2_X1 U608 ( .A1(n555), .A2(n582), .ZN(n546) );
  XNOR2_X1 U609 ( .A(n547), .B(n546), .ZN(G1340GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n549) );
  NAND2_X1 U611 ( .A1(n555), .A2(n571), .ZN(n548) );
  XNOR2_X1 U612 ( .A(n549), .B(n548), .ZN(n551) );
  XOR2_X1 U613 ( .A(G120GAT), .B(KEYINPUT114), .Z(n550) );
  XNOR2_X1 U614 ( .A(n551), .B(n550), .ZN(G1341GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n553) );
  NAND2_X1 U616 ( .A1(n555), .A2(n591), .ZN(n552) );
  XNOR2_X1 U617 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U618 ( .A(G127GAT), .B(n554), .Z(G1342GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n557) );
  NAND2_X1 U620 ( .A1(n555), .A2(n567), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n557), .B(n556), .ZN(n559) );
  XOR2_X1 U622 ( .A(G134GAT), .B(KEYINPUT117), .Z(n558) );
  XNOR2_X1 U623 ( .A(n559), .B(n558), .ZN(G1343GAT) );
  NOR2_X1 U624 ( .A1(n581), .A2(n560), .ZN(n561) );
  XOR2_X1 U625 ( .A(KEYINPUT119), .B(n561), .Z(n568) );
  NAND2_X1 U626 ( .A1(n568), .A2(n582), .ZN(n562) );
  XNOR2_X1 U627 ( .A(G141GAT), .B(n562), .ZN(G1344GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n564) );
  NAND2_X1 U629 ( .A1(n568), .A2(n571), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(G148GAT), .B(n565), .ZN(G1345GAT) );
  NAND2_X1 U632 ( .A1(n568), .A2(n591), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n566), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U636 ( .A1(n576), .A2(n582), .ZN(n570) );
  XNOR2_X1 U637 ( .A(G169GAT), .B(n570), .ZN(G1348GAT) );
  XOR2_X1 U638 ( .A(G176GAT), .B(KEYINPUT57), .Z(n573) );
  NAND2_X1 U639 ( .A1(n576), .A2(n571), .ZN(n572) );
  XNOR2_X1 U640 ( .A(n573), .B(n572), .ZN(n575) );
  XOR2_X1 U641 ( .A(KEYINPUT121), .B(KEYINPUT56), .Z(n574) );
  XNOR2_X1 U642 ( .A(n575), .B(n574), .ZN(G1349GAT) );
  NAND2_X1 U643 ( .A1(n576), .A2(n591), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n577), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U645 ( .A(G197GAT), .B(KEYINPUT123), .Z(n584) );
  NAND2_X1 U646 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U647 ( .A1(n581), .A2(n580), .ZN(n596) );
  NAND2_X1 U648 ( .A1(n596), .A2(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(n586) );
  XOR2_X1 U650 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1352GAT) );
  XOR2_X1 U652 ( .A(KEYINPUT61), .B(KEYINPUT124), .Z(n589) );
  NAND2_X1 U653 ( .A1(n596), .A2(n587), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U655 ( .A(G204GAT), .B(n590), .ZN(G1353GAT) );
  XOR2_X1 U656 ( .A(G211GAT), .B(KEYINPUT125), .Z(n593) );
  NAND2_X1 U657 ( .A1(n596), .A2(n591), .ZN(n592) );
  XNOR2_X1 U658 ( .A(n593), .B(n592), .ZN(G1354GAT) );
  XOR2_X1 U659 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n595) );
  XNOR2_X1 U660 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n594) );
  XNOR2_X1 U661 ( .A(n595), .B(n594), .ZN(n600) );
  INV_X1 U662 ( .A(n596), .ZN(n597) );
  NOR2_X1 U663 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X1 U664 ( .A(n600), .B(n599), .Z(G1355GAT) );
endmodule

