//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 1 1 0 1 1 1 0 1 1 1 1 0 0 1 1 0 0 1 1 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n450, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n609, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187, new_n1188;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT64), .B(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT65), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n453), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI211_X1 g043(.A(G137), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n463), .A2(G101), .A3(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n468), .A2(new_n471), .ZN(G160));
  NOR2_X1   g047(.A1(new_n464), .A2(new_n465), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  OR2_X1    g049(.A1(new_n474), .A2(KEYINPUT66), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(KEYINPUT66), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  NOR2_X1   g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT67), .ZN(new_n481));
  INV_X1    g056(.A(G2104), .ZN(new_n482));
  INV_X1    g057(.A(G112), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(new_n465), .ZN(new_n485));
  NAND2_X1  g060(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n463), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AOI22_X1  g062(.A1(new_n481), .A2(new_n484), .B1(new_n487), .B2(G124), .ZN(new_n488));
  AND2_X1   g063(.A1(new_n479), .A2(new_n488), .ZN(G162));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(KEYINPUT70), .C1(new_n465), .C2(new_n464), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT69), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n491), .B(new_n494), .C1(new_n465), .C2(new_n464), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n493), .A2(KEYINPUT4), .A3(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n492), .A2(KEYINPUT69), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT68), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n463), .A2(G114), .ZN(new_n500));
  OAI21_X1  g075(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OR2_X1    g077(.A1(G102), .A2(G2105), .ZN(new_n503));
  INV_X1    g078(.A(G114), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G2105), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n503), .A2(new_n505), .A3(KEYINPUT68), .A4(G2104), .ZN(new_n506));
  AOI22_X1  g081(.A1(G126), .A2(new_n487), .B1(new_n502), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n496), .A2(new_n498), .A3(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT71), .B1(new_n510), .B2(KEYINPUT6), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(new_n513), .A3(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n510), .A2(KEYINPUT6), .ZN(new_n516));
  NAND4_X1  g091(.A1(new_n515), .A2(G50), .A3(G543), .A4(new_n516), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT72), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  OR2_X1    g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G62), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n519), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n515), .A2(new_n516), .A3(new_n522), .ZN(new_n526));
  AOI22_X1  g101(.A1(G651), .A2(new_n525), .B1(new_n526), .B2(G88), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n518), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(KEYINPUT73), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT73), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n518), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n529), .A2(new_n531), .ZN(G166));
  NAND2_X1  g107(.A1(new_n526), .A2(G89), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n515), .A2(G51), .A3(G543), .A4(new_n516), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n537));
  AND2_X1   g112(.A1(G63), .A2(G651), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n536), .A2(new_n537), .B1(new_n522), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n533), .A2(new_n534), .A3(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(G168));
  AOI22_X1  g116(.A1(new_n522), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(new_n510), .ZN(new_n543));
  XOR2_X1   g118(.A(KEYINPUT74), .B(G90), .Z(new_n544));
  NAND2_X1  g119(.A1(new_n526), .A2(new_n544), .ZN(new_n545));
  AND3_X1   g120(.A1(new_n515), .A2(G543), .A3(new_n516), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G52), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n543), .A2(new_n545), .A3(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  AOI22_X1  g124(.A1(new_n522), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(new_n510), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n546), .A2(G43), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n515), .A2(G81), .A3(new_n516), .A4(new_n522), .ZN(new_n553));
  AND3_X1   g128(.A1(new_n552), .A2(KEYINPUT75), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g129(.A(KEYINPUT75), .B1(new_n552), .B2(new_n553), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n551), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(new_n522), .A2(G65), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT76), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G651), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(KEYINPUT77), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n510), .B1(new_n563), .B2(new_n565), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT77), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n568), .A2(new_n571), .B1(G91), .B2(new_n526), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n515), .A2(G53), .A3(G543), .A4(new_n516), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT9), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n574), .ZN(G299));
  XNOR2_X1  g150(.A(new_n540), .B(KEYINPUT78), .ZN(G286));
  INV_X1    g151(.A(G166), .ZN(G303));
  NAND2_X1  g152(.A1(new_n546), .A2(G49), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n526), .A2(G87), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n522), .B2(G74), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G288));
  NAND2_X1  g156(.A1(new_n526), .A2(G86), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n546), .A2(G48), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n522), .A2(G61), .ZN(new_n585));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n584), .B1(new_n587), .B2(G651), .ZN(new_n588));
  AOI211_X1 g163(.A(KEYINPUT79), .B(new_n510), .C1(new_n585), .C2(new_n586), .ZN(new_n589));
  OAI211_X1 g164(.A(new_n582), .B(new_n583), .C1(new_n588), .C2(new_n589), .ZN(G305));
  AOI22_X1  g165(.A1(new_n522), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  OR2_X1    g166(.A1(new_n591), .A2(new_n510), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n526), .A2(G85), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n546), .A2(G47), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(G301), .A2(G868), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n515), .A2(G92), .A3(new_n516), .A4(new_n522), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n597), .B(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n523), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(G651), .A2(new_n602), .B1(new_n546), .B2(G54), .ZN(new_n603));
  AND2_X1   g178(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n596), .B1(new_n604), .B2(G868), .ZN(G321));
  XOR2_X1   g180(.A(G321), .B(KEYINPUT80), .Z(G284));
  MUX2_X1   g181(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g182(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n604), .B1(new_n609), .B2(G860), .ZN(G148));
  NAND2_X1  g185(.A1(new_n599), .A2(new_n603), .ZN(new_n611));
  OAI21_X1  g186(.A(G868), .B1(new_n611), .B2(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G868), .B2(new_n557), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g189(.A1(new_n478), .A2(G135), .ZN(new_n615));
  OR3_X1    g190(.A1(new_n463), .A2(KEYINPUT83), .A3(G111), .ZN(new_n616));
  OAI21_X1  g191(.A(KEYINPUT83), .B1(new_n463), .B2(G111), .ZN(new_n617));
  OR2_X1    g192(.A1(G99), .A2(G2105), .ZN(new_n618));
  NAND4_X1  g193(.A1(new_n616), .A2(G2104), .A3(new_n617), .A4(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n487), .A2(G123), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT82), .Z(new_n621));
  AND3_X1   g196(.A1(new_n615), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n623), .A2(G2096), .ZN(new_n624));
  XOR2_X1   g199(.A(KEYINPUT81), .B(KEYINPUT12), .Z(new_n625));
  NAND3_X1  g200(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2100), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n623), .A2(G2096), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n624), .A2(new_n629), .A3(new_n630), .ZN(G156));
  INV_X1    g206(.A(KEYINPUT14), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2427), .B(G2438), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2430), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2435), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n632), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(new_n635), .B2(new_n634), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT85), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n637), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2451), .B(G2454), .Z(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n642), .A2(new_n645), .ZN(new_n647));
  AND3_X1   g222(.A1(new_n646), .A2(G14), .A3(new_n647), .ZN(G401));
  XNOR2_X1  g223(.A(G2067), .B(G2678), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT86), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2084), .B(G2090), .ZN(new_n652));
  NOR2_X1   g227(.A1(G2072), .A2(G2078), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n442), .A2(new_n653), .ZN(new_n654));
  NOR3_X1   g229(.A1(new_n651), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT87), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT18), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n654), .B(KEYINPUT17), .Z(new_n658));
  NOR3_X1   g233(.A1(new_n658), .A2(new_n650), .A3(new_n652), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT89), .Z(new_n660));
  INV_X1    g235(.A(new_n652), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(new_n651), .B2(new_n654), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT88), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n658), .A2(new_n650), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n660), .B1(new_n664), .B2(new_n667), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n657), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(G2100), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT90), .B(G2096), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G227));
  XOR2_X1   g247(.A(G1971), .B(G1976), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  XOR2_X1   g249(.A(G1956), .B(G2474), .Z(new_n675));
  XOR2_X1   g250(.A(G1961), .B(G1966), .Z(new_n676));
  AND2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT20), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n675), .A2(new_n676), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  MUX2_X1   g257(.A(new_n682), .B(new_n681), .S(new_n674), .Z(new_n683));
  NOR2_X1   g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1991), .B(G1996), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(G229));
  INV_X1    g266(.A(G29), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n692), .A2(KEYINPUT91), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(KEYINPUT91), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n695), .A2(G35), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(G162), .B2(new_n695), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT29), .ZN(new_n698));
  AND2_X1   g273(.A1(new_n698), .A2(G2090), .ZN(new_n699));
  INV_X1    g274(.A(new_n695), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G27), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(G164), .B2(new_n700), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(G2078), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n692), .A2(G33), .ZN(new_n704));
  NAND2_X1  g279(.A1(G115), .A2(G2104), .ZN(new_n705));
  INV_X1    g280(.A(G127), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(new_n473), .B2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT25), .ZN(new_n708));
  NAND2_X1  g283(.A1(G103), .A2(G2104), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(G2105), .ZN(new_n710));
  NAND4_X1  g285(.A1(new_n463), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n711));
  AOI22_X1  g286(.A1(new_n707), .A2(G2105), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G139), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n477), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n704), .B1(new_n714), .B2(G29), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G2072), .ZN(new_n716));
  NAND2_X1  g291(.A1(G160), .A2(G29), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT24), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n718), .A2(G34), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(G34), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n700), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n717), .A2(G2084), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n622), .A2(new_n695), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT31), .B(G11), .Z(new_n724));
  XOR2_X1   g299(.A(KEYINPUT102), .B(G28), .Z(new_n725));
  NOR2_X1   g300(.A1(new_n725), .A2(KEYINPUT30), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n726), .A2(G29), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n725), .A2(KEYINPUT30), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n724), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n716), .A2(new_n722), .A3(new_n723), .A4(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n604), .A2(G16), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G4), .B2(G16), .ZN(new_n732));
  INV_X1    g307(.A(G1348), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR4_X1   g309(.A1(new_n699), .A2(new_n703), .A3(new_n730), .A4(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n732), .A2(new_n733), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n478), .A2(G141), .ZN(new_n737));
  NAND3_X1  g312(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT100), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT26), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n487), .A2(G129), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n463), .A2(G105), .A3(G2104), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n739), .A2(new_n740), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n737), .A2(G29), .A3(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT101), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n747), .B(new_n748), .C1(G29), .C2(G32), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n748), .B2(new_n747), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT27), .B(G1996), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n736), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n752), .B2(new_n750), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT104), .ZN(new_n755));
  OR3_X1    g330(.A1(new_n698), .A2(new_n755), .A3(G2090), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n755), .B1(new_n698), .B2(G2090), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n754), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G16), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G20), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT23), .Z(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G299), .B2(G16), .ZN(new_n762));
  INV_X1    g337(.A(G1956), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(G16), .A2(G19), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n557), .B2(G16), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n766), .A2(G1341), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n766), .A2(G1341), .ZN(new_n768));
  NOR3_X1   g343(.A1(new_n764), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  AND3_X1   g344(.A1(new_n700), .A2(KEYINPUT28), .A3(G26), .ZN(new_n770));
  AOI21_X1  g345(.A(KEYINPUT28), .B1(new_n700), .B2(G26), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n487), .A2(G128), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT97), .Z(new_n773));
  OAI21_X1  g348(.A(KEYINPUT98), .B1(G104), .B2(G2105), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  NOR3_X1   g350(.A1(KEYINPUT98), .A2(G104), .A3(G2105), .ZN(new_n776));
  OAI221_X1 g351(.A(G2104), .B1(G116), .B2(new_n463), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(G140), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n773), .B(new_n777), .C1(new_n778), .C2(new_n477), .ZN(new_n779));
  AOI211_X1 g354(.A(new_n770), .B(new_n771), .C1(new_n779), .C2(G29), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT99), .B(G2067), .Z(new_n781));
  AND2_X1   g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n759), .A2(G5), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G171), .B2(new_n759), .ZN(new_n784));
  OAI22_X1  g359(.A1(new_n780), .A2(new_n781), .B1(G1961), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n759), .A2(G21), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G168), .B2(new_n759), .ZN(new_n787));
  AOI22_X1  g362(.A1(new_n784), .A2(G1961), .B1(new_n787), .B2(G1966), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G1966), .B2(new_n787), .ZN(new_n789));
  AOI21_X1  g364(.A(G2084), .B1(new_n717), .B2(new_n721), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT103), .ZN(new_n791));
  NOR4_X1   g366(.A1(new_n782), .A2(new_n785), .A3(new_n789), .A4(new_n791), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n735), .A2(new_n758), .A3(new_n769), .A4(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT105), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n759), .A2(G6), .ZN(new_n797));
  INV_X1    g372(.A(G305), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(new_n798), .B2(new_n759), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT94), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT32), .B(G1981), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(G16), .A2(G22), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G166), .B2(G16), .ZN(new_n804));
  INV_X1    g379(.A(G1971), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n759), .A2(G23), .ZN(new_n807));
  NAND2_X1  g382(.A1(G288), .A2(KEYINPUT95), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT95), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n578), .A2(new_n579), .A3(new_n809), .A4(new_n580), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n807), .B1(new_n812), .B2(new_n759), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT33), .B(G1976), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT96), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n813), .B(new_n815), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n802), .A2(new_n806), .A3(new_n816), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT93), .B(KEYINPUT34), .Z(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n817), .A2(new_n819), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n695), .A2(G25), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n478), .A2(G131), .ZN(new_n823));
  OAI21_X1  g398(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n824));
  INV_X1    g399(.A(G107), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n824), .B1(new_n825), .B2(G2105), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(new_n487), .B2(G119), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n823), .A2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n822), .B1(new_n829), .B2(new_n695), .ZN(new_n830));
  XOR2_X1   g405(.A(KEYINPUT35), .B(G1991), .Z(new_n831));
  XOR2_X1   g406(.A(new_n830), .B(new_n831), .Z(new_n832));
  NAND2_X1  g407(.A1(new_n759), .A2(G24), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT92), .ZN(new_n834));
  INV_X1    g409(.A(G290), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n835), .B2(new_n759), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G1986), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n832), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n820), .A2(new_n821), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(KEYINPUT36), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT36), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n820), .A2(new_n841), .A3(new_n821), .A4(new_n838), .ZN(new_n842));
  AOI22_X1  g417(.A1(new_n795), .A2(new_n796), .B1(new_n840), .B2(new_n842), .ZN(G311));
  NAND2_X1  g418(.A1(new_n795), .A2(new_n796), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n840), .A2(new_n842), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(G150));
  XOR2_X1   g421(.A(KEYINPUT106), .B(KEYINPUT38), .Z(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n556), .A2(KEYINPUT107), .ZN(new_n849));
  AOI22_X1  g424(.A1(new_n522), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n850), .A2(new_n510), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n526), .A2(G93), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n546), .A2(G55), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT107), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n856), .B(new_n551), .C1(new_n554), .C2(new_n555), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n849), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n611), .A2(new_n609), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n556), .A2(KEYINPUT107), .A3(new_n854), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n858), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n860), .B1(new_n858), .B2(new_n861), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n848), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n864), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n866), .A2(new_n847), .A3(new_n862), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(KEYINPUT39), .ZN(new_n869));
  INV_X1    g444(.A(G860), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT39), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n865), .A2(new_n867), .A3(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n869), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(KEYINPUT108), .Z(new_n874));
  NAND2_X1  g449(.A1(new_n854), .A2(G860), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n875), .B(KEYINPUT109), .Z(new_n876));
  XOR2_X1   g451(.A(new_n876), .B(KEYINPUT37), .Z(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(G145));
  XNOR2_X1  g453(.A(KEYINPUT111), .B(G37), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n737), .A2(new_n746), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n714), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n828), .B(new_n627), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n881), .B(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n779), .B(new_n508), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n487), .A2(G130), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n463), .A2(G118), .ZN(new_n886));
  OAI21_X1  g461(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n888), .B1(new_n478), .B2(G142), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n884), .B(new_n889), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n883), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n883), .A2(new_n890), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XOR2_X1   g468(.A(G160), .B(KEYINPUT110), .Z(new_n894));
  XNOR2_X1  g469(.A(G162), .B(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(new_n623), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n896), .B1(new_n891), .B2(new_n892), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n879), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g476(.A1(new_n526), .A2(G91), .ZN(new_n902));
  INV_X1    g477(.A(new_n571), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n569), .A2(new_n570), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n902), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n574), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n604), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n572), .A2(new_n611), .A3(new_n574), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(KEYINPUT112), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT112), .ZN(new_n910));
  NAND3_X1  g485(.A1(G299), .A2(new_n910), .A3(new_n604), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n909), .A2(KEYINPUT41), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT41), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n907), .A2(new_n913), .A3(new_n908), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n611), .A2(G559), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n858), .A2(new_n916), .A3(new_n861), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n916), .B1(new_n858), .B2(new_n861), .ZN(new_n919));
  OR3_X1    g494(.A1(new_n915), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n909), .A2(new_n911), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n922), .B1(new_n918), .B2(new_n919), .ZN(new_n923));
  AOI21_X1  g498(.A(KEYINPUT113), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(G303), .A2(G290), .ZN(new_n925));
  NAND2_X1  g500(.A1(G166), .A2(new_n835), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n812), .A2(G305), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n811), .A2(new_n798), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n925), .A2(new_n926), .A3(new_n928), .A4(new_n929), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n933), .B(KEYINPUT42), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n920), .A2(KEYINPUT113), .A3(new_n923), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n924), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n924), .B1(new_n935), .B2(new_n934), .ZN(new_n937));
  OAI21_X1  g512(.A(G868), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n938), .B1(G868), .B2(new_n855), .ZN(G295));
  OAI21_X1  g514(.A(new_n938), .B1(G868), .B2(new_n855), .ZN(G331));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n858), .A2(new_n861), .ZN(new_n942));
  NAND2_X1  g517(.A1(G301), .A2(new_n540), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n943), .B1(G286), .B2(G301), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n858), .A2(new_n861), .A3(new_n944), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n915), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n858), .A2(new_n861), .A3(new_n944), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n944), .B1(new_n858), .B2(new_n861), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n921), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n933), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n907), .A2(new_n908), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n946), .A2(KEYINPUT41), .A3(new_n955), .A4(new_n947), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n949), .A2(new_n950), .A3(new_n913), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n933), .B(new_n956), .C1(new_n957), .C2(new_n922), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT43), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n954), .A2(new_n958), .A3(new_n959), .A4(new_n879), .ZN(new_n960));
  AOI21_X1  g535(.A(G37), .B1(new_n952), .B2(new_n953), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n933), .A2(new_n948), .A3(new_n951), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT114), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n960), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  AOI211_X1 g540(.A(KEYINPUT114), .B(new_n959), .C1(new_n961), .C2(new_n962), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n941), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n954), .A2(new_n958), .A3(new_n879), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n941), .B1(new_n968), .B2(KEYINPUT43), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT115), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n961), .A2(new_n959), .A3(new_n962), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n970), .B1(new_n969), .B2(new_n971), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n967), .B1(new_n972), .B2(new_n973), .ZN(G397));
  XOR2_X1   g549(.A(KEYINPUT116), .B(G1384), .Z(new_n975));
  NAND2_X1  g550(.A1(new_n508), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT45), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G40), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n468), .A2(new_n471), .A3(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G1996), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n880), .B(new_n983), .ZN(new_n984));
  OR2_X1    g559(.A1(new_n829), .A2(new_n831), .ZN(new_n985));
  INV_X1    g560(.A(G2067), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n779), .B(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n829), .A2(new_n831), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n984), .A2(new_n985), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  XNOR2_X1  g564(.A(G290), .B(G1986), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n982), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G1384), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n993), .B1(KEYINPUT69), .B2(new_n492), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n502), .A2(new_n506), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n487), .A2(G126), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n498), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n992), .B(new_n980), .C1(new_n994), .C2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G8), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n808), .A2(G1976), .A3(new_n810), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT52), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n587), .A2(G651), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n582), .A2(new_n583), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(G1981), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(G305), .B2(G1981), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT49), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1007), .B(KEYINPUT49), .C1(G305), .C2(G1981), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1010), .A2(new_n1001), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1976), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT52), .B1(G288), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1001), .A2(new_n1002), .A3(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1004), .A2(new_n1012), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT120), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1004), .A2(new_n1012), .A3(KEYINPUT120), .A4(new_n1015), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n992), .B1(new_n994), .B2(new_n997), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n981), .B1(new_n1021), .B2(new_n977), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n508), .A2(KEYINPUT45), .A3(new_n975), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n805), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT119), .ZN(new_n1026));
  XOR2_X1   g601(.A(KEYINPUT117), .B(KEYINPUT50), .Z(new_n1027));
  AOI21_X1  g602(.A(new_n1027), .B1(new_n508), .B2(new_n992), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1026), .B1(new_n1028), .B2(new_n981), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n498), .A2(new_n995), .A3(new_n996), .ZN(new_n1030));
  AOI21_X1  g605(.A(G1384), .B1(new_n1030), .B2(new_n496), .ZN(new_n1031));
  OAI211_X1 g606(.A(KEYINPUT119), .B(new_n980), .C1(new_n1031), .C2(new_n1027), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1021), .A2(KEYINPUT50), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1029), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1025), .B1(new_n1035), .B2(G2090), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(G8), .ZN(new_n1037));
  XNOR2_X1  g612(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n529), .A2(G8), .A3(new_n531), .A4(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n529), .A2(G8), .A3(new_n531), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1038), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1037), .A2(new_n1039), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1021), .A2(KEYINPUT50), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n992), .B(new_n1027), .C1(new_n994), .C2(new_n997), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1044), .A2(new_n980), .A3(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1025), .B1(G2090), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1042), .A2(new_n1039), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1047), .A2(new_n1048), .A3(G8), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1020), .A2(new_n1043), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1045), .A2(new_n980), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT50), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1054), .B1(new_n508), .B2(new_n992), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT122), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G1961), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT122), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1044), .A2(new_n1058), .A3(new_n980), .A4(new_n1045), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1056), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1061), .B1(new_n1024), .B2(G2078), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1031), .A2(KEYINPUT45), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1061), .A2(G2078), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1022), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1060), .A2(new_n1062), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(G171), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n978), .A2(new_n980), .A3(new_n1023), .A4(new_n1064), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1060), .A2(new_n1062), .A3(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1067), .B1(new_n1069), .B2(G171), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1069), .A2(G171), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1073), .B(KEYINPUT54), .C1(G171), .C2(new_n1066), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1022), .A2(new_n1063), .ZN(new_n1075));
  INV_X1    g650(.A(G1966), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G2084), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1044), .A2(new_n1078), .A3(new_n980), .A4(new_n1045), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1077), .A2(G168), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(G8), .ZN(new_n1081));
  AOI21_X1  g656(.A(G168), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT51), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT51), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1080), .A2(new_n1084), .A3(G8), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1052), .A2(new_n1072), .A3(new_n1074), .A4(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1056), .A2(new_n733), .A3(new_n1059), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n999), .A2(new_n986), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT60), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT127), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1092), .A2(new_n1093), .A3(new_n604), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT60), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1096));
  OAI21_X1  g671(.A(KEYINPUT127), .B1(new_n1096), .B2(new_n611), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1094), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1095), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1021), .A2(new_n977), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1102), .A2(new_n983), .A3(new_n980), .A4(new_n1023), .ZN(new_n1103));
  XOR2_X1   g678(.A(KEYINPUT58), .B(G1341), .Z(new_n1104));
  NAND2_X1  g679(.A1(new_n998), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(KEYINPUT124), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT124), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n998), .A2(new_n1107), .A3(new_n1104), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1103), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT125), .ZN(new_n1110));
  AND3_X1   g685(.A1(new_n1109), .A2(new_n1110), .A3(new_n557), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1110), .B1(new_n1109), .B2(new_n557), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1101), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1109), .A2(new_n557), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT125), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1109), .A2(new_n1110), .A3(new_n557), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1115), .A2(KEYINPUT59), .A3(new_n1116), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1113), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT57), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n572), .A2(new_n1120), .A3(new_n574), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1027), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n981), .B1(new_n1021), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1033), .B1(new_n1124), .B2(KEYINPUT119), .ZN(new_n1125));
  AOI21_X1  g700(.A(G1956), .B1(new_n1125), .B2(new_n1029), .ZN(new_n1126));
  XNOR2_X1  g701(.A(KEYINPUT56), .B(G2072), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1022), .A2(new_n1023), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1122), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1035), .A2(new_n763), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1122), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1131), .A2(new_n1132), .A3(new_n1128), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT61), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1130), .A2(new_n1133), .A3(KEYINPUT61), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1118), .A2(KEYINPUT126), .A3(new_n1135), .A4(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT126), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1136), .A2(new_n1113), .A3(new_n1117), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1138), .B1(new_n1139), .B2(new_n1134), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1100), .A2(new_n1137), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1130), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n611), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1133), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1144), .B(KEYINPUT123), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1087), .B1(new_n1141), .B2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(G305), .A2(G1981), .ZN(new_n1147));
  NOR2_X1   g722(.A1(G288), .A2(G1976), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1147), .B1(new_n1012), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1001), .ZN(new_n1150));
  OAI22_X1  g725(.A1(new_n1050), .A2(new_n1016), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1048), .B1(new_n1047), .B2(G8), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1049), .A2(new_n1152), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n1154), .A2(new_n1000), .A3(G286), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT63), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1016), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1153), .A2(new_n1155), .A3(new_n1157), .ZN(new_n1158));
  XOR2_X1   g733(.A(KEYINPUT121), .B(KEYINPUT63), .Z(new_n1159));
  AOI21_X1  g734(.A(new_n1151), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1155), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1161), .B1(new_n1153), .B2(new_n1157), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1067), .B1(new_n1086), .B2(KEYINPUT62), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT62), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1083), .A2(new_n1164), .A3(new_n1085), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1162), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1160), .B1(new_n1166), .B2(new_n1051), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n991), .B1(new_n1146), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(G1986), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n982), .A2(new_n1169), .A3(new_n835), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT48), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  AND2_X1   g747(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1173));
  AOI211_X1 g748(.A(new_n1172), .B(new_n1173), .C1(new_n982), .C2(new_n989), .ZN(new_n1174));
  INV_X1    g749(.A(new_n987), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n982), .B1(new_n1175), .B2(new_n880), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n982), .A2(new_n983), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1177), .B(KEYINPUT46), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  XOR2_X1   g754(.A(new_n1179), .B(KEYINPUT47), .Z(new_n1180));
  NAND2_X1  g755(.A1(new_n984), .A2(new_n987), .ZN(new_n1181));
  OAI22_X1  g756(.A1(new_n1181), .A2(new_n988), .B1(G2067), .B2(new_n779), .ZN(new_n1182));
  AOI211_X1 g757(.A(new_n1174), .B(new_n1180), .C1(new_n982), .C2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1168), .A2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g759(.A1(G401), .A2(new_n461), .ZN(new_n1186));
  NAND2_X1  g760(.A1(new_n690), .A2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g761(.A1(new_n1187), .A2(G227), .ZN(new_n1188));
  OAI211_X1 g762(.A(new_n1188), .B(new_n900), .C1(new_n965), .C2(new_n966), .ZN(G225));
  INV_X1    g763(.A(G225), .ZN(G308));
endmodule


