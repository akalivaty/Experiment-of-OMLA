//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 1 0 0 0 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 1 0 0 1 0 1 1 1 1 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n746, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n859, new_n860, new_n861, new_n862, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984, new_n985, new_n986;
  XOR2_X1   g000(.A(G8gat), .B(G36gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G64gat), .ZN(new_n203));
  INV_X1    g002(.A(G92gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G226gat), .A2(G233gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208));
  INV_X1    g007(.A(G169gat), .ZN(new_n209));
  INV_X1    g008(.A(G176gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  OR2_X1    g010(.A1(new_n211), .A2(KEYINPUT26), .ZN(new_n212));
  NAND2_X1  g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(KEYINPUT26), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(KEYINPUT27), .B(G183gat), .ZN(new_n216));
  INV_X1    g015(.A(G190gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(KEYINPUT28), .A3(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT69), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n218), .B(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT67), .ZN(new_n221));
  INV_X1    g020(.A(G183gat), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT27), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT27), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n224), .A2(KEYINPUT67), .A3(G183gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n223), .A2(new_n217), .A3(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT68), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT28), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n223), .A2(KEYINPUT68), .A3(new_n217), .A4(new_n225), .ZN(new_n230));
  AND3_X1   g029(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n208), .B(new_n215), .C1(new_n220), .C2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT24), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n208), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n222), .A2(new_n217), .ZN(new_n237));
  NAND3_X1  g036(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n238));
  AND2_X1   g037(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n236), .B(new_n237), .C1(new_n239), .C2(new_n235), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n213), .A2(KEYINPUT23), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(new_n211), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n209), .A2(new_n210), .A3(KEYINPUT23), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n240), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT64), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n239), .A2(new_n245), .A3(new_n237), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n234), .A2(new_n238), .A3(new_n237), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT64), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT25), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  XOR2_X1   g048(.A(KEYINPUT65), .B(G169gat), .Z(new_n250));
  AND2_X1   g049(.A1(new_n210), .A2(KEYINPUT23), .ZN(new_n251));
  AOI22_X1  g050(.A1(new_n250), .A2(new_n251), .B1(new_n211), .B2(new_n241), .ZN(new_n252));
  AOI22_X1  g051(.A1(new_n244), .A2(KEYINPUT25), .B1(new_n249), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT73), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n232), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n254), .B1(new_n232), .B2(new_n253), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n207), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n232), .A2(new_n253), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n207), .A2(KEYINPUT29), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G197gat), .B(G204gat), .ZN(new_n262));
  INV_X1    g061(.A(G211gat), .ZN(new_n263));
  INV_X1    g062(.A(G218gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n262), .B1(KEYINPUT22), .B2(new_n265), .ZN(new_n266));
  XOR2_X1   g065(.A(G211gat), .B(G218gat), .Z(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n261), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n258), .A2(KEYINPUT73), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n232), .A2(new_n253), .A3(new_n254), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n271), .A2(new_n272), .A3(new_n259), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n232), .A2(new_n253), .A3(new_n207), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n273), .A2(new_n268), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n205), .B1(new_n270), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT74), .B1(new_n276), .B2(KEYINPUT30), .ZN(new_n277));
  INV_X1    g076(.A(new_n205), .ZN(new_n278));
  INV_X1    g077(.A(new_n275), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n268), .B1(new_n257), .B2(new_n260), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT74), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT30), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n276), .A2(KEYINPUT30), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n270), .A2(new_n275), .A3(new_n205), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n277), .A2(new_n284), .A3(new_n285), .A4(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G155gat), .A2(G162gat), .ZN(new_n288));
  INV_X1    g087(.A(G155gat), .ZN(new_n289));
  INV_X1    g088(.A(G162gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n288), .B1(new_n291), .B2(KEYINPUT2), .ZN(new_n292));
  XOR2_X1   g091(.A(G141gat), .B(G148gat), .Z(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT75), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT75), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n292), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n291), .A2(new_n288), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT2), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n299), .B1(new_n293), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT3), .ZN(new_n304));
  INV_X1    g103(.A(G113gat), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT70), .B1(new_n305), .B2(G120gat), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT70), .ZN(new_n307));
  INV_X1    g106(.A(G120gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(new_n308), .A3(G113gat), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n306), .B(new_n309), .C1(G113gat), .C2(new_n308), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT1), .ZN(new_n311));
  XNOR2_X1  g110(.A(G127gat), .B(G134gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n312), .ZN(new_n314));
  XNOR2_X1  g113(.A(G113gat), .B(G120gat), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n314), .B1(KEYINPUT1), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n301), .B1(new_n295), .B2(new_n297), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT3), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n317), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT4), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n317), .A2(KEYINPUT71), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT71), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n313), .A2(new_n324), .A3(new_n316), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n322), .B1(new_n326), .B2(new_n303), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n318), .A2(KEYINPUT4), .A3(new_n316), .A4(new_n313), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n321), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G225gat), .A2(G233gat), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n303), .B(new_n317), .ZN(new_n333));
  OR2_X1    g132(.A1(new_n333), .A2(new_n331), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n332), .A2(KEYINPUT39), .A3(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(KEYINPUT0), .B(G57gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n336), .B(G85gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(G1gat), .B(G29gat), .ZN(new_n338));
  XOR2_X1   g137(.A(new_n337), .B(new_n338), .Z(new_n339));
  OAI21_X1  g138(.A(new_n339), .B1(new_n332), .B2(KEYINPUT39), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT40), .ZN(new_n341));
  NOR3_X1   g140(.A1(new_n335), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n318), .A2(new_n319), .ZN(new_n343));
  AOI211_X1 g142(.A(KEYINPUT3), .B(new_n301), .C1(new_n295), .C2(new_n297), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n331), .B1(new_n345), .B2(new_n317), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT76), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n322), .B1(new_n303), .B2(new_n317), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n323), .A2(new_n318), .A3(KEYINPUT4), .A4(new_n325), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n346), .A2(new_n347), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n321), .A2(new_n330), .A3(new_n348), .A4(new_n349), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT76), .ZN(new_n352));
  XOR2_X1   g151(.A(KEYINPUT77), .B(KEYINPUT5), .Z(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n354), .B1(new_n333), .B2(new_n331), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n350), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n321), .A2(new_n327), .A3(new_n328), .A4(new_n330), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT78), .B1(new_n357), .B2(new_n353), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n321), .A2(new_n327), .A3(new_n328), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT78), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n359), .A2(new_n360), .A3(new_n354), .A4(new_n330), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n356), .A2(new_n358), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n339), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT83), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n362), .A2(KEYINPUT83), .A3(new_n363), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n342), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n341), .B1(new_n335), .B2(new_n340), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n287), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT84), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AND2_X1   g171(.A1(G228gat), .A2(G233gat), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n269), .B1(new_n344), .B2(KEYINPUT29), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT29), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n268), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n318), .B1(new_n377), .B2(new_n319), .ZN(new_n378));
  OAI211_X1 g177(.A(KEYINPUT81), .B(new_n373), .C1(new_n375), .C2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n378), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n373), .A2(KEYINPUT81), .ZN(new_n381));
  OR2_X1    g180(.A1(new_n373), .A2(KEYINPUT81), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n380), .A2(new_n381), .A3(new_n382), .A4(new_n374), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n379), .A2(new_n383), .A3(G22gat), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT82), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G78gat), .B(G106gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT31), .B(G50gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n387), .B(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n379), .A2(new_n383), .ZN(new_n391));
  INV_X1    g190(.A(G22gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(new_n384), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n386), .A2(new_n389), .B1(new_n393), .B2(new_n384), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n366), .A2(new_n367), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n356), .A2(new_n339), .A3(new_n358), .A4(new_n361), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT6), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n364), .A2(new_n401), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT37), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n407), .B1(new_n279), .B2(new_n280), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n270), .A2(KEYINPUT37), .A3(new_n275), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(new_n409), .A3(new_n205), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n276), .B1(new_n410), .B2(KEYINPUT38), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n257), .A2(new_n268), .A3(new_n260), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n273), .A2(new_n274), .ZN(new_n413));
  OAI211_X1 g212(.A(KEYINPUT37), .B(new_n412), .C1(new_n413), .C2(new_n268), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT38), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n408), .A2(new_n414), .A3(new_n415), .A4(new_n205), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n404), .A2(new_n406), .A3(new_n411), .A4(new_n416), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n287), .A2(new_n368), .A3(KEYINPUT84), .A4(new_n369), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n372), .A2(new_n398), .A3(new_n417), .A4(new_n418), .ZN(new_n419));
  XOR2_X1   g218(.A(G15gat), .B(G43gat), .Z(new_n420));
  XNOR2_X1  g219(.A(G71gat), .B(G99gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n420), .B(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(G227gat), .ZN(new_n423));
  INV_X1    g222(.A(G233gat), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n258), .A2(new_n326), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n232), .A2(new_n253), .A3(new_n323), .A4(new_n325), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n422), .B1(new_n429), .B2(KEYINPUT33), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT32), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  OR2_X1    g231(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n427), .A2(new_n426), .A3(new_n428), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n434), .B(KEYINPUT34), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n427), .A2(new_n428), .ZN(new_n437));
  AOI221_X4 g236(.A(new_n431), .B1(KEYINPUT33), .B2(new_n422), .C1(new_n437), .C2(new_n425), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n433), .A2(new_n436), .A3(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n430), .A2(new_n432), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n435), .B1(new_n441), .B2(new_n438), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT36), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n440), .A2(new_n442), .A3(KEYINPUT72), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT72), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n445), .B(new_n435), .C1(new_n441), .C2(new_n438), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n443), .B1(new_n447), .B2(KEYINPUT36), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT79), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n402), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n364), .A2(KEYINPUT80), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n400), .A2(KEYINPUT79), .A3(new_n401), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT80), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n362), .A2(new_n453), .A3(new_n363), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n450), .A2(new_n451), .A3(new_n452), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n406), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n285), .A2(new_n286), .ZN(new_n457));
  NOR3_X1   g256(.A1(new_n276), .A2(KEYINPUT74), .A3(KEYINPUT30), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n282), .B1(new_n281), .B2(new_n283), .ZN(new_n459));
  NOR3_X1   g258(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n448), .B1(new_n461), .B2(new_n397), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n419), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n440), .A2(new_n442), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n464), .A2(new_n397), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n402), .B1(new_n366), .B2(new_n367), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n460), .B(new_n465), .C1(new_n405), .C2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT35), .ZN(new_n468));
  AOI211_X1 g267(.A(new_n468), .B(new_n397), .C1(new_n444), .C2(new_n446), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n287), .B1(new_n455), .B2(new_n406), .ZN(new_n470));
  AOI22_X1  g269(.A1(new_n467), .A2(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n463), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(G15gat), .B(G22gat), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT16), .ZN(new_n474));
  OR2_X1    g273(.A1(new_n474), .A2(G1gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n476), .B1(G1gat), .B2(new_n473), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(G8gat), .ZN(new_n478));
  INV_X1    g277(.A(G8gat), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n476), .B(new_n479), .C1(G1gat), .C2(new_n473), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  XOR2_X1   g280(.A(G57gat), .B(G64gat), .Z(new_n482));
  OR2_X1    g281(.A1(G71gat), .A2(G78gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(G71gat), .A2(G78gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT9), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n482), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(G57gat), .B(G64gat), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n484), .B(new_n483), .C1(new_n489), .C2(new_n486), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n481), .B1(KEYINPUT21), .B2(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n492), .B(G183gat), .ZN(new_n493));
  XOR2_X1   g292(.A(KEYINPUT91), .B(KEYINPUT21), .Z(new_n494));
  NOR2_X1   g293(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n493), .B(new_n495), .ZN(new_n496));
  XOR2_X1   g295(.A(G127gat), .B(G155gat), .Z(new_n497));
  XNOR2_X1  g296(.A(new_n497), .B(KEYINPUT20), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n496), .A2(new_n498), .ZN(new_n500));
  XNOR2_X1  g299(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n501), .B(G211gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(G231gat), .A2(G233gat), .ZN(new_n503));
  XOR2_X1   g302(.A(new_n502), .B(new_n503), .Z(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  OR3_X1    g304(.A1(new_n499), .A2(new_n500), .A3(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n505), .B1(new_n499), .B2(new_n500), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT95), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT17), .ZN(new_n510));
  INV_X1    g309(.A(G50gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(G43gat), .ZN(new_n512));
  INV_X1    g311(.A(G43gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(G50gat), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT86), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n512), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n515), .B1(new_n512), .B2(new_n514), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT14), .ZN(new_n519));
  INV_X1    g318(.A(G29gat), .ZN(new_n520));
  INV_X1    g319(.A(G36gat), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(KEYINPUT87), .A3(new_n523), .ZN(new_n524));
  NOR3_X1   g323(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT87), .ZN(new_n526));
  AOI22_X1  g325(.A1(new_n525), .A2(new_n526), .B1(G29gat), .B2(G36gat), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n518), .A2(KEYINPUT15), .A3(new_n524), .A4(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n514), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(KEYINPUT86), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n512), .A2(new_n514), .A3(new_n515), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n530), .A2(KEYINPUT15), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n522), .A2(new_n523), .ZN(new_n533));
  NAND2_X1  g332(.A1(G29gat), .A2(G36gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(G43gat), .B(G50gat), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n533), .B(new_n534), .C1(KEYINPUT15), .C2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n510), .B1(new_n528), .B2(new_n537), .ZN(new_n538));
  AND3_X1   g337(.A1(KEYINPUT93), .A2(G85gat), .A3(G92gat), .ZN(new_n539));
  OR2_X1    g338(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n540));
  NAND2_X1  g339(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(KEYINPUT93), .A2(G85gat), .A3(G92gat), .ZN(new_n543));
  AND2_X1   g342(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n544));
  NOR2_X1   g343(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(G99gat), .A2(G106gat), .ZN(new_n547));
  INV_X1    g346(.A(G85gat), .ZN(new_n548));
  AOI22_X1  g347(.A1(KEYINPUT8), .A2(new_n547), .B1(new_n548), .B2(new_n204), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n542), .A2(new_n546), .A3(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(G99gat), .B(G106gat), .Z(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n542), .A2(new_n551), .A3(new_n546), .A4(new_n549), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n528), .A2(new_n510), .A3(new_n537), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT88), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n528), .A2(new_n537), .A3(KEYINPUT88), .A4(new_n510), .ZN(new_n559));
  AOI211_X1 g358(.A(new_n538), .B(new_n555), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(G190gat), .B(G218gat), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  AND2_X1   g361(.A1(G232gat), .A2(G233gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT41), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n528), .A2(new_n537), .ZN(new_n565));
  INV_X1    g364(.A(new_n555), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NOR3_X1   g366(.A1(new_n560), .A2(new_n562), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n558), .A2(new_n559), .ZN(new_n569));
  INV_X1    g368(.A(new_n538), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n569), .A2(new_n570), .A3(new_n566), .ZN(new_n571));
  INV_X1    g370(.A(new_n567), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n561), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n509), .B1(new_n568), .B2(new_n573), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n562), .B1(new_n560), .B2(new_n567), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n571), .A2(new_n561), .A3(new_n572), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n575), .A2(KEYINPUT95), .A3(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n563), .A2(KEYINPUT41), .ZN(new_n578));
  XNOR2_X1  g377(.A(G134gat), .B(G162gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n574), .A2(new_n577), .A3(new_n581), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n575), .A2(KEYINPUT95), .A3(new_n576), .A4(new_n580), .ZN(new_n583));
  AND2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n508), .A2(new_n584), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n472), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n538), .A2(new_n481), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n569), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n481), .A2(new_n528), .A3(new_n537), .ZN(new_n589));
  NAND2_X1  g388(.A1(G229gat), .A2(G233gat), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT18), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(KEYINPUT89), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n478), .A2(new_n480), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n595), .A2(new_n565), .ZN(new_n596));
  INV_X1    g395(.A(new_n590), .ZN(new_n597));
  AOI211_X1 g396(.A(new_n596), .B(new_n597), .C1(new_n569), .C2(new_n587), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n595), .A2(new_n565), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(new_n589), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n590), .B(KEYINPUT13), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  AOI22_X1  g401(.A1(new_n598), .A2(KEYINPUT18), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT89), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n591), .A2(new_n604), .A3(new_n592), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n594), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(KEYINPUT11), .B(G169gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(G197gat), .ZN(new_n608));
  XOR2_X1   g407(.A(G113gat), .B(G141gat), .Z(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n610), .A2(KEYINPUT85), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(KEYINPUT85), .ZN(new_n612));
  AND3_X1   g411(.A1(new_n611), .A2(KEYINPUT12), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT12), .B1(new_n611), .B2(new_n612), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n606), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT90), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n593), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n591), .A2(KEYINPUT90), .A3(new_n592), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n619), .A2(new_n603), .A3(new_n615), .A4(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(G230gat), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n624), .A2(new_n424), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n550), .A2(KEYINPUT96), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n627), .A2(new_n490), .A3(new_n488), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(new_n555), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n491), .A2(new_n553), .A3(new_n554), .A4(new_n627), .ZN(new_n630));
  AOI21_X1  g429(.A(KEYINPUT10), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n555), .A2(KEYINPUT10), .A3(new_n491), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n626), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n629), .A2(new_n630), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n634), .B1(new_n626), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT97), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G120gat), .B(G148gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(new_n210), .ZN(new_n640));
  INV_X1    g439(.A(G204gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n636), .A2(new_n637), .A3(new_n642), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n623), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n586), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n648), .A2(new_n456), .ZN(new_n649));
  XOR2_X1   g448(.A(KEYINPUT98), .B(G1gat), .Z(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(G1324gat));
  OAI21_X1  g450(.A(G8gat), .B1(new_n648), .B2(new_n460), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT99), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n648), .A2(new_n460), .ZN(new_n655));
  NAND2_X1  g454(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n474), .A2(new_n479), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n658), .A2(KEYINPUT42), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(KEYINPUT42), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n654), .B1(new_n659), .B2(new_n660), .ZN(G1325gat));
  INV_X1    g460(.A(G15gat), .ZN(new_n662));
  INV_X1    g461(.A(new_n448), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n648), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n464), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n586), .A2(new_n647), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n664), .B1(new_n662), .B2(new_n666), .ZN(G1326gat));
  NOR2_X1   g466(.A1(new_n648), .A2(new_n398), .ZN(new_n668));
  XOR2_X1   g467(.A(KEYINPUT43), .B(G22gat), .Z(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(G1327gat));
  INV_X1    g469(.A(new_n647), .ZN(new_n671));
  AND3_X1   g470(.A1(new_n506), .A2(new_n507), .A3(KEYINPUT101), .ZN(new_n672));
  AOI21_X1  g471(.A(KEYINPUT101), .B1(new_n506), .B2(new_n507), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n467), .A2(new_n468), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n469), .A2(new_n470), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n678), .B1(new_n462), .B2(new_n419), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n582), .A2(new_n583), .ZN(new_n680));
  OAI21_X1  g479(.A(KEYINPUT44), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n680), .B1(new_n463), .B2(new_n471), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AOI211_X1 g483(.A(new_n671), .B(new_n675), .C1(new_n681), .C2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n456), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n685), .A2(KEYINPUT102), .A3(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT102), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n682), .A2(new_n683), .ZN(new_n689));
  AOI211_X1 g488(.A(KEYINPUT44), .B(new_n680), .C1(new_n463), .C2(new_n471), .ZN(new_n690));
  OAI211_X1 g489(.A(new_n647), .B(new_n674), .C1(new_n689), .C2(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n688), .B1(new_n691), .B2(new_n456), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n687), .A2(G29gat), .A3(new_n692), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n682), .A2(new_n686), .A3(new_n647), .A4(new_n508), .ZN(new_n694));
  OR3_X1    g493(.A1(new_n694), .A2(KEYINPUT100), .A3(G29gat), .ZN(new_n695));
  OAI21_X1  g494(.A(KEYINPUT100), .B1(new_n694), .B2(G29gat), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n695), .A2(KEYINPUT45), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n696), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT45), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n693), .A2(new_n697), .A3(new_n700), .ZN(G1328gat));
  NAND3_X1  g500(.A1(new_n682), .A2(new_n647), .A3(new_n508), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n702), .A2(G36gat), .A3(new_n460), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT46), .ZN(new_n704));
  OAI21_X1  g503(.A(G36gat), .B1(new_n691), .B2(new_n460), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(G1329gat));
  OAI21_X1  g505(.A(G43gat), .B1(new_n691), .B2(new_n663), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT47), .ZN(new_n708));
  OR3_X1    g507(.A1(new_n702), .A2(G43gat), .A3(new_n464), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n708), .B1(new_n707), .B2(new_n709), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(G1330gat));
  INV_X1    g511(.A(KEYINPUT104), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n713), .B1(new_n691), .B2(new_n398), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n671), .B1(new_n681), .B2(new_n684), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n715), .A2(KEYINPUT104), .A3(new_n397), .A4(new_n674), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n714), .A2(new_n716), .A3(G50gat), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT48), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT103), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n682), .A2(new_n719), .A3(new_n647), .A4(new_n508), .ZN(new_n720));
  AND3_X1   g519(.A1(new_n720), .A2(new_n511), .A3(new_n397), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n702), .A2(KEYINPUT103), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n718), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n717), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n511), .B1(new_n685), .B2(new_n397), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n721), .A2(new_n722), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n718), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n724), .A2(new_n727), .ZN(G1331gat));
  INV_X1    g527(.A(new_n646), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n622), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n586), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n686), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g533(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n586), .A2(new_n287), .A3(new_n730), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT105), .ZN(new_n737));
  OR2_X1    g536(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(G1333gat));
  INV_X1    g538(.A(G71gat), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n732), .A2(new_n740), .A3(new_n665), .ZN(new_n741));
  OAI21_X1  g540(.A(G71gat), .B1(new_n731), .B2(new_n663), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT50), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(G1334gat));
  NOR2_X1   g544(.A1(new_n731), .A2(new_n398), .ZN(new_n746));
  XNOR2_X1  g545(.A(KEYINPUT106), .B(G78gat), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(G1335gat));
  NAND2_X1  g547(.A1(new_n508), .A2(new_n623), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT107), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n682), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT51), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n682), .A2(KEYINPUT51), .A3(new_n751), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n729), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(G85gat), .B1(new_n756), .B2(new_n686), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n681), .A2(new_n684), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n750), .A2(new_n729), .ZN(new_n759));
  AND3_X1   g558(.A1(new_n758), .A2(G85gat), .A3(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n757), .B1(new_n686), .B2(new_n760), .ZN(G1336gat));
  NAND3_X1  g560(.A1(new_n756), .A2(new_n204), .A3(new_n287), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n758), .A2(new_n287), .A3(new_n759), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G92gat), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(KEYINPUT52), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n762), .A2(new_n764), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n768), .ZN(G1337gat));
  INV_X1    g568(.A(G99gat), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n756), .A2(new_n770), .A3(new_n665), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n758), .A2(new_n448), .A3(new_n759), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(G99gat), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(KEYINPUT108), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT108), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n771), .A2(new_n773), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(G1338gat));
  NAND2_X1  g577(.A1(new_n756), .A2(new_n397), .ZN(new_n779));
  INV_X1    g578(.A(G106gat), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n758), .A2(G106gat), .A3(new_n397), .A4(new_n759), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n781), .A2(KEYINPUT53), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n784));
  AOI21_X1  g583(.A(G106gat), .B1(new_n756), .B2(new_n397), .ZN(new_n785));
  INV_X1    g584(.A(new_n782), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n783), .A2(new_n787), .ZN(G1339gat));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT10), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n628), .A2(new_n555), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n491), .A2(new_n627), .B1(new_n553), .B2(new_n554), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n793), .A2(new_n625), .A3(new_n632), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n794), .A2(new_n634), .A3(KEYINPUT54), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n625), .B1(new_n793), .B2(new_n632), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n795), .A2(new_n798), .A3(new_n642), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n795), .A2(new_n798), .A3(KEYINPUT55), .A4(new_n642), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n635), .A2(new_n626), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n796), .A2(new_n803), .A3(new_n642), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n801), .A2(new_n802), .A3(new_n805), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n598), .A2(new_n618), .A3(KEYINPUT18), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT90), .B1(new_n591), .B2(new_n592), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n596), .B1(new_n569), .B2(new_n587), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n810), .A2(KEYINPUT18), .A3(new_n590), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n600), .A2(new_n602), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n615), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  AOI211_X1 g613(.A(new_n481), .B(new_n538), .C1(new_n558), .C2(new_n559), .ZN(new_n815));
  OAI211_X1 g614(.A(KEYINPUT109), .B(new_n597), .C1(new_n815), .C2(new_n596), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT109), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n817), .B1(new_n810), .B2(new_n590), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n599), .A2(new_n589), .A3(new_n601), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n819), .B(KEYINPUT110), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n816), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  AOI22_X1  g620(.A1(new_n809), .A2(new_n814), .B1(new_n610), .B2(new_n821), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n584), .A2(new_n789), .A3(new_n806), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n610), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n804), .B1(new_n799), .B2(new_n800), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n621), .A2(new_n802), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(KEYINPUT111), .B1(new_n826), .B2(new_n680), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n823), .A2(new_n827), .ZN(new_n828));
  AOI211_X1 g627(.A(KEYINPUT89), .B(KEYINPUT18), .C1(new_n810), .C2(new_n590), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n604), .B1(new_n591), .B2(new_n592), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n615), .B1(new_n831), .B2(new_n603), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n813), .A2(new_n807), .A3(new_n808), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n806), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n822), .A2(new_n646), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n584), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT112), .B1(new_n828), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n825), .A2(new_n802), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n838), .B1(new_n617), .B2(new_n621), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n621), .A2(new_n646), .A3(new_n824), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n680), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT112), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n841), .A2(new_n842), .A3(new_n827), .A4(new_n823), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n837), .A2(new_n674), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n585), .A2(new_n623), .A3(new_n729), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n456), .A2(new_n287), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n447), .A2(new_n398), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n851), .A2(new_n305), .A3(new_n622), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n848), .A2(new_n465), .ZN(new_n853));
  OAI21_X1  g652(.A(G113gat), .B1(new_n853), .B2(new_n623), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(new_n854), .ZN(G1340gat));
  NAND3_X1  g654(.A1(new_n851), .A2(new_n308), .A3(new_n646), .ZN(new_n856));
  OAI21_X1  g655(.A(G120gat), .B1(new_n853), .B2(new_n729), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(G1341gat));
  INV_X1    g657(.A(new_n508), .ZN(new_n859));
  AOI21_X1  g658(.A(G127gat), .B1(new_n851), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(G127gat), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n853), .A2(new_n861), .A3(new_n674), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n860), .A2(new_n862), .ZN(G1342gat));
  INV_X1    g662(.A(G134gat), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n851), .A2(new_n864), .A3(new_n584), .ZN(new_n865));
  XOR2_X1   g664(.A(new_n865), .B(KEYINPUT56), .Z(new_n866));
  OAI21_X1  g665(.A(G134gat), .B1(new_n853), .B2(new_n680), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(G1343gat));
  NAND2_X1  g667(.A1(new_n846), .A2(new_n397), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n869), .A2(KEYINPUT113), .A3(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT113), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n398), .B1(new_n844), .B2(new_n845), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n872), .B1(new_n873), .B2(KEYINPUT57), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n799), .A2(KEYINPUT114), .A3(new_n800), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n800), .A2(KEYINPUT114), .ZN(new_n876));
  OR2_X1    g675(.A1(new_n799), .A2(new_n876), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n622), .A2(new_n805), .A3(new_n875), .A4(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n584), .B1(new_n878), .B2(new_n835), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n879), .A2(new_n828), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n845), .B1(new_n880), .B2(new_n859), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(KEYINPUT57), .A3(new_n397), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n871), .A2(new_n874), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n663), .A2(new_n847), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n883), .A2(new_n622), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(G141gat), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT115), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(G141gat), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n448), .A2(new_n398), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n848), .A2(new_n890), .A3(new_n622), .A4(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n887), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n889), .A2(new_n893), .A3(KEYINPUT58), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT58), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n887), .B(new_n892), .C1(new_n888), .C2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(new_n896), .ZN(G1344gat));
  NAND3_X1  g696(.A1(new_n873), .A2(KEYINPUT118), .A3(KEYINPUT57), .ZN(new_n898));
  AOI211_X1 g697(.A(new_n870), .B(new_n398), .C1(new_n844), .C2(new_n845), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT118), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n826), .A2(new_n680), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n508), .B1(new_n879), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n398), .B1(new_n902), .B2(new_n845), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n900), .B1(new_n903), .B2(KEYINPUT57), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n898), .B(new_n646), .C1(new_n899), .C2(new_n904), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n884), .A2(KEYINPUT117), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n884), .A2(KEYINPUT117), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(G148gat), .ZN(new_n909));
  OAI21_X1  g708(.A(KEYINPUT59), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n883), .A2(new_n646), .A3(new_n885), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n909), .A2(KEYINPUT59), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n911), .A2(KEYINPUT116), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(KEYINPUT116), .B1(new_n911), .B2(new_n912), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n910), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n848), .A2(new_n891), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n917), .A2(new_n909), .A3(new_n646), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n915), .A2(new_n918), .ZN(G1345gat));
  AOI21_X1  g718(.A(G155gat), .B1(new_n917), .B2(new_n859), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n883), .A2(new_n885), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n674), .A2(new_n289), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n920), .B1(new_n922), .B2(new_n923), .ZN(G1346gat));
  NAND3_X1  g723(.A1(new_n922), .A2(KEYINPUT119), .A3(new_n584), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT119), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n926), .B1(new_n921), .B2(new_n680), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n925), .A2(G162gat), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n917), .A2(new_n290), .A3(new_n584), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(G1347gat));
  NOR2_X1   g729(.A1(new_n686), .A2(new_n460), .ZN(new_n931));
  AND3_X1   g730(.A1(new_n846), .A2(new_n465), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n622), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(G169gat), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT122), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n933), .A2(KEYINPUT122), .A3(G169gat), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n846), .A2(new_n931), .ZN(new_n939));
  OAI21_X1  g738(.A(KEYINPUT120), .B1(new_n939), .B2(new_n849), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT120), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n846), .A2(new_n941), .A3(new_n850), .A4(new_n931), .ZN(new_n942));
  NAND4_X1  g741(.A1(new_n940), .A2(new_n622), .A3(new_n250), .A4(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT121), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n943), .A2(new_n944), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n938), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(KEYINPUT123), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT123), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n938), .B(new_n949), .C1(new_n945), .C2(new_n946), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(G1348gat));
  AND2_X1   g750(.A1(new_n940), .A2(new_n942), .ZN(new_n952));
  AOI21_X1  g751(.A(G176gat), .B1(new_n952), .B2(new_n646), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n729), .A2(new_n210), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n953), .B1(new_n932), .B2(new_n954), .ZN(G1349gat));
  AOI21_X1  g754(.A(new_n222), .B1(new_n932), .B2(new_n675), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n859), .A2(new_n216), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n939), .A2(new_n849), .A3(new_n957), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n956), .A2(KEYINPUT124), .A3(new_n958), .ZN(new_n959));
  XOR2_X1   g758(.A(new_n959), .B(KEYINPUT60), .Z(G1350gat));
  AOI21_X1  g759(.A(new_n217), .B1(new_n932), .B2(new_n584), .ZN(new_n961));
  XOR2_X1   g760(.A(new_n961), .B(KEYINPUT61), .Z(new_n962));
  NAND3_X1  g761(.A1(new_n952), .A2(new_n217), .A3(new_n584), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(G1351gat));
  NAND2_X1  g763(.A1(new_n931), .A2(new_n663), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  OAI211_X1 g765(.A(new_n898), .B(new_n966), .C1(new_n899), .C2(new_n904), .ZN(new_n967));
  OAI21_X1  g766(.A(G197gat), .B1(new_n967), .B2(new_n623), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n869), .A2(new_n965), .ZN(new_n969));
  INV_X1    g768(.A(G197gat), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n969), .A2(new_n970), .A3(new_n622), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n968), .A2(new_n971), .ZN(G1352gat));
  NAND3_X1  g771(.A1(new_n969), .A2(new_n641), .A3(new_n646), .ZN(new_n973));
  XOR2_X1   g772(.A(new_n973), .B(KEYINPUT62), .Z(new_n974));
  OAI21_X1  g773(.A(G204gat), .B1(new_n905), .B2(new_n965), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(G1353gat));
  OAI21_X1  g775(.A(G211gat), .B1(new_n967), .B2(new_n508), .ZN(new_n977));
  OR2_X1    g776(.A1(new_n977), .A2(KEYINPUT63), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n969), .A2(new_n263), .A3(new_n859), .ZN(new_n979));
  XOR2_X1   g778(.A(new_n979), .B(KEYINPUT125), .Z(new_n980));
  NAND2_X1  g779(.A1(new_n977), .A2(KEYINPUT63), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n978), .A2(new_n980), .A3(new_n981), .ZN(G1354gat));
  NOR2_X1   g781(.A1(new_n680), .A2(new_n264), .ZN(new_n983));
  XNOR2_X1  g782(.A(new_n983), .B(KEYINPUT126), .ZN(new_n984));
  NOR3_X1   g783(.A1(new_n869), .A2(new_n680), .A3(new_n965), .ZN(new_n985));
  OAI22_X1  g784(.A1(new_n967), .A2(new_n984), .B1(G218gat), .B2(new_n985), .ZN(new_n986));
  XOR2_X1   g785(.A(new_n986), .B(KEYINPUT127), .Z(G1355gat));
endmodule


