//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 0 0 1 1 0 1 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 0 0 1 1 0 0 0 0 1 1 0 0 0 1 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n786, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n813,
    new_n814, new_n815, new_n816, new_n818, new_n819, new_n820, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1016, new_n1017, new_n1018, new_n1019;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202));
  INV_X1    g001(.A(G183gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT27), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT27), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G183gat), .ZN(new_n206));
  INV_X1    g005(.A(G190gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT69), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT28), .ZN(new_n210));
  AND3_X1   g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n210), .B1(new_n208), .B2(new_n209), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n202), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G169gat), .ZN(new_n214));
  INV_X1    g013(.A(G176gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n214), .A2(new_n215), .A3(KEYINPUT67), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT67), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(G169gat), .B2(G176gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT26), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n216), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT70), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n216), .A2(new_n218), .A3(KEYINPUT70), .A4(new_n219), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n214), .A2(new_n215), .ZN(new_n224));
  NAND2_X1  g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(new_n219), .ZN(new_n226));
  AOI22_X1  g025(.A1(new_n222), .A2(new_n223), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n228), .A2(new_n203), .A3(new_n207), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT24), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n202), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT64), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT64), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n236), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n231), .A2(new_n233), .A3(new_n235), .A4(new_n237), .ZN(new_n238));
  AND2_X1   g037(.A1(KEYINPUT66), .A2(G176gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(KEYINPUT66), .A2(G176gat), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT23), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n242), .A2(G169gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n225), .A2(KEYINPUT23), .ZN(new_n244));
  AOI22_X1  g043(.A1(new_n241), .A2(new_n243), .B1(new_n224), .B2(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT25), .B1(new_n238), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n203), .A2(new_n207), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n202), .B1(new_n248), .B2(KEYINPUT24), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n232), .A2(KEYINPUT68), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n247), .B(new_n234), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n216), .A2(new_n218), .A3(KEYINPUT23), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT25), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n253), .B1(new_n244), .B2(new_n224), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n251), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  OAI22_X1  g054(.A1(new_n213), .A2(new_n227), .B1(new_n246), .B2(new_n255), .ZN(new_n256));
  OR2_X1    g055(.A1(KEYINPUT72), .A2(G120gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(KEYINPUT72), .A2(G120gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n257), .A2(G113gat), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT73), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(G113gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT74), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT74), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(G113gat), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n263), .A2(new_n265), .A3(G120gat), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n257), .A2(KEYINPUT73), .A3(G113gat), .A4(new_n258), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n261), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G127gat), .B(G134gat), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT1), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  XOR2_X1   g071(.A(G113gat), .B(G120gat), .Z(new_n273));
  INV_X1    g072(.A(G134gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(G127gat), .ZN(new_n275));
  INV_X1    g074(.A(G127gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(G134gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n273), .A2(new_n270), .B1(new_n278), .B2(KEYINPUT71), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n269), .A2(new_n280), .ZN(new_n281));
  AOI22_X1  g080(.A1(new_n268), .A2(new_n272), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n256), .B(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT34), .ZN(new_n284));
  NAND2_X1  g083(.A1(G227gat), .A2(G233gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n284), .B1(new_n283), .B2(new_n285), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT32), .B1(new_n283), .B2(new_n285), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT33), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n291), .B1(new_n283), .B2(new_n285), .ZN(new_n292));
  XOR2_X1   g091(.A(G15gat), .B(G43gat), .Z(new_n293));
  XNOR2_X1  g092(.A(G71gat), .B(G99gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  AND3_X1   g094(.A1(new_n290), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n295), .ZN(new_n297));
  OAI221_X1 g096(.A(KEYINPUT32), .B1(new_n291), .B2(new_n297), .C1(new_n283), .C2(new_n285), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  OAI211_X1 g098(.A(KEYINPUT75), .B(new_n289), .C1(new_n296), .C2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT75), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n301), .B1(new_n287), .B2(new_n288), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n283), .A2(new_n285), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT34), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n304), .A2(KEYINPUT75), .A3(new_n286), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n290), .A2(new_n292), .A3(new_n295), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n302), .A2(new_n305), .A3(new_n298), .A4(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n300), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(KEYINPUT76), .A2(KEYINPUT36), .ZN(new_n309));
  OR2_X1    g108(.A1(KEYINPUT76), .A2(KEYINPUT36), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n300), .A2(new_n307), .A3(KEYINPUT76), .A4(KEYINPUT36), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(G8gat), .B(G36gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(G64gat), .B(G92gat), .ZN(new_n315));
  XOR2_X1   g114(.A(new_n314), .B(new_n315), .Z(new_n316));
  INV_X1    g115(.A(KEYINPUT81), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT80), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n256), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n222), .A2(new_n223), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n226), .A2(new_n224), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n208), .A2(new_n209), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT28), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n322), .A2(new_n202), .A3(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n251), .A2(new_n252), .A3(new_n254), .ZN(new_n328));
  OR2_X1    g127(.A1(KEYINPUT66), .A2(G176gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(KEYINPUT66), .A2(G176gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n243), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n244), .A2(new_n224), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI22_X1  g132(.A1(new_n229), .A2(new_n230), .B1(new_n232), .B2(new_n202), .ZN(new_n334));
  AND2_X1   g133(.A1(new_n235), .A2(new_n237), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n328), .B1(new_n336), .B2(KEYINPUT25), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n327), .A2(new_n337), .A3(KEYINPUT80), .ZN(new_n338));
  NAND2_X1  g137(.A1(G226gat), .A2(G233gat), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n319), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT79), .ZN(new_n342));
  INV_X1    g141(.A(G204gat), .ZN(new_n343));
  AND2_X1   g142(.A1(KEYINPUT77), .A2(G197gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(KEYINPUT77), .A2(G197gat), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n343), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT77), .ZN(new_n347));
  INV_X1    g146(.A(G197gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(KEYINPUT77), .A2(G197gat), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(G204gat), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(G211gat), .ZN(new_n353));
  INV_X1    g152(.A(G218gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G211gat), .A2(G218gat), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(KEYINPUT78), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT22), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n352), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n357), .B1(new_n352), .B2(new_n359), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n342), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NOR3_X1   g161(.A1(new_n344), .A2(new_n345), .A3(new_n343), .ZN(new_n363));
  AOI21_X1  g162(.A(G204gat), .B1(new_n349), .B2(new_n350), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n359), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n357), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n346), .A2(new_n351), .B1(new_n358), .B2(new_n356), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(new_n357), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n367), .A2(new_n369), .A3(KEYINPUT79), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n362), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT29), .B1(new_n327), .B2(new_n337), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n371), .B1(new_n372), .B2(new_n340), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n317), .B1(new_n341), .B2(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n340), .A2(KEYINPUT29), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n319), .A2(new_n338), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n327), .A2(new_n337), .A3(new_n340), .ZN(new_n377));
  INV_X1    g176(.A(new_n371), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n319), .A2(new_n338), .A3(new_n340), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT29), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n256), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n339), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n380), .A2(new_n383), .A3(KEYINPUT81), .A4(new_n371), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n374), .A2(new_n379), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n316), .B1(new_n385), .B2(KEYINPUT37), .ZN(new_n386));
  OAI22_X1  g185(.A1(new_n386), .A2(KEYINPUT94), .B1(KEYINPUT37), .B2(new_n385), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n384), .A2(new_n379), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n378), .B1(new_n339), .B2(new_n382), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT81), .B1(new_n389), .B2(new_n380), .ZN(new_n390));
  OAI21_X1  g189(.A(KEYINPUT37), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n316), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT94), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT38), .B1(new_n387), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(KEYINPUT83), .A2(KEYINPUT2), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(G141gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(G148gat), .ZN(new_n400));
  INV_X1    g199(.A(G148gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(G141gat), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n398), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(G155gat), .A2(G162gat), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT83), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(G155gat), .ZN(new_n407));
  INV_X1    g206(.A(G162gat), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(KEYINPUT83), .A2(G155gat), .A3(G162gat), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n406), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n403), .A2(new_n411), .ZN(new_n412));
  OR2_X1    g211(.A1(KEYINPUT84), .A2(G148gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(KEYINPUT84), .A2(G148gat), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n413), .A2(G141gat), .A3(new_n414), .ZN(new_n415));
  NOR2_X1   g214(.A1(G155gat), .A2(G162gat), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT2), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI22_X1  g217(.A1(new_n415), .A2(new_n400), .B1(new_n404), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT85), .B1(new_n412), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n404), .ZN(new_n421));
  AND2_X1   g220(.A1(KEYINPUT84), .A2(G148gat), .ZN(new_n422));
  NOR2_X1   g221(.A1(KEYINPUT84), .A2(G148gat), .ZN(new_n423));
  NOR3_X1   g222(.A1(new_n422), .A2(new_n423), .A3(new_n399), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n401), .A2(G141gat), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n421), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n416), .B1(new_n405), .B2(new_n404), .ZN(new_n427));
  XNOR2_X1  g226(.A(G141gat), .B(G148gat), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n427), .B(new_n410), .C1(new_n428), .C2(new_n398), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT85), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n426), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n282), .A2(KEYINPUT4), .A3(new_n420), .A4(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n267), .A2(new_n266), .ZN(new_n433));
  AND2_X1   g232(.A1(KEYINPUT72), .A2(G120gat), .ZN(new_n434));
  NOR2_X1   g233(.A1(KEYINPUT72), .A2(G120gat), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT73), .B1(new_n436), .B2(G113gat), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n272), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n415), .A2(new_n400), .ZN(new_n439));
  AND3_X1   g238(.A1(new_n406), .A2(new_n409), .A3(new_n410), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n399), .A2(G148gat), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n397), .B1(new_n425), .B2(new_n441), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n439), .A2(new_n421), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n279), .A2(new_n281), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n438), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT4), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(G225gat), .A2(G233gat), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT3), .B1(new_n412), .B2(new_n419), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT3), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n426), .A2(new_n429), .A3(new_n450), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n267), .A2(new_n266), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n271), .B1(new_n452), .B2(new_n261), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n273), .A2(new_n270), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n278), .A2(KEYINPUT71), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n454), .A2(new_n455), .A3(new_n281), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n449), .B(new_n451), .C1(new_n453), .C2(new_n456), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n432), .A2(new_n447), .A3(new_n448), .A4(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n448), .ZN(new_n459));
  INV_X1    g258(.A(new_n445), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n443), .B1(new_n438), .B2(new_n444), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n458), .A2(KEYINPUT5), .A3(new_n462), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n282), .A2(new_n446), .A3(new_n420), .A4(new_n431), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n445), .A2(KEYINPUT4), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT5), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n466), .A2(new_n467), .A3(new_n448), .A4(new_n457), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  XOR2_X1   g268(.A(G1gat), .B(G29gat), .Z(new_n470));
  XNOR2_X1  g269(.A(G57gat), .B(G85gat), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n470), .B(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(KEYINPUT86), .B(KEYINPUT0), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n472), .B(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n469), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT6), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n463), .A2(new_n474), .A3(new_n468), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n469), .A2(KEYINPUT6), .A3(new_n475), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n374), .A2(new_n316), .A3(new_n379), .A4(new_n384), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n385), .A2(KEYINPUT37), .ZN(new_n483));
  XOR2_X1   g282(.A(new_n316), .B(KEYINPUT82), .Z(new_n484));
  NOR3_X1   g283(.A1(new_n483), .A2(KEYINPUT38), .A3(new_n484), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n376), .A2(new_n377), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n371), .B1(new_n380), .B2(new_n383), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT93), .ZN(new_n488));
  OAI22_X1  g287(.A1(new_n486), .A2(new_n378), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n487), .A2(new_n488), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT37), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n482), .B1(new_n485), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n396), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n451), .A2(new_n381), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n362), .A2(new_n370), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(G228gat), .A2(G233gat), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n450), .B1(new_n426), .B2(new_n429), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n367), .A2(new_n369), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT29), .B1(new_n426), .B2(new_n429), .ZN(new_n501));
  AOI211_X1 g300(.A(KEYINPUT90), .B(new_n499), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT90), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n501), .B1(new_n360), .B2(new_n361), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n503), .B1(new_n504), .B2(new_n449), .ZN(new_n505));
  NOR3_X1   g304(.A1(new_n498), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  XOR2_X1   g305(.A(new_n496), .B(KEYINPUT89), .Z(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n420), .A2(new_n431), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n355), .A2(new_n356), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n365), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n368), .A2(new_n510), .ZN(new_n513));
  AND3_X1   g312(.A1(new_n512), .A2(new_n381), .A3(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n509), .B1(new_n514), .B2(KEYINPUT3), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n508), .B1(new_n515), .B2(new_n495), .ZN(new_n516));
  OAI21_X1  g315(.A(G22gat), .B1(new_n506), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n495), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(new_n507), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n449), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT90), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n504), .A2(new_n503), .A3(new_n449), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n521), .A2(new_n522), .A3(new_n495), .A4(new_n497), .ZN(new_n523));
  INV_X1    g322(.A(G22gat), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n519), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G78gat), .B(G106gat), .ZN(new_n526));
  INV_X1    g325(.A(G50gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(KEYINPUT88), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(KEYINPUT31), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n517), .A2(new_n525), .A3(KEYINPUT91), .A4(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n517), .A2(KEYINPUT91), .A3(new_n525), .ZN(new_n532));
  INV_X1    g331(.A(new_n530), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT91), .B1(new_n517), .B2(new_n525), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n531), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n481), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT30), .ZN(new_n538));
  INV_X1    g337(.A(new_n484), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n385), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT30), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n481), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n538), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n448), .B1(new_n466), .B2(new_n457), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT39), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n461), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n547), .A2(new_n448), .A3(new_n445), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT92), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n547), .A2(KEYINPUT92), .A3(new_n448), .A4(new_n445), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n546), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n475), .B1(new_n544), .B2(new_n545), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n553), .A2(KEYINPUT40), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(KEYINPUT40), .B1(new_n553), .B2(new_n554), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n474), .B1(new_n463), .B2(new_n468), .ZN(new_n557));
  NOR3_X1   g356(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n536), .B1(new_n543), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n313), .B1(new_n493), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT87), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n478), .A2(new_n477), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n562), .A2(new_n557), .ZN(new_n563));
  INV_X1    g362(.A(new_n480), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n542), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n540), .B1(new_n541), .B2(new_n481), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n561), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AOI22_X1  g366(.A1(new_n537), .A2(KEYINPUT30), .B1(new_n539), .B2(new_n385), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n479), .A2(new_n480), .B1(new_n541), .B2(new_n481), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n568), .A2(new_n569), .A3(KEYINPUT87), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n567), .A2(new_n570), .A3(new_n536), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n560), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n567), .A2(new_n570), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n536), .B1(new_n300), .B2(new_n307), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT35), .ZN(new_n576));
  NOR3_X1   g375(.A1(new_n565), .A2(new_n566), .A3(KEYINPUT35), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n572), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT99), .ZN(new_n581));
  XNOR2_X1  g380(.A(G57gat), .B(G64gat), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G71gat), .B(G78gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT21), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G127gat), .B(G155gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT20), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n590), .B(new_n592), .ZN(new_n593));
  XOR2_X1   g392(.A(G183gat), .B(G211gat), .Z(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G15gat), .B(G22gat), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT16), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n596), .B1(new_n597), .B2(G1gat), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n598), .B1(G1gat), .B2(new_n596), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(G8gat), .ZN(new_n600));
  INV_X1    g399(.A(G8gat), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n598), .B(new_n601), .C1(G1gat), .C2(new_n596), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n586), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n603), .B1(new_n604), .B2(KEYINPUT21), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT103), .ZN(new_n606));
  XOR2_X1   g405(.A(KEYINPUT100), .B(KEYINPUT101), .Z(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT102), .B(KEYINPUT19), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n606), .B(new_n609), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n595), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n610), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G99gat), .A2(G106gat), .ZN(new_n614));
  INV_X1    g413(.A(G85gat), .ZN(new_n615));
  INV_X1    g414(.A(G92gat), .ZN(new_n616));
  AOI22_X1  g415(.A1(KEYINPUT8), .A2(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT104), .ZN(new_n618));
  NAND2_X1  g417(.A1(G85gat), .A2(G92gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT7), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(G99gat), .B(G106gat), .Z(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n622), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n618), .A2(new_n624), .A3(new_n620), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(G43gat), .B(G50gat), .Z(new_n628));
  INV_X1    g427(.A(KEYINPUT15), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G43gat), .B(G50gat), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(KEYINPUT15), .ZN(new_n632));
  INV_X1    g431(.A(G29gat), .ZN(new_n633));
  INV_X1    g432(.A(G36gat), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(G29gat), .A2(G36gat), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n635), .B1(KEYINPUT14), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT14), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n638), .B1(G29gat), .B2(G36gat), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n630), .A2(new_n632), .A3(new_n637), .A4(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n636), .A2(KEYINPUT14), .ZN(new_n641));
  OAI211_X1 g440(.A(new_n641), .B(new_n639), .C1(new_n633), .C2(new_n634), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n642), .A2(KEYINPUT15), .A3(new_n631), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g443(.A1(G232gat), .A2(G233gat), .ZN(new_n645));
  AOI22_X1  g444(.A1(new_n627), .A2(new_n644), .B1(KEYINPUT41), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n626), .A2(KEYINPUT105), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n640), .A2(KEYINPUT17), .A3(new_n643), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT17), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n644), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n647), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n626), .A2(KEYINPUT105), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n646), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(G190gat), .B(G218gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n645), .A2(KEYINPUT41), .ZN(new_n656));
  XNOR2_X1  g455(.A(G134gat), .B(G162gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n655), .B(new_n658), .Z(new_n659));
  NOR2_X1   g458(.A1(new_n613), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n626), .A2(new_n586), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT10), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n604), .A2(new_n623), .A3(new_n625), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n627), .A2(KEYINPUT10), .A3(new_n604), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(G230gat), .A2(G233gat), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n661), .A2(new_n663), .ZN(new_n669));
  INV_X1    g468(.A(new_n667), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(G120gat), .B(G148gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(G176gat), .B(G204gat), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n673), .B(new_n674), .Z(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n668), .A2(new_n671), .A3(new_n675), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n660), .A2(new_n680), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n600), .A2(new_n602), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(new_n644), .ZN(new_n683));
  NAND2_X1  g482(.A1(G229gat), .A2(G233gat), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n684), .B(KEYINPUT13), .Z(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n682), .A2(new_n650), .A3(KEYINPUT96), .A4(new_n648), .ZN(new_n688));
  INV_X1    g487(.A(new_n648), .ZN(new_n689));
  AOI21_X1  g488(.A(KEYINPUT17), .B1(new_n640), .B2(new_n643), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n689), .A2(new_n603), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n603), .A2(new_n644), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT96), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n688), .B1(new_n691), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(new_n684), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT18), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n687), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n695), .A2(KEYINPUT18), .A3(new_n684), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(KEYINPUT97), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT97), .ZN(new_n701));
  INV_X1    g500(.A(new_n684), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n682), .A2(new_n648), .A3(new_n650), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n703), .A2(new_n693), .A3(new_n692), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n702), .B1(new_n704), .B2(new_n688), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n701), .B1(new_n705), .B2(KEYINPUT18), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n698), .B1(new_n700), .B2(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(G113gat), .B(G141gat), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT95), .B(G197gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(KEYINPUT11), .B(G169gat), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n712), .B(KEYINPUT12), .Z(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n696), .A2(new_n697), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT98), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n707), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n705), .A2(KEYINPUT18), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n713), .B1(new_n719), .B2(KEYINPUT98), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n699), .A2(KEYINPUT97), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n705), .A2(new_n701), .A3(KEYINPUT18), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n720), .A2(new_n723), .A3(new_n698), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n718), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n681), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n580), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n479), .A2(new_n480), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XOR2_X1   g529(.A(new_n730), .B(G1gat), .Z(G1324gat));
  INV_X1    g530(.A(new_n728), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n601), .B1(new_n732), .B2(new_n543), .ZN(new_n733));
  INV_X1    g532(.A(new_n543), .ZN(new_n734));
  XNOR2_X1  g533(.A(KEYINPUT16), .B(G8gat), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n728), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(KEYINPUT42), .B1(new_n733), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(KEYINPUT42), .B2(new_n736), .ZN(G1325gat));
  AND2_X1   g537(.A1(new_n311), .A2(new_n312), .ZN(new_n739));
  OAI21_X1  g538(.A(G15gat), .B1(new_n728), .B2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n308), .ZN(new_n741));
  OR2_X1    g540(.A1(new_n741), .A2(G15gat), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n740), .B1(new_n728), .B2(new_n742), .ZN(G1326gat));
  INV_X1    g542(.A(new_n536), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n728), .A2(new_n744), .ZN(new_n745));
  XOR2_X1   g544(.A(KEYINPUT43), .B(G22gat), .Z(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1327gat));
  NAND2_X1  g546(.A1(new_n571), .A2(KEYINPUT106), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT38), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n483), .B1(new_n393), .B2(new_n394), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n386), .A2(KEYINPUT94), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n484), .A2(KEYINPUT38), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n491), .B(new_n753), .C1(KEYINPUT37), .C2(new_n385), .ZN(new_n754));
  INV_X1    g553(.A(new_n482), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n559), .B1(new_n752), .B2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT106), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n567), .A2(new_n570), .A3(new_n758), .A4(new_n536), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n748), .A2(new_n757), .A3(new_n739), .A4(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT107), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n560), .A2(KEYINPUT107), .A3(new_n748), .A4(new_n759), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n579), .ZN(new_n765));
  INV_X1    g564(.A(new_n659), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n766), .A2(KEYINPUT44), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n765), .A2(KEYINPUT108), .A3(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT108), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n576), .A2(new_n578), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n770), .B1(new_n762), .B2(new_n763), .ZN(new_n771));
  INV_X1    g570(.A(new_n767), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n769), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n766), .B1(new_n572), .B2(new_n579), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT44), .ZN(new_n775));
  OR2_X1    g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n768), .A2(new_n773), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n613), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n778), .A2(new_n726), .A3(new_n679), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(G29gat), .B1(new_n780), .B2(new_n729), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n774), .A2(new_n779), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n782), .A2(G29gat), .A3(new_n729), .ZN(new_n783));
  XOR2_X1   g582(.A(new_n783), .B(KEYINPUT45), .Z(new_n784));
  NAND2_X1  g583(.A1(new_n781), .A2(new_n784), .ZN(G1328gat));
  OAI21_X1  g584(.A(G36gat), .B1(new_n780), .B2(new_n734), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n782), .A2(G36gat), .A3(new_n734), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT46), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(G1329gat));
  NAND2_X1  g588(.A1(new_n313), .A2(G43gat), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n782), .A2(new_n741), .ZN(new_n791));
  OAI22_X1  g590(.A1(new_n780), .A2(new_n790), .B1(G43gat), .B2(new_n791), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g592(.A(new_n527), .B1(new_n782), .B2(new_n744), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n536), .A2(G50gat), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n794), .B1(new_n780), .B2(new_n795), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT48), .ZN(G1331gat));
  NOR4_X1   g596(.A1(new_n613), .A2(new_n659), .A3(new_n725), .A4(new_n680), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n765), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n729), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(G57gat), .ZN(G1332gat));
  OR2_X1    g602(.A1(new_n543), .A2(KEYINPUT109), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n543), .A2(KEYINPUT109), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n799), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n809));
  AND2_X1   g608(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n808), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n811), .B1(new_n808), .B2(new_n809), .ZN(G1333gat));
  XOR2_X1   g611(.A(new_n308), .B(KEYINPUT110), .Z(new_n813));
  AOI21_X1  g612(.A(G71gat), .B1(new_n800), .B2(new_n813), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n313), .A2(G71gat), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n814), .B1(new_n800), .B2(new_n815), .ZN(new_n816));
  XOR2_X1   g615(.A(new_n816), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g616(.A1(new_n800), .A2(new_n536), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(KEYINPUT112), .ZN(new_n819));
  XNOR2_X1  g618(.A(KEYINPUT111), .B(G78gat), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n819), .B(new_n820), .ZN(G1335gat));
  NOR3_X1   g620(.A1(new_n778), .A2(new_n766), .A3(new_n725), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n765), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n823), .B(KEYINPUT51), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n824), .B(KEYINPUT113), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n801), .A2(new_n615), .A3(new_n679), .ZN(new_n826));
  XOR2_X1   g625(.A(new_n826), .B(KEYINPUT114), .Z(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n778), .A2(new_n725), .A3(new_n680), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n777), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(G85gat), .B1(new_n830), .B2(new_n729), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n828), .A2(new_n831), .ZN(G1336gat));
  OAI21_X1  g631(.A(G92gat), .B1(new_n830), .B2(new_n807), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n806), .A2(new_n616), .A3(new_n679), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n833), .B(new_n834), .C1(new_n824), .C2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n777), .A2(new_n543), .A3(new_n829), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n837), .A2(KEYINPUT115), .A3(G92gat), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT115), .B1(new_n837), .B2(G92gat), .ZN(new_n839));
  XOR2_X1   g638(.A(new_n835), .B(KEYINPUT116), .Z(new_n840));
  NOR2_X1   g639(.A1(new_n824), .A2(new_n840), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n838), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n836), .B1(new_n842), .B2(new_n834), .ZN(G1337gat));
  NOR3_X1   g642(.A1(new_n741), .A2(G99gat), .A3(new_n680), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n825), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(G99gat), .B1(new_n830), .B2(new_n739), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(G1338gat));
  OAI21_X1  g646(.A(G106gat), .B1(new_n830), .B2(new_n744), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT51), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n823), .B(new_n849), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n744), .A2(G106gat), .A3(new_n680), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  XOR2_X1   g652(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n854));
  XNOR2_X1  g653(.A(new_n853), .B(new_n854), .ZN(G1339gat));
  NAND3_X1  g654(.A1(new_n660), .A2(new_n726), .A3(new_n680), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n664), .A2(new_n665), .A3(new_n670), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n668), .A2(KEYINPUT54), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n670), .B1(new_n664), .B2(new_n665), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n675), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n858), .A2(KEYINPUT55), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n678), .ZN(new_n863));
  AOI21_X1  g662(.A(KEYINPUT55), .B1(new_n858), .B2(new_n861), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n725), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n723), .A2(new_n714), .A3(new_n698), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n683), .A2(new_n686), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n868), .B1(new_n684), .B2(new_n695), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n712), .ZN(new_n870));
  AND3_X1   g669(.A1(new_n679), .A2(new_n867), .A3(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n659), .B1(new_n866), .B2(new_n872), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n867), .A2(new_n870), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n659), .A2(new_n874), .A3(new_n865), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n856), .B1(new_n877), .B2(new_n778), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(KEYINPUT118), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT118), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n880), .B(new_n856), .C1(new_n877), .C2(new_n778), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(new_n801), .A3(new_n574), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n883), .A2(new_n806), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n884), .A2(new_n263), .A3(new_n265), .A4(new_n725), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n806), .A2(new_n729), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n882), .A2(new_n744), .A3(new_n308), .A4(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(G113gat), .B1(new_n887), .B2(new_n726), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n885), .A2(new_n888), .ZN(G1340gat));
  NAND3_X1  g688(.A1(new_n884), .A2(new_n436), .A3(new_n679), .ZN(new_n890));
  OAI21_X1  g689(.A(G120gat), .B1(new_n887), .B2(new_n680), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(G1341gat));
  NAND3_X1  g691(.A1(new_n884), .A2(new_n276), .A3(new_n778), .ZN(new_n893));
  OAI21_X1  g692(.A(G127gat), .B1(new_n887), .B2(new_n613), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(G1342gat));
  NAND3_X1  g694(.A1(new_n659), .A2(new_n274), .A3(new_n734), .ZN(new_n896));
  OR3_X1    g695(.A1(new_n883), .A2(KEYINPUT56), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(G134gat), .B1(new_n887), .B2(new_n766), .ZN(new_n898));
  OAI21_X1  g697(.A(KEYINPUT56), .B1(new_n883), .B2(new_n896), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(G1343gat));
  NAND3_X1  g699(.A1(new_n879), .A2(new_n536), .A3(new_n881), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT57), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n744), .A2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT119), .ZN(new_n904));
  AND3_X1   g703(.A1(new_n664), .A2(new_n665), .A3(new_n670), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n905), .A2(new_n859), .A3(new_n860), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n666), .A2(new_n860), .A3(new_n667), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n676), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n904), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT55), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n858), .A2(KEYINPUT119), .A3(new_n861), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n862), .A2(new_n678), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n725), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n872), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n659), .B1(new_n915), .B2(KEYINPUT120), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n863), .B1(new_n724), .B2(new_n718), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n871), .B1(new_n917), .B2(new_n912), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT120), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n876), .B1(new_n916), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n856), .B1(new_n921), .B2(new_n778), .ZN(new_n922));
  AOI22_X1  g721(.A1(new_n901), .A2(new_n902), .B1(new_n903), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n886), .A2(new_n739), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n399), .B1(new_n925), .B2(new_n725), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n313), .A2(new_n744), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n882), .A2(new_n801), .A3(new_n927), .ZN(new_n928));
  NOR4_X1   g727(.A1(new_n928), .A2(G141gat), .A3(new_n726), .A4(new_n806), .ZN(new_n929));
  OR3_X1    g728(.A1(new_n926), .A2(KEYINPUT58), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(KEYINPUT58), .B1(new_n926), .B2(new_n929), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(G1344gat));
  INV_X1    g731(.A(new_n928), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n413), .A2(new_n414), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n933), .A2(new_n935), .A3(new_n679), .A4(new_n807), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT59), .ZN(new_n937));
  INV_X1    g736(.A(new_n924), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n882), .A2(new_n903), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT121), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n744), .B1(new_n922), .B2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(new_n856), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n766), .B1(new_n918), .B2(new_n919), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n915), .A2(KEYINPUT120), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n875), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n942), .B1(new_n945), .B2(new_n613), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(KEYINPUT121), .ZN(new_n947));
  AOI21_X1  g746(.A(KEYINPUT57), .B1(new_n941), .B2(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT122), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n939), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n536), .B1(new_n946), .B2(KEYINPUT121), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n922), .A2(new_n940), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n902), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n953), .A2(KEYINPUT122), .ZN(new_n954));
  OAI211_X1 g753(.A(new_n679), .B(new_n938), .C1(new_n950), .C2(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n937), .B1(new_n955), .B2(G148gat), .ZN(new_n956));
  AOI211_X1 g755(.A(KEYINPUT59), .B(new_n935), .C1(new_n925), .C2(new_n679), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n936), .B1(new_n956), .B2(new_n957), .ZN(G1345gat));
  NAND2_X1  g757(.A1(new_n933), .A2(new_n807), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n778), .A2(new_n407), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n923), .A2(new_n613), .A3(new_n924), .ZN(new_n961));
  OAI22_X1  g760(.A1(new_n959), .A2(new_n960), .B1(new_n961), .B2(new_n407), .ZN(G1346gat));
  NOR3_X1   g761(.A1(new_n923), .A2(new_n766), .A3(new_n924), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n659), .A2(new_n408), .A3(new_n734), .ZN(new_n964));
  OAI22_X1  g763(.A1(new_n963), .A2(new_n408), .B1(new_n928), .B2(new_n964), .ZN(G1347gat));
  NOR2_X1   g764(.A1(new_n734), .A2(new_n801), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n813), .A2(new_n966), .ZN(new_n967));
  NAND4_X1  g766(.A1(new_n879), .A2(new_n744), .A3(new_n881), .A4(new_n967), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n968), .A2(new_n214), .A3(new_n726), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n882), .A2(new_n729), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n970), .A2(new_n574), .A3(new_n806), .ZN(new_n971));
  OR2_X1    g770(.A1(new_n971), .A2(new_n726), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n969), .B1(new_n972), .B2(new_n214), .ZN(G1348gat));
  NOR3_X1   g772(.A1(new_n968), .A2(new_n241), .A3(new_n680), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n215), .B1(new_n971), .B2(new_n680), .ZN(new_n975));
  OR2_X1    g774(.A1(new_n975), .A2(KEYINPUT123), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(KEYINPUT123), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n974), .B1(new_n976), .B2(new_n977), .ZN(G1349gat));
  NAND3_X1  g777(.A1(new_n778), .A2(new_n204), .A3(new_n206), .ZN(new_n979));
  OAI21_X1  g778(.A(KEYINPUT124), .B1(new_n968), .B2(new_n613), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(G183gat), .ZN(new_n981));
  NOR3_X1   g780(.A1(new_n968), .A2(KEYINPUT124), .A3(new_n613), .ZN(new_n982));
  OAI22_X1  g781(.A1(new_n971), .A2(new_n979), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  XNOR2_X1  g782(.A(new_n983), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g783(.A(G190gat), .B1(new_n968), .B2(new_n766), .ZN(new_n985));
  OR2_X1    g784(.A1(new_n985), .A2(KEYINPUT61), .ZN(new_n986));
  INV_X1    g785(.A(new_n986), .ZN(new_n987));
  AND2_X1   g786(.A1(new_n985), .A2(KEYINPUT61), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n659), .A2(new_n207), .ZN(new_n989));
  OAI22_X1  g788(.A1(new_n987), .A2(new_n988), .B1(new_n971), .B2(new_n989), .ZN(G1351gat));
  AND3_X1   g789(.A1(new_n970), .A2(new_n806), .A3(new_n927), .ZN(new_n991));
  AOI21_X1  g790(.A(G197gat), .B1(new_n991), .B2(new_n725), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n953), .A2(KEYINPUT122), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n948), .A2(new_n949), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n993), .A2(new_n994), .A3(new_n939), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n739), .A2(new_n966), .ZN(new_n996));
  XOR2_X1   g795(.A(new_n996), .B(KEYINPUT125), .Z(new_n997));
  NOR3_X1   g796(.A1(new_n997), .A2(new_n348), .A3(new_n726), .ZN(new_n998));
  AOI21_X1  g797(.A(new_n992), .B1(new_n995), .B2(new_n998), .ZN(G1352gat));
  NAND2_X1  g798(.A1(new_n995), .A2(new_n679), .ZN(new_n1000));
  OAI21_X1  g799(.A(G204gat), .B1(new_n1000), .B2(new_n997), .ZN(new_n1001));
  NOR2_X1   g800(.A1(new_n680), .A2(G204gat), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n991), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1003), .A2(KEYINPUT62), .ZN(new_n1004));
  OR2_X1    g803(.A1(new_n1003), .A2(KEYINPUT62), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n1001), .A2(new_n1004), .A3(new_n1005), .ZN(G1353gat));
  NAND3_X1  g805(.A1(new_n991), .A2(new_n353), .A3(new_n778), .ZN(new_n1007));
  NOR2_X1   g806(.A1(new_n996), .A2(new_n613), .ZN(new_n1008));
  OAI21_X1  g807(.A(new_n1008), .B1(new_n950), .B2(new_n954), .ZN(new_n1009));
  INV_X1    g808(.A(KEYINPUT63), .ZN(new_n1010));
  NOR2_X1   g809(.A1(new_n1010), .A2(KEYINPUT126), .ZN(new_n1011));
  AOI21_X1  g810(.A(new_n353), .B1(KEYINPUT126), .B2(new_n1010), .ZN(new_n1012));
  AND3_X1   g811(.A1(new_n1009), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g812(.A(new_n1011), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1014));
  OAI21_X1  g813(.A(new_n1007), .B1(new_n1013), .B2(new_n1014), .ZN(G1354gat));
  AOI21_X1  g814(.A(G218gat), .B1(new_n991), .B2(new_n659), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n659), .A2(G218gat), .ZN(new_n1017));
  XNOR2_X1  g816(.A(new_n1017), .B(KEYINPUT127), .ZN(new_n1018));
  NOR2_X1   g817(.A1(new_n997), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g818(.A(new_n1016), .B1(new_n995), .B2(new_n1019), .ZN(G1355gat));
endmodule


