//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 1 0 0 0 0 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n777, new_n778,
    new_n779, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT11), .ZN(new_n192));
  INV_X1    g006(.A(G134), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(G137), .ZN(new_n194));
  INV_X1    g008(.A(G137), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(KEYINPUT11), .A3(G134), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n193), .A2(G137), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G131), .ZN(new_n199));
  INV_X1    g013(.A(G131), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n194), .A2(new_n196), .A3(new_n200), .A4(new_n197), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT12), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  AND2_X1   g019(.A1(KEYINPUT66), .A2(G143), .ZN(new_n206));
  NOR2_X1   g020(.A1(KEYINPUT66), .A2(G143), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n205), .A2(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT1), .ZN(new_n212));
  AOI22_X1  g026(.A1(new_n208), .A2(new_n210), .B1(new_n212), .B2(G128), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(new_n209), .ZN(new_n215));
  NAND2_X1  g029(.A1(KEYINPUT66), .A2(G143), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(G146), .A3(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G128), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n217), .A2(new_n211), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT68), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT68), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n217), .A2(new_n222), .A3(new_n211), .A4(new_n219), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n213), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G104), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G107), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n225), .A2(G107), .ZN(new_n228));
  OAI21_X1  g042(.A(G101), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(KEYINPUT3), .B1(new_n225), .B2(G107), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n231));
  INV_X1    g045(.A(G107), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(new_n232), .A3(G104), .ZN(new_n233));
  INV_X1    g047(.A(G101), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n230), .A2(new_n233), .A3(new_n234), .A4(new_n226), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n229), .A2(new_n235), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n224), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n221), .A2(new_n223), .ZN(new_n238));
  AOI21_X1  g052(.A(G146), .B1(new_n215), .B2(new_n216), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT1), .ZN(new_n240));
  OAI21_X1  g054(.A(G128), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n217), .A2(new_n211), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n236), .B1(new_n238), .B2(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n204), .B1(new_n237), .B2(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(KEYINPUT71), .B1(new_n199), .B2(new_n201), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n199), .A2(KEYINPUT71), .A3(new_n201), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n211), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n206), .A2(new_n207), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n250), .B1(new_n251), .B2(G146), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n222), .B1(new_n252), .B2(new_n219), .ZN(new_n253));
  INV_X1    g067(.A(new_n223), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n243), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n236), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n224), .A2(new_n236), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n249), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n245), .B1(new_n259), .B2(KEYINPUT12), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT10), .ZN(new_n261));
  AOI22_X1  g075(.A1(new_n221), .A2(new_n223), .B1(new_n241), .B2(new_n242), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n261), .B1(new_n262), .B2(new_n236), .ZN(new_n263));
  INV_X1    g077(.A(new_n213), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n238), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n236), .A2(new_n261), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT0), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n268), .A2(new_n218), .A3(KEYINPUT64), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT64), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n270), .B1(KEYINPUT0), .B2(G128), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  AND3_X1   g086(.A1(KEYINPUT65), .A2(KEYINPUT0), .A3(G128), .ZN(new_n273));
  AOI21_X1  g087(.A(KEYINPUT65), .B1(KEYINPUT0), .B2(G128), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n208), .A2(new_n210), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n268), .A2(new_n218), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n276), .A2(new_n277), .B1(new_n252), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n230), .A2(new_n233), .A3(new_n226), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT4), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n281), .A3(G101), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(G101), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n283), .A2(KEYINPUT4), .A3(new_n235), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n279), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n263), .A2(new_n267), .A3(new_n249), .A4(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n260), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G953), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G227), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n289), .B(KEYINPUT85), .ZN(new_n290));
  XNOR2_X1  g104(.A(G110), .B(G140), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n290), .B(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n287), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT87), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n199), .A2(KEYINPUT71), .A3(new_n201), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n295), .A2(new_n246), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n244), .A2(KEYINPUT10), .ZN(new_n297));
  INV_X1    g111(.A(new_n266), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n284), .A2(new_n282), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n277), .A2(new_n272), .A3(new_n275), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n252), .A2(new_n278), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI22_X1  g116(.A1(new_n298), .A2(new_n224), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n294), .B(new_n296), .C1(new_n297), .C2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n263), .A2(new_n267), .A3(new_n285), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n294), .B1(new_n306), .B2(new_n296), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT86), .ZN(new_n308));
  INV_X1    g122(.A(new_n292), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n286), .A2(new_n309), .ZN(new_n310));
  OAI22_X1  g124(.A1(new_n305), .A2(new_n307), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  AND2_X1   g125(.A1(new_n286), .A2(new_n309), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n312), .A2(KEYINPUT86), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n293), .B(G469), .C1(new_n311), .C2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(G469), .A2(G902), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G469), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n306), .A2(new_n296), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT87), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n304), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n309), .B1(new_n320), .B2(new_n286), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n258), .B1(new_n236), .B2(new_n262), .ZN(new_n322));
  AOI21_X1  g136(.A(KEYINPUT12), .B1(new_n322), .B2(new_n296), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n203), .B1(new_n257), .B2(new_n258), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT88), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT88), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n245), .B(new_n326), .C1(new_n259), .C2(KEYINPUT12), .ZN(new_n327));
  AND3_X1   g141(.A1(new_n325), .A2(new_n327), .A3(new_n312), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n317), .B(new_n190), .C1(new_n321), .C2(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n191), .B1(new_n316), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G475), .ZN(new_n332));
  INV_X1    g146(.A(G140), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G125), .ZN(new_n334));
  INV_X1    g148(.A(G125), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G140), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT81), .ZN(new_n338));
  XNOR2_X1  g152(.A(G125), .B(G140), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT81), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n338), .A2(new_n341), .A3(new_n205), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n339), .A2(new_n205), .ZN(new_n343));
  INV_X1    g157(.A(G237), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(new_n288), .A3(G214), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(new_n215), .A3(new_n216), .ZN(new_n346));
  NAND2_X1  g160(.A1(KEYINPUT18), .A2(G131), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n344), .A2(new_n288), .A3(G143), .A4(G214), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n346), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n348), .B1(new_n346), .B2(new_n349), .ZN(new_n352));
  OAI22_X1  g166(.A1(new_n342), .A2(new_n343), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n346), .A2(new_n200), .A3(new_n349), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n200), .B1(new_n346), .B2(new_n349), .ZN(new_n356));
  NOR3_X1   g170(.A1(new_n355), .A2(new_n356), .A3(KEYINPUT17), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n346), .A2(new_n349), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n358), .A2(KEYINPUT17), .A3(G131), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n334), .A2(new_n336), .A3(KEYINPUT16), .ZN(new_n360));
  OR3_X1    g174(.A1(new_n335), .A2(KEYINPUT16), .A3(G140), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n205), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n360), .A2(new_n361), .A3(G146), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n359), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n353), .B1(new_n357), .B2(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(G113), .B(G122), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n367), .B(new_n225), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n353), .B(new_n368), .C1(new_n357), .C2(new_n365), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n332), .B1(new_n372), .B2(new_n190), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n371), .ZN(new_n375));
  INV_X1    g189(.A(new_n364), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n358), .A2(G131), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n376), .B1(new_n377), .B2(new_n354), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT19), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n338), .A2(new_n341), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n337), .A2(KEYINPUT19), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n205), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n358), .A2(new_n347), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n350), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n338), .A2(new_n341), .A3(new_n205), .ZN(new_n385));
  INV_X1    g199(.A(new_n343), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI22_X1  g201(.A1(new_n378), .A2(new_n382), .B1(new_n384), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n368), .B1(new_n388), .B2(KEYINPUT91), .ZN(new_n389));
  INV_X1    g203(.A(new_n382), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n364), .B1(new_n355), .B2(new_n356), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n353), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT91), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n375), .B1(new_n389), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(G475), .A2(G902), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NOR3_X1   g211(.A1(new_n395), .A2(KEYINPUT20), .A3(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT20), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n353), .B(KEYINPUT91), .C1(new_n390), .C2(new_n391), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n369), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n378), .A2(new_n382), .ZN(new_n402));
  AOI21_X1  g216(.A(KEYINPUT91), .B1(new_n402), .B2(new_n353), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n371), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n399), .B1(new_n404), .B2(new_n396), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n374), .B1(new_n398), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT92), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(KEYINPUT20), .B1(new_n395), .B2(new_n397), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n404), .A2(new_n399), .A3(new_n396), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(KEYINPUT92), .A3(new_n374), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n408), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G116), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G122), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n414), .A2(G122), .ZN(new_n417));
  NOR3_X1   g231(.A1(new_n416), .A2(new_n417), .A3(G107), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n415), .A2(KEYINPUT14), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n415), .B1(new_n417), .B2(KEYINPUT14), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n419), .B1(new_n420), .B2(KEYINPUT95), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n421), .B1(KEYINPUT95), .B2(new_n420), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n418), .B1(new_n422), .B2(G107), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n215), .A2(new_n216), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n424), .A2(new_n218), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n209), .A2(G128), .ZN(new_n426));
  OAI21_X1  g240(.A(G134), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n251), .A2(G128), .ZN(new_n428));
  INV_X1    g242(.A(new_n426), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n428), .A2(new_n193), .A3(new_n429), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n427), .A2(KEYINPUT94), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(KEYINPUT94), .B1(new_n427), .B2(new_n430), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n423), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n416), .A2(new_n417), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n434), .A2(new_n232), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT93), .ZN(new_n436));
  OR3_X1    g250(.A1(new_n435), .A2(new_n436), .A3(new_n418), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n428), .A2(KEYINPUT13), .A3(new_n429), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n438), .B(G134), .C1(KEYINPUT13), .C2(new_n428), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n436), .B1(new_n435), .B2(new_n418), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n437), .A2(new_n439), .A3(new_n430), .A4(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G217), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n188), .A2(new_n442), .A3(G953), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n433), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n443), .B1(new_n433), .B2(new_n441), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n190), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(G478), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n447), .A2(KEYINPUT15), .ZN(new_n448));
  XOR2_X1   g262(.A(new_n446), .B(new_n448), .Z(new_n449));
  NAND2_X1  g263(.A1(new_n413), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(G110), .B(G122), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n414), .A2(G119), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(G113), .B1(new_n454), .B2(KEYINPUT5), .ZN(new_n455));
  INV_X1    g269(.A(G119), .ZN(new_n456));
  OAI21_X1  g270(.A(KEYINPUT69), .B1(new_n456), .B2(G116), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT69), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n458), .A2(new_n414), .A3(G119), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n454), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT70), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n453), .B1(new_n457), .B2(new_n459), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT70), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n455), .B1(new_n466), .B2(KEYINPUT5), .ZN(new_n467));
  XNOR2_X1  g281(.A(KEYINPUT2), .B(G113), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n464), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n256), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n463), .A2(new_n465), .A3(new_n468), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n299), .B1(new_n473), .B2(new_n470), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n452), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n473), .A2(new_n470), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n476), .A2(new_n282), .A3(new_n284), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n477), .B(new_n451), .C1(new_n467), .C2(new_n471), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n475), .A2(new_n478), .A3(KEYINPUT6), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n302), .A2(G125), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n480), .B1(new_n265), .B2(G125), .ZN(new_n481));
  INV_X1    g295(.A(G224), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n482), .A2(G953), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n483), .B(KEYINPUT89), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n481), .B(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT6), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n486), .B(new_n452), .C1(new_n472), .C2(new_n474), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n479), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n470), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n236), .B1(new_n467), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n455), .B1(new_n464), .B2(KEYINPUT5), .ZN(new_n491));
  OR2_X1    g305(.A1(new_n471), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  XOR2_X1   g307(.A(new_n451), .B(KEYINPUT8), .Z(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(KEYINPUT7), .B1(new_n482), .B2(G953), .ZN(new_n497));
  OR2_X1    g311(.A1(new_n481), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n481), .A2(new_n497), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n496), .A2(new_n478), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n488), .A2(new_n500), .A3(new_n190), .ZN(new_n501));
  OAI21_X1  g315(.A(G210), .B1(G237), .B2(G902), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n488), .A2(new_n500), .A3(new_n190), .A4(new_n502), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n504), .A2(KEYINPUT90), .A3(new_n505), .ZN(new_n506));
  OR2_X1    g320(.A1(new_n505), .A2(KEYINPUT90), .ZN(new_n507));
  NAND2_X1  g321(.A1(G234), .A2(G237), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n508), .A2(G952), .A3(new_n288), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n508), .A2(G902), .A3(G953), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT21), .B(G898), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(G214), .B1(G237), .B2(G902), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n506), .A2(new_n507), .A3(new_n515), .A4(new_n516), .ZN(new_n517));
  OR3_X1    g331(.A1(new_n331), .A2(new_n450), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n442), .B1(G234), .B2(new_n190), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT82), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n521), .A2(KEYINPUT25), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT22), .B(G137), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n288), .A2(G221), .A3(G234), .ZN(new_n524));
  XOR2_X1   g338(.A(new_n523), .B(new_n524), .Z(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n385), .A2(new_n364), .ZN(new_n527));
  XNOR2_X1  g341(.A(KEYINPUT24), .B(G110), .ZN(new_n528));
  AOI21_X1  g342(.A(KEYINPUT77), .B1(new_n456), .B2(G128), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n456), .A2(KEYINPUT77), .A3(G128), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n456), .A2(G128), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n532), .A2(KEYINPUT78), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(KEYINPUT78), .B1(new_n532), .B2(new_n534), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n528), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n456), .A2(G128), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n538), .A2(KEYINPUT79), .A3(KEYINPUT23), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n539), .B(new_n533), .C1(KEYINPUT79), .C2(KEYINPUT23), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n540), .B1(new_n533), .B2(new_n539), .ZN(new_n541));
  INV_X1    g355(.A(G110), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n537), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT80), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT80), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n537), .A2(new_n546), .A3(new_n543), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n527), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n363), .A2(new_n364), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n549), .B1(new_n541), .B2(new_n542), .ZN(new_n550));
  NOR3_X1   g364(.A1(new_n535), .A2(new_n536), .A3(new_n528), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n526), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n552), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n537), .A2(new_n546), .A3(new_n543), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n546), .B1(new_n537), .B2(new_n543), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n554), .B(new_n525), .C1(new_n557), .C2(new_n527), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n522), .B1(new_n559), .B2(G902), .ZN(new_n560));
  INV_X1    g374(.A(new_n522), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n553), .A2(new_n558), .A3(new_n190), .A4(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n520), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n519), .A2(G902), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n553), .A2(new_n558), .A3(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(KEYINPUT83), .ZN(new_n566));
  OR2_X1    g380(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n473), .A2(KEYINPUT72), .A3(new_n470), .ZN(new_n569));
  AOI21_X1  g383(.A(KEYINPUT72), .B1(new_n473), .B2(new_n470), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n195), .A2(G134), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n200), .B1(new_n572), .B2(new_n197), .ZN(new_n573));
  OR2_X1    g387(.A1(new_n573), .A2(KEYINPUT67), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(KEYINPUT67), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(new_n201), .A3(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  AOI22_X1  g391(.A1(new_n279), .A2(new_n296), .B1(new_n265), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n202), .A2(new_n300), .A3(new_n301), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n579), .B1(new_n224), .B2(new_n576), .ZN(new_n580));
  AOI22_X1  g394(.A1(new_n571), .A2(new_n578), .B1(new_n476), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT28), .ZN(new_n582));
  OAI21_X1  g396(.A(KEYINPUT73), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n265), .A2(new_n577), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT72), .ZN(new_n585));
  AOI211_X1 g399(.A(new_n462), .B(new_n453), .C1(new_n459), .C2(new_n457), .ZN(new_n586));
  AOI21_X1  g400(.A(KEYINPUT70), .B1(new_n460), .B2(new_n454), .ZN(new_n587));
  NOR3_X1   g401(.A1(new_n586), .A2(new_n587), .A3(new_n469), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n585), .B1(new_n588), .B2(new_n489), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n247), .A2(new_n279), .A3(new_n248), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n473), .A2(KEYINPUT72), .A3(new_n470), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n584), .A2(new_n589), .A3(new_n590), .A4(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n580), .A2(new_n476), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT73), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(new_n595), .A3(KEYINPUT28), .ZN(new_n596));
  AOI21_X1  g410(.A(KEYINPUT28), .B1(new_n571), .B2(new_n578), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n583), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n344), .A2(new_n288), .A3(G210), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(KEYINPUT27), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT26), .B(G101), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n599), .A2(KEYINPUT74), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n584), .A2(KEYINPUT30), .A3(new_n590), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT30), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n580), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n606), .A2(new_n476), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n609), .A2(new_n603), .A3(new_n592), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT31), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n605), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(KEYINPUT74), .B1(new_n599), .B2(new_n604), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(G472), .A2(G902), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(KEYINPUT32), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n590), .B1(new_n224), .B2(new_n576), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n589), .A2(new_n591), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n620), .A2(KEYINPUT76), .A3(new_n592), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT76), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n618), .A2(new_n619), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n621), .A2(KEYINPUT28), .A3(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT29), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n597), .A2(new_n625), .A3(new_n604), .ZN(new_n626));
  AOI21_X1  g440(.A(G902), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n609), .A2(new_n592), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n604), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n625), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n597), .A2(new_n604), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n583), .A2(new_n632), .A3(new_n596), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n631), .B1(KEYINPUT75), .B2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT75), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n583), .A2(new_n632), .A3(new_n635), .A4(new_n596), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n628), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(G472), .ZN(new_n638));
  OAI22_X1  g452(.A1(new_n615), .A2(new_n617), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT74), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n595), .B1(new_n594), .B2(KEYINPUT28), .ZN(new_n641));
  AOI211_X1 g455(.A(KEYINPUT73), .B(new_n582), .C1(new_n592), .C2(new_n593), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n641), .A2(new_n642), .A3(new_n597), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n640), .B1(new_n643), .B2(new_n603), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n644), .A2(new_n612), .A3(new_n605), .ZN(new_n645));
  AOI21_X1  g459(.A(KEYINPUT32), .B1(new_n645), .B2(new_n616), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n568), .B1(new_n639), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(KEYINPUT84), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n616), .B1(new_n613), .B2(new_n614), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT32), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n617), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n645), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n633), .A2(KEYINPUT75), .ZN(new_n654));
  INV_X1    g468(.A(new_n631), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n654), .A2(new_n636), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n627), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(G472), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n651), .A2(new_n653), .A3(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT84), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n659), .A2(new_n660), .A3(new_n568), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n518), .B1(new_n648), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT96), .B(G101), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G3));
  NAND2_X1  g478(.A1(new_n645), .A2(new_n190), .ZN(new_n665));
  AOI22_X1  g479(.A1(new_n665), .A2(G472), .B1(new_n616), .B2(new_n645), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n666), .A2(new_n568), .A3(new_n330), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n516), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n669), .B1(new_n504), .B2(new_n505), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n515), .ZN(new_n671));
  AOI21_X1  g485(.A(KEYINPUT92), .B1(new_n411), .B2(new_n374), .ZN(new_n672));
  AOI211_X1 g486(.A(new_n407), .B(new_n373), .C1(new_n409), .C2(new_n410), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OAI211_X1 g488(.A(new_n447), .B(new_n190), .C1(new_n444), .C2(new_n445), .ZN(new_n675));
  NAND2_X1  g489(.A1(G478), .A2(G902), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g491(.A(KEYINPUT33), .B1(new_n444), .B2(new_n445), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n433), .A2(new_n441), .ZN(new_n679));
  INV_X1    g493(.A(new_n443), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT33), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n433), .A2(new_n441), .A3(new_n443), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n681), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n678), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n677), .B1(new_n685), .B2(G478), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n674), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(KEYINPUT97), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT97), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n674), .A2(new_n689), .A3(new_n686), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n671), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n668), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(KEYINPUT98), .ZN(new_n693));
  XOR2_X1   g507(.A(KEYINPUT34), .B(G104), .Z(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G6));
  NOR3_X1   g509(.A1(new_n671), .A2(new_n449), .A3(new_n406), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n668), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g511(.A(KEYINPUT35), .B(G107), .Z(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G9));
  NOR2_X1   g513(.A1(new_n548), .A2(new_n552), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n526), .A2(KEYINPUT36), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n700), .B(new_n702), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n703), .A2(new_n564), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n563), .A2(new_n704), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n517), .A2(new_n450), .A3(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n706), .A2(new_n666), .A3(new_n330), .ZN(new_n707));
  XOR2_X1   g521(.A(KEYINPUT37), .B(G110), .Z(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(KEYINPUT99), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(KEYINPUT100), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n707), .B(new_n710), .ZN(G12));
  OR2_X1    g525(.A1(new_n563), .A2(new_n704), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n712), .A2(new_n330), .A3(new_n670), .ZN(new_n713));
  INV_X1    g527(.A(new_n449), .ZN(new_n714));
  INV_X1    g528(.A(new_n406), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n509), .B1(new_n511), .B2(G900), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n659), .A2(new_n713), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G128), .ZN(G30));
  NAND2_X1  g534(.A1(new_n506), .A2(new_n507), .ZN(new_n721));
  XOR2_X1   g535(.A(new_n721), .B(KEYINPUT38), .Z(new_n722));
  NAND2_X1  g536(.A1(new_n674), .A2(new_n714), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  AND4_X1   g538(.A1(new_n516), .A2(new_n722), .A3(new_n705), .A4(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(KEYINPUT102), .B(KEYINPUT39), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n716), .B(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n330), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT40), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n729), .A2(KEYINPUT40), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n629), .A2(new_n603), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n621), .A2(new_n623), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n190), .B(new_n732), .C1(new_n733), .C2(new_n603), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(G472), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(KEYINPUT101), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n651), .A2(new_n736), .A3(new_n653), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n725), .A2(new_n730), .A3(new_n731), .A4(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n424), .ZN(G45));
  INV_X1    g553(.A(KEYINPUT103), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n674), .A2(new_n740), .A3(new_n686), .A4(new_n716), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n408), .A2(new_n686), .A3(new_n412), .A4(new_n716), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(KEYINPUT103), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(new_n659), .A3(new_n713), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G146), .ZN(G48));
  AOI22_X1  g561(.A1(G472), .A2(new_n657), .B1(new_n645), .B2(new_n652), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n567), .B1(new_n748), .B2(new_n651), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n286), .B1(new_n305), .B2(new_n307), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n310), .B1(new_n260), .B2(KEYINPUT88), .ZN(new_n751));
  AOI22_X1  g565(.A1(new_n750), .A2(new_n292), .B1(new_n751), .B2(new_n327), .ZN(new_n752));
  OAI21_X1  g566(.A(G469), .B1(new_n752), .B2(G902), .ZN(new_n753));
  INV_X1    g567(.A(new_n191), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(new_n754), .A3(new_n329), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(KEYINPUT104), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT104), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n753), .A2(new_n757), .A3(new_n329), .A4(new_n754), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n749), .A2(new_n691), .A3(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(KEYINPUT41), .B(G113), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n760), .B(new_n761), .ZN(G15));
  NAND4_X1  g576(.A1(new_n759), .A2(new_n659), .A3(new_n568), .A4(new_n696), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G116), .ZN(G18));
  AND4_X1   g578(.A1(new_n515), .A2(new_n756), .A3(new_n670), .A4(new_n758), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n413), .B(new_n449), .C1(new_n563), .C2(new_n704), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n766), .B1(new_n748), .B2(new_n651), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G119), .ZN(G21));
  AOI21_X1  g583(.A(new_n638), .B1(new_n645), .B2(new_n190), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n624), .A2(new_n598), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n604), .ZN(new_n772));
  AOI211_X1 g586(.A(G472), .B(G902), .C1(new_n772), .C2(new_n612), .ZN(new_n773));
  NOR4_X1   g587(.A1(new_n770), .A2(new_n567), .A3(new_n723), .A4(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n765), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G122), .ZN(G24));
  AND3_X1   g590(.A1(new_n756), .A2(new_n670), .A3(new_n758), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n770), .A2(new_n705), .A3(new_n773), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(new_n778), .A3(new_n745), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G125), .ZN(G27));
  INV_X1    g594(.A(KEYINPUT105), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n781), .A2(KEYINPUT42), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n669), .B1(new_n506), .B2(new_n507), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n741), .A2(new_n743), .A3(new_n783), .A4(new_n330), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n782), .B1(new_n647), .B2(new_n784), .ZN(new_n785));
  AND4_X1   g599(.A1(new_n330), .A2(new_n741), .A3(new_n743), .A4(new_n783), .ZN(new_n786));
  INV_X1    g600(.A(new_n782), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n749), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G131), .ZN(G33));
  INV_X1    g604(.A(new_n783), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(new_n331), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n717), .B(KEYINPUT106), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n749), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G134), .ZN(G36));
  INV_X1    g609(.A(new_n666), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n413), .A2(new_n686), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT43), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n796), .A2(new_n799), .A3(new_n712), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT44), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n802), .A2(new_n803), .A3(new_n791), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n293), .B1(new_n311), .B2(new_n313), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT45), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n317), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n807), .B1(new_n806), .B2(new_n805), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n808), .A2(KEYINPUT46), .A3(new_n315), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n315), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT46), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n809), .A2(new_n329), .A3(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n813), .A2(new_n754), .A3(new_n728), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(KEYINPUT107), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n804), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G137), .ZN(G39));
  AND2_X1   g631(.A1(new_n813), .A2(new_n754), .ZN(new_n818));
  OR2_X1    g632(.A1(new_n818), .A2(KEYINPUT47), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(KEYINPUT47), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NOR4_X1   g635(.A1(new_n659), .A2(new_n744), .A3(new_n568), .A4(new_n791), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(G140), .ZN(G42));
  NAND2_X1  g638(.A1(new_n799), .A2(new_n510), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n759), .A2(new_n783), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n825), .A2(new_n826), .A3(new_n647), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n827), .A2(KEYINPUT48), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n288), .A2(G952), .ZN(new_n829));
  NOR4_X1   g643(.A1(new_n826), .A2(new_n737), .A3(new_n567), .A4(new_n509), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n688), .A2(new_n690), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n770), .A2(new_n773), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n568), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n825), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n777), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n827), .A2(KEYINPUT48), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n828), .A2(new_n832), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n835), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(new_n722), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n759), .A2(new_n669), .ZN(new_n841));
  XOR2_X1   g655(.A(new_n841), .B(KEYINPUT111), .Z(new_n842));
  AND3_X1   g656(.A1(new_n840), .A2(new_n842), .A3(KEYINPUT50), .ZN(new_n843));
  AOI21_X1  g657(.A(KEYINPUT50), .B1(new_n840), .B2(new_n842), .ZN(new_n844));
  OR2_X1    g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n753), .A2(new_n329), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n819), .B(new_n820), .C1(new_n754), .C2(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n839), .A2(new_n791), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n845), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n674), .A2(new_n686), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n825), .A2(new_n826), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n830), .A2(new_n851), .B1(new_n778), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(KEYINPUT51), .B1(new_n853), .B2(KEYINPUT113), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n854), .B1(KEYINPUT113), .B2(new_n853), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n838), .B1(new_n850), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT112), .B1(new_n845), .B2(new_n853), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n853), .B(KEYINPUT112), .C1(new_n843), .C2(new_n844), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT110), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n849), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n847), .A2(KEYINPUT110), .A3(new_n848), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n858), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n856), .B1(new_n863), .B2(KEYINPUT51), .ZN(new_n864));
  INV_X1    g678(.A(new_n685), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n865), .A2(new_n447), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n408), .B(new_n412), .C1(new_n866), .C2(new_n677), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n450), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(new_n517), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n869), .A2(new_n666), .A3(new_n568), .A4(new_n330), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n775), .A2(new_n768), .A3(new_n763), .A4(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n760), .A2(new_n707), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n871), .A2(new_n662), .A3(new_n872), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n779), .A2(new_n719), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT52), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n716), .B(KEYINPUT109), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n331), .A2(new_n712), .A3(new_n876), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n724), .A2(new_n670), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n877), .A2(new_n737), .A3(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n874), .A2(new_n875), .A3(new_n746), .A4(new_n879), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n744), .A2(new_n770), .A3(new_n773), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n449), .A2(new_n715), .A3(new_n716), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n882), .B1(new_n748), .B2(new_n651), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n712), .B(new_n792), .C1(new_n881), .C2(new_n883), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n789), .A2(new_n794), .A3(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n879), .A2(new_n779), .A3(new_n719), .A4(new_n746), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(KEYINPUT52), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n873), .A2(new_n880), .A3(new_n885), .A4(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT53), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n874), .A2(new_n875), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n891), .A2(KEYINPUT53), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n890), .B1(new_n888), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(KEYINPUT54), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n789), .A2(new_n794), .A3(new_n884), .ZN(new_n895));
  NOR4_X1   g709(.A1(new_n895), .A2(new_n871), .A3(new_n662), .A4(new_n872), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n891), .A2(new_n889), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n896), .A2(new_n880), .A3(new_n887), .A4(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n890), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n894), .B1(KEYINPUT54), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n864), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(G952), .A2(G953), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT49), .ZN(new_n903));
  INV_X1    g717(.A(new_n846), .ZN(new_n904));
  AOI211_X1 g718(.A(new_n797), .B(new_n722), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n567), .A2(new_n191), .A3(new_n669), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT108), .ZN(new_n907));
  AOI22_X1  g721(.A1(new_n906), .A2(new_n907), .B1(new_n846), .B2(KEYINPUT49), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n905), .B(new_n908), .C1(new_n907), .C2(new_n906), .ZN(new_n909));
  OAI22_X1  g723(.A1(new_n901), .A2(new_n902), .B1(new_n737), .B2(new_n909), .ZN(G75));
  NOR2_X1   g724(.A1(new_n288), .A2(G952), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT115), .Z(new_n912));
  AND2_X1   g726(.A1(new_n888), .A2(new_n889), .ZN(new_n913));
  INV_X1    g727(.A(new_n897), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n888), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(G902), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT56), .B1(new_n917), .B2(G210), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n479), .A2(new_n487), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(new_n485), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT55), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n912), .B1(new_n918), .B2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT114), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n923), .B1(new_n899), .B2(G902), .ZN(new_n924));
  AOI211_X1 g738(.A(KEYINPUT114), .B(new_n190), .C1(new_n898), .C2(new_n890), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n503), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT56), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n921), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n922), .B1(new_n927), .B2(new_n929), .ZN(G51));
  NAND2_X1  g744(.A1(new_n916), .A2(KEYINPUT114), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n899), .A2(new_n923), .A3(G902), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n808), .B(KEYINPUT116), .Z(new_n933));
  NAND3_X1  g747(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n934), .A2(KEYINPUT117), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n315), .B(KEYINPUT57), .Z(new_n936));
  NOR2_X1   g750(.A1(new_n899), .A2(KEYINPUT54), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT54), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n938), .B1(new_n898), .B2(new_n890), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n936), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n752), .ZN(new_n941));
  AOI22_X1  g755(.A1(new_n934), .A2(KEYINPUT117), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n911), .B1(new_n935), .B2(new_n942), .ZN(G54));
  INV_X1    g757(.A(KEYINPUT118), .ZN(new_n944));
  AND2_X1   g758(.A1(KEYINPUT58), .A2(G475), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n404), .B1(new_n926), .B2(new_n945), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n404), .A2(new_n945), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n931), .A2(new_n932), .A3(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n911), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n944), .B1(new_n946), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n931), .A2(new_n932), .A3(new_n945), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n395), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n953), .A2(KEYINPUT118), .A3(new_n949), .A4(new_n948), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n951), .A2(new_n954), .ZN(G60));
  XNOR2_X1  g769(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(new_n676), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n865), .B(new_n957), .C1(new_n937), .C2(new_n939), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n912), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n865), .B1(new_n900), .B2(new_n957), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n959), .A2(new_n960), .ZN(G63));
  XNOR2_X1  g775(.A(new_n559), .B(KEYINPUT121), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n913), .A2(new_n915), .ZN(new_n963));
  NAND2_X1  g777(.A1(G217), .A2(G902), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT60), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n962), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  OR2_X1    g780(.A1(new_n963), .A2(new_n965), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n703), .B(KEYINPUT120), .Z(new_n968));
  OAI211_X1 g782(.A(new_n912), .B(new_n966), .C1(new_n967), .C2(new_n968), .ZN(new_n969));
  XNOR2_X1  g783(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(G66));
  OAI21_X1  g785(.A(G953), .B1(new_n513), .B2(new_n482), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n972), .B1(new_n873), .B2(G953), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n919), .B1(G898), .B2(new_n288), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n973), .B(new_n974), .ZN(G69));
  NAND2_X1  g789(.A1(new_n606), .A2(new_n608), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n380), .A2(new_n381), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n976), .B(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n874), .A2(new_n746), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n738), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT62), .ZN(new_n982));
  AOI22_X1  g796(.A1(new_n821), .A2(new_n822), .B1(new_n804), .B2(new_n815), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n648), .A2(new_n661), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n868), .B(KEYINPUT123), .Z(new_n985));
  NAND4_X1  g799(.A1(new_n984), .A2(new_n728), .A3(new_n792), .A4(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n983), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(KEYINPUT124), .B1(new_n982), .B2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT62), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n981), .B(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT124), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n990), .A2(new_n991), .A3(new_n983), .A4(new_n986), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n988), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n979), .B1(new_n993), .B2(G953), .ZN(new_n994));
  NAND2_X1  g808(.A1(G227), .A2(G900), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(G953), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n288), .A2(G900), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT125), .Z(new_n998));
  NAND3_X1  g812(.A1(new_n815), .A2(new_n749), .A3(new_n878), .ZN(new_n999));
  AND3_X1   g813(.A1(new_n980), .A2(new_n789), .A3(new_n794), .ZN(new_n1000));
  AND3_X1   g814(.A1(new_n983), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n998), .B1(new_n1001), .B2(G953), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(new_n978), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n994), .A2(new_n996), .A3(new_n1003), .ZN(new_n1004));
  OAI211_X1 g818(.A(G953), .B(new_n995), .C1(new_n1002), .C2(new_n979), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(G72));
  NAND3_X1  g820(.A1(new_n988), .A2(new_n992), .A3(new_n873), .ZN(new_n1007));
  NAND2_X1  g821(.A1(G472), .A2(G902), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT63), .Z(new_n1009));
  NAND2_X1  g823(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g824(.A(new_n732), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n609), .A2(new_n604), .A3(new_n592), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n893), .A2(new_n732), .A3(new_n1013), .A4(new_n1009), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n1014), .B(KEYINPUT127), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n983), .A2(new_n873), .A3(new_n999), .A4(new_n1000), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1013), .B1(new_n1016), .B2(new_n1009), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n1017), .A2(new_n911), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1018), .A2(KEYINPUT126), .ZN(new_n1019));
  AND2_X1   g833(.A1(new_n1018), .A2(KEYINPUT126), .ZN(new_n1020));
  OAI211_X1 g834(.A(new_n1012), .B(new_n1015), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  INV_X1    g835(.A(new_n1021), .ZN(G57));
endmodule


