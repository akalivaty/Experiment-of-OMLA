

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U554 ( .A1(G2104), .A2(G2105), .ZN(n524) );
  OR2_X1 U555 ( .A1(n724), .A2(n723), .ZN(n734) );
  NOR2_X1 U556 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U557 ( .A1(n933), .A2(n714), .ZN(n696) );
  AND2_X1 U558 ( .A1(n749), .A2(n748), .ZN(n751) );
  AND2_X1 U559 ( .A1(n520), .A2(n530), .ZN(G164) );
  NOR2_X1 U560 ( .A1(n538), .A2(n537), .ZN(G160) );
  NOR2_X2 U561 ( .A1(n769), .A2(n770), .ZN(n720) );
  XNOR2_X2 U562 ( .A(n521), .B(KEYINPUT66), .ZN(n893) );
  AND2_X1 U563 ( .A1(n523), .A2(n522), .ZN(n520) );
  INV_X1 U564 ( .A(KEYINPUT32), .ZN(n750) );
  XNOR2_X1 U565 ( .A(n751), .B(n750), .ZN(n752) );
  INV_X1 U566 ( .A(KEYINPUT100), .ZN(n757) );
  INV_X1 U567 ( .A(KEYINPUT88), .ZN(n528) );
  AND2_X1 U568 ( .A1(G2104), .A2(G2105), .ZN(n896) );
  NAND2_X1 U569 ( .A1(n896), .A2(G114), .ZN(n523) );
  INV_X1 U570 ( .A(G2105), .ZN(n525) );
  NOR2_X1 U571 ( .A1(n525), .A2(G2104), .ZN(n521) );
  NAND2_X1 U572 ( .A1(G126), .A2(n893), .ZN(n522) );
  XOR2_X2 U573 ( .A(KEYINPUT17), .B(n524), .Z(n887) );
  NAND2_X1 U574 ( .A1(G138), .A2(n887), .ZN(n527) );
  AND2_X2 U575 ( .A1(n525), .A2(G2104), .ZN(n889) );
  NAND2_X1 U576 ( .A1(G102), .A2(n889), .ZN(n526) );
  NAND2_X1 U577 ( .A1(n527), .A2(n526), .ZN(n529) );
  XNOR2_X1 U578 ( .A(n529), .B(n528), .ZN(n530) );
  NAND2_X1 U579 ( .A1(G101), .A2(n889), .ZN(n531) );
  XNOR2_X1 U580 ( .A(n531), .B(KEYINPUT67), .ZN(n532) );
  XNOR2_X1 U581 ( .A(n532), .B(KEYINPUT23), .ZN(n534) );
  NAND2_X1 U582 ( .A1(G137), .A2(n887), .ZN(n533) );
  NAND2_X1 U583 ( .A1(n534), .A2(n533), .ZN(n538) );
  NAND2_X1 U584 ( .A1(n896), .A2(G113), .ZN(n536) );
  NAND2_X1 U585 ( .A1(G125), .A2(n893), .ZN(n535) );
  NAND2_X1 U586 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U587 ( .A(G2430), .B(G2451), .Z(n540) );
  XNOR2_X1 U588 ( .A(KEYINPUT105), .B(G2443), .ZN(n539) );
  XNOR2_X1 U589 ( .A(n540), .B(n539), .ZN(n547) );
  XOR2_X1 U590 ( .A(G2435), .B(G2446), .Z(n542) );
  XNOR2_X1 U591 ( .A(G2427), .B(G2454), .ZN(n541) );
  XNOR2_X1 U592 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U593 ( .A(n543), .B(G2438), .Z(n545) );
  XNOR2_X1 U594 ( .A(G1348), .B(G1341), .ZN(n544) );
  XNOR2_X1 U595 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U596 ( .A(n547), .B(n546), .ZN(n548) );
  AND2_X1 U597 ( .A1(n548), .A2(G14), .ZN(G401) );
  INV_X1 U598 ( .A(G651), .ZN(n553) );
  NOR2_X1 U599 ( .A1(G543), .A2(n553), .ZN(n549) );
  XOR2_X1 U600 ( .A(KEYINPUT1), .B(n549), .Z(n661) );
  NAND2_X1 U601 ( .A1(G64), .A2(n661), .ZN(n552) );
  XOR2_X1 U602 ( .A(KEYINPUT0), .B(G543), .Z(n655) );
  NOR2_X1 U603 ( .A1(n655), .A2(G651), .ZN(n550) );
  XOR2_X2 U604 ( .A(KEYINPUT65), .B(n550), .Z(n657) );
  NAND2_X1 U605 ( .A1(G52), .A2(n657), .ZN(n551) );
  NAND2_X1 U606 ( .A1(n552), .A2(n551), .ZN(n558) );
  NOR2_X1 U607 ( .A1(n655), .A2(n553), .ZN(n649) );
  NAND2_X1 U608 ( .A1(G77), .A2(n649), .ZN(n555) );
  NOR2_X1 U609 ( .A1(G543), .A2(G651), .ZN(n646) );
  NAND2_X1 U610 ( .A1(G90), .A2(n646), .ZN(n554) );
  NAND2_X1 U611 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U612 ( .A(KEYINPUT9), .B(n556), .Z(n557) );
  NOR2_X1 U613 ( .A1(n558), .A2(n557), .ZN(G171) );
  AND2_X1 U614 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U615 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U616 ( .A(KEYINPUT76), .B(KEYINPUT6), .ZN(n562) );
  NAND2_X1 U617 ( .A1(G63), .A2(n661), .ZN(n560) );
  NAND2_X1 U618 ( .A1(G51), .A2(n657), .ZN(n559) );
  NAND2_X1 U619 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U620 ( .A(n562), .B(n561), .ZN(n570) );
  NAND2_X1 U621 ( .A1(G89), .A2(n646), .ZN(n563) );
  XNOR2_X1 U622 ( .A(n563), .B(KEYINPUT74), .ZN(n564) );
  XNOR2_X1 U623 ( .A(n564), .B(KEYINPUT4), .ZN(n566) );
  NAND2_X1 U624 ( .A1(G76), .A2(n649), .ZN(n565) );
  NAND2_X1 U625 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U626 ( .A(KEYINPUT5), .B(n567), .ZN(n568) );
  XNOR2_X1 U627 ( .A(KEYINPUT75), .B(n568), .ZN(n569) );
  NOR2_X1 U628 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U629 ( .A(KEYINPUT7), .B(n571), .Z(G168) );
  XNOR2_X1 U630 ( .A(G168), .B(KEYINPUT8), .ZN(n572) );
  XNOR2_X1 U631 ( .A(n572), .B(KEYINPUT77), .ZN(G286) );
  NAND2_X1 U632 ( .A1(G7), .A2(G661), .ZN(n573) );
  XNOR2_X1 U633 ( .A(n573), .B(KEYINPUT70), .ZN(n574) );
  XNOR2_X1 U634 ( .A(KEYINPUT10), .B(n574), .ZN(G223) );
  INV_X1 U635 ( .A(G223), .ZN(n839) );
  NAND2_X1 U636 ( .A1(n839), .A2(G567), .ZN(n575) );
  XOR2_X1 U637 ( .A(KEYINPUT11), .B(n575), .Z(G234) );
  NAND2_X1 U638 ( .A1(n646), .A2(G81), .ZN(n576) );
  XNOR2_X1 U639 ( .A(KEYINPUT12), .B(n576), .ZN(n579) );
  NAND2_X1 U640 ( .A1(n649), .A2(G68), .ZN(n577) );
  XOR2_X1 U641 ( .A(KEYINPUT71), .B(n577), .Z(n578) );
  NAND2_X1 U642 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U643 ( .A(n580), .B(KEYINPUT13), .ZN(n582) );
  NAND2_X1 U644 ( .A1(G43), .A2(n657), .ZN(n581) );
  NAND2_X1 U645 ( .A1(n582), .A2(n581), .ZN(n585) );
  NAND2_X1 U646 ( .A1(n661), .A2(G56), .ZN(n583) );
  XOR2_X1 U647 ( .A(KEYINPUT14), .B(n583), .Z(n584) );
  NOR2_X1 U648 ( .A1(n585), .A2(n584), .ZN(n935) );
  NAND2_X1 U649 ( .A1(n935), .A2(G860), .ZN(G153) );
  XOR2_X1 U650 ( .A(G171), .B(KEYINPUT72), .Z(G301) );
  NAND2_X1 U651 ( .A1(G868), .A2(G301), .ZN(n595) );
  NAND2_X1 U652 ( .A1(G66), .A2(n661), .ZN(n587) );
  NAND2_X1 U653 ( .A1(G79), .A2(n649), .ZN(n586) );
  NAND2_X1 U654 ( .A1(n587), .A2(n586), .ZN(n591) );
  NAND2_X1 U655 ( .A1(G92), .A2(n646), .ZN(n589) );
  NAND2_X1 U656 ( .A1(G54), .A2(n657), .ZN(n588) );
  NAND2_X1 U657 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U658 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U659 ( .A(KEYINPUT15), .B(n592), .Z(n593) );
  XNOR2_X1 U660 ( .A(KEYINPUT73), .B(n593), .ZN(n930) );
  INV_X1 U661 ( .A(G868), .ZN(n674) );
  NAND2_X1 U662 ( .A1(n930), .A2(n674), .ZN(n594) );
  NAND2_X1 U663 ( .A1(n595), .A2(n594), .ZN(G284) );
  NAND2_X1 U664 ( .A1(G65), .A2(n661), .ZN(n597) );
  NAND2_X1 U665 ( .A1(G91), .A2(n646), .ZN(n596) );
  NAND2_X1 U666 ( .A1(n597), .A2(n596), .ZN(n600) );
  NAND2_X1 U667 ( .A1(G78), .A2(n649), .ZN(n598) );
  XNOR2_X1 U668 ( .A(KEYINPUT69), .B(n598), .ZN(n599) );
  NOR2_X1 U669 ( .A1(n600), .A2(n599), .ZN(n602) );
  NAND2_X1 U670 ( .A1(n657), .A2(G53), .ZN(n601) );
  NAND2_X1 U671 ( .A1(n602), .A2(n601), .ZN(G299) );
  NOR2_X1 U672 ( .A1(G286), .A2(n674), .ZN(n604) );
  NOR2_X1 U673 ( .A1(G868), .A2(G299), .ZN(n603) );
  NOR2_X1 U674 ( .A1(n604), .A2(n603), .ZN(G297) );
  INV_X1 U675 ( .A(G860), .ZN(n624) );
  NAND2_X1 U676 ( .A1(n624), .A2(G559), .ZN(n605) );
  INV_X1 U677 ( .A(n930), .ZN(n847) );
  NAND2_X1 U678 ( .A1(n605), .A2(n847), .ZN(n606) );
  XNOR2_X1 U679 ( .A(n606), .B(KEYINPUT78), .ZN(n607) );
  XNOR2_X1 U680 ( .A(KEYINPUT16), .B(n607), .ZN(G148) );
  NAND2_X1 U681 ( .A1(n847), .A2(G868), .ZN(n608) );
  NOR2_X1 U682 ( .A1(G559), .A2(n608), .ZN(n610) );
  AND2_X1 U683 ( .A1(n674), .A2(n935), .ZN(n609) );
  NOR2_X1 U684 ( .A1(n610), .A2(n609), .ZN(G282) );
  NAND2_X1 U685 ( .A1(n893), .A2(G123), .ZN(n611) );
  XNOR2_X1 U686 ( .A(n611), .B(KEYINPUT18), .ZN(n618) );
  NAND2_X1 U687 ( .A1(G135), .A2(n887), .ZN(n613) );
  NAND2_X1 U688 ( .A1(G111), .A2(n896), .ZN(n612) );
  NAND2_X1 U689 ( .A1(n613), .A2(n612), .ZN(n616) );
  NAND2_X1 U690 ( .A1(G99), .A2(n889), .ZN(n614) );
  XNOR2_X1 U691 ( .A(KEYINPUT79), .B(n614), .ZN(n615) );
  NOR2_X1 U692 ( .A1(n616), .A2(n615), .ZN(n617) );
  NAND2_X1 U693 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U694 ( .A(KEYINPUT80), .B(n619), .ZN(n980) );
  XNOR2_X1 U695 ( .A(n980), .B(G2096), .ZN(n620) );
  XNOR2_X1 U696 ( .A(n620), .B(KEYINPUT81), .ZN(n622) );
  INV_X1 U697 ( .A(G2100), .ZN(n621) );
  NAND2_X1 U698 ( .A1(n622), .A2(n621), .ZN(G156) );
  NAND2_X1 U699 ( .A1(G559), .A2(n847), .ZN(n623) );
  XNOR2_X1 U700 ( .A(n623), .B(n935), .ZN(n670) );
  NAND2_X1 U701 ( .A1(n624), .A2(n670), .ZN(n631) );
  NAND2_X1 U702 ( .A1(G67), .A2(n661), .ZN(n626) );
  NAND2_X1 U703 ( .A1(G55), .A2(n657), .ZN(n625) );
  NAND2_X1 U704 ( .A1(n626), .A2(n625), .ZN(n630) );
  NAND2_X1 U705 ( .A1(G80), .A2(n649), .ZN(n628) );
  NAND2_X1 U706 ( .A1(G93), .A2(n646), .ZN(n627) );
  NAND2_X1 U707 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n673) );
  XOR2_X1 U709 ( .A(n631), .B(n673), .Z(G145) );
  NAND2_X1 U710 ( .A1(G62), .A2(n661), .ZN(n633) );
  NAND2_X1 U711 ( .A1(G75), .A2(n649), .ZN(n632) );
  NAND2_X1 U712 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U713 ( .A1(n646), .A2(G88), .ZN(n634) );
  XOR2_X1 U714 ( .A(KEYINPUT84), .B(n634), .Z(n635) );
  NOR2_X1 U715 ( .A1(n636), .A2(n635), .ZN(n638) );
  NAND2_X1 U716 ( .A1(n657), .A2(G50), .ZN(n637) );
  NAND2_X1 U717 ( .A1(n638), .A2(n637), .ZN(G303) );
  INV_X1 U718 ( .A(G303), .ZN(G166) );
  NAND2_X1 U719 ( .A1(n649), .A2(G72), .ZN(n640) );
  NAND2_X1 U720 ( .A1(n661), .A2(G60), .ZN(n639) );
  NAND2_X1 U721 ( .A1(n640), .A2(n639), .ZN(n644) );
  NAND2_X1 U722 ( .A1(G85), .A2(n646), .ZN(n642) );
  NAND2_X1 U723 ( .A1(G47), .A2(n657), .ZN(n641) );
  NAND2_X1 U724 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U725 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U726 ( .A(KEYINPUT68), .B(n645), .Z(G290) );
  NAND2_X1 U727 ( .A1(G61), .A2(n661), .ZN(n648) );
  NAND2_X1 U728 ( .A1(G86), .A2(n646), .ZN(n647) );
  NAND2_X1 U729 ( .A1(n648), .A2(n647), .ZN(n652) );
  NAND2_X1 U730 ( .A1(n649), .A2(G73), .ZN(n650) );
  XOR2_X1 U731 ( .A(KEYINPUT2), .B(n650), .Z(n651) );
  NOR2_X1 U732 ( .A1(n652), .A2(n651), .ZN(n654) );
  NAND2_X1 U733 ( .A1(n657), .A2(G48), .ZN(n653) );
  NAND2_X1 U734 ( .A1(n654), .A2(n653), .ZN(G305) );
  NAND2_X1 U735 ( .A1(G87), .A2(n655), .ZN(n656) );
  XNOR2_X1 U736 ( .A(n656), .B(KEYINPUT82), .ZN(n663) );
  NAND2_X1 U737 ( .A1(G49), .A2(n657), .ZN(n659) );
  NAND2_X1 U738 ( .A1(G74), .A2(G651), .ZN(n658) );
  NAND2_X1 U739 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U740 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U741 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U742 ( .A(KEYINPUT83), .B(n664), .Z(G288) );
  XNOR2_X1 U743 ( .A(G166), .B(KEYINPUT19), .ZN(n669) );
  INV_X1 U744 ( .A(G299), .ZN(n933) );
  XNOR2_X1 U745 ( .A(n933), .B(n673), .ZN(n667) );
  XNOR2_X1 U746 ( .A(G290), .B(G305), .ZN(n665) );
  XNOR2_X1 U747 ( .A(n665), .B(G288), .ZN(n666) );
  XNOR2_X1 U748 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U749 ( .A(n669), .B(n668), .ZN(n846) );
  XNOR2_X1 U750 ( .A(n670), .B(n846), .ZN(n671) );
  XNOR2_X1 U751 ( .A(KEYINPUT85), .B(n671), .ZN(n672) );
  NOR2_X1 U752 ( .A1(n674), .A2(n672), .ZN(n676) );
  AND2_X1 U753 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U754 ( .A1(n676), .A2(n675), .ZN(G295) );
  NAND2_X1 U755 ( .A1(G2078), .A2(G2084), .ZN(n677) );
  XOR2_X1 U756 ( .A(KEYINPUT20), .B(n677), .Z(n678) );
  NAND2_X1 U757 ( .A1(G2090), .A2(n678), .ZN(n679) );
  XNOR2_X1 U758 ( .A(KEYINPUT21), .B(n679), .ZN(n680) );
  NAND2_X1 U759 ( .A1(n680), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U760 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U761 ( .A(KEYINPUT86), .B(KEYINPUT22), .Z(n682) );
  NAND2_X1 U762 ( .A1(G132), .A2(G82), .ZN(n681) );
  XNOR2_X1 U763 ( .A(n682), .B(n681), .ZN(n683) );
  NAND2_X1 U764 ( .A1(n683), .A2(G96), .ZN(n684) );
  NOR2_X1 U765 ( .A1(n684), .A2(G218), .ZN(n685) );
  XNOR2_X1 U766 ( .A(n685), .B(KEYINPUT87), .ZN(n844) );
  NAND2_X1 U767 ( .A1(n844), .A2(G2106), .ZN(n689) );
  NAND2_X1 U768 ( .A1(G108), .A2(G120), .ZN(n686) );
  NOR2_X1 U769 ( .A1(G237), .A2(n686), .ZN(n687) );
  NAND2_X1 U770 ( .A1(G69), .A2(n687), .ZN(n845) );
  NAND2_X1 U771 ( .A1(n845), .A2(G567), .ZN(n688) );
  NAND2_X1 U772 ( .A1(n689), .A2(n688), .ZN(n919) );
  NAND2_X1 U773 ( .A1(G483), .A2(G661), .ZN(n690) );
  NOR2_X1 U774 ( .A1(n919), .A2(n690), .ZN(n841) );
  NAND2_X1 U775 ( .A1(n841), .A2(G36), .ZN(G176) );
  NOR2_X1 U776 ( .A1(G164), .A2(G1384), .ZN(n691) );
  INV_X1 U777 ( .A(n691), .ZN(n769) );
  NAND2_X1 U778 ( .A1(G160), .A2(G40), .ZN(n770) );
  INV_X1 U779 ( .A(n720), .ZN(n697) );
  NAND2_X1 U780 ( .A1(n697), .A2(G8), .ZN(n814) );
  NOR2_X1 U781 ( .A1(G1966), .A2(n814), .ZN(n738) );
  INV_X1 U782 ( .A(n720), .ZN(n740) );
  NAND2_X1 U783 ( .A1(G1956), .A2(n740), .ZN(n694) );
  NAND2_X1 U784 ( .A1(n720), .A2(G2072), .ZN(n692) );
  XOR2_X1 U785 ( .A(n692), .B(KEYINPUT27), .Z(n693) );
  NAND2_X1 U786 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U787 ( .A(n695), .B(KEYINPUT94), .Z(n714) );
  XOR2_X1 U788 ( .A(n696), .B(KEYINPUT28), .Z(n718) );
  NAND2_X1 U789 ( .A1(G1348), .A2(n697), .ZN(n699) );
  NAND2_X1 U790 ( .A1(G2067), .A2(n720), .ZN(n698) );
  NAND2_X1 U791 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U792 ( .A(n700), .B(KEYINPUT95), .ZN(n701) );
  AND2_X1 U793 ( .A1(n847), .A2(n701), .ZN(n713) );
  XNOR2_X1 U794 ( .A(KEYINPUT64), .B(KEYINPUT26), .ZN(n703) );
  NOR2_X1 U795 ( .A1(G1996), .A2(n703), .ZN(n711) );
  NOR2_X1 U796 ( .A1(n847), .A2(n701), .ZN(n708) );
  INV_X1 U797 ( .A(G1341), .ZN(n959) );
  NAND2_X1 U798 ( .A1(n959), .A2(n703), .ZN(n702) );
  NAND2_X1 U799 ( .A1(n702), .A2(n740), .ZN(n706) );
  INV_X1 U800 ( .A(G1996), .ZN(n1011) );
  NOR2_X1 U801 ( .A1(n1011), .A2(n740), .ZN(n704) );
  NAND2_X1 U802 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U803 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U804 ( .A1(n935), .A2(n709), .ZN(n710) );
  NOR2_X1 U805 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U806 ( .A1(n713), .A2(n712), .ZN(n716) );
  NAND2_X1 U807 ( .A1(n933), .A2(n714), .ZN(n715) );
  NAND2_X1 U808 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U809 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U810 ( .A(n719), .B(KEYINPUT29), .ZN(n724) );
  INV_X1 U811 ( .A(G1961), .ZN(n948) );
  NAND2_X1 U812 ( .A1(n740), .A2(n948), .ZN(n722) );
  XNOR2_X1 U813 ( .A(G2078), .B(KEYINPUT25), .ZN(n1010) );
  NAND2_X1 U814 ( .A1(n720), .A2(n1010), .ZN(n721) );
  NAND2_X1 U815 ( .A1(n722), .A2(n721), .ZN(n729) );
  AND2_X1 U816 ( .A1(n729), .A2(G171), .ZN(n723) );
  NOR2_X1 U817 ( .A1(G2084), .A2(n740), .ZN(n735) );
  NOR2_X1 U818 ( .A1(n738), .A2(n735), .ZN(n725) );
  NAND2_X1 U819 ( .A1(G8), .A2(n725), .ZN(n726) );
  XNOR2_X1 U820 ( .A(KEYINPUT96), .B(n726), .ZN(n727) );
  XNOR2_X1 U821 ( .A(KEYINPUT30), .B(n727), .ZN(n728) );
  NOR2_X1 U822 ( .A1(G168), .A2(n728), .ZN(n731) );
  NOR2_X1 U823 ( .A1(G171), .A2(n729), .ZN(n730) );
  NOR2_X1 U824 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U825 ( .A(KEYINPUT31), .B(n732), .Z(n733) );
  NAND2_X1 U826 ( .A1(n734), .A2(n733), .ZN(n739) );
  NAND2_X1 U827 ( .A1(G8), .A2(n735), .ZN(n736) );
  NAND2_X1 U828 ( .A1(n739), .A2(n736), .ZN(n737) );
  NOR2_X1 U829 ( .A1(n738), .A2(n737), .ZN(n753) );
  NAND2_X1 U830 ( .A1(n739), .A2(G286), .ZN(n749) );
  INV_X1 U831 ( .A(G8), .ZN(n747) );
  NOR2_X1 U832 ( .A1(G2090), .A2(n740), .ZN(n741) );
  XNOR2_X1 U833 ( .A(KEYINPUT97), .B(n741), .ZN(n744) );
  NOR2_X1 U834 ( .A1(G1971), .A2(n814), .ZN(n742) );
  NOR2_X1 U835 ( .A1(G166), .A2(n742), .ZN(n743) );
  NAND2_X1 U836 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U837 ( .A(n745), .B(KEYINPUT98), .ZN(n746) );
  OR2_X1 U838 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U839 ( .A1(n753), .A2(n752), .ZN(n806) );
  NOR2_X1 U840 ( .A1(G1971), .A2(G303), .ZN(n754) );
  NOR2_X1 U841 ( .A1(n806), .A2(n754), .ZN(n756) );
  NOR2_X1 U842 ( .A1(G1976), .A2(G288), .ZN(n755) );
  XNOR2_X1 U843 ( .A(KEYINPUT99), .B(n755), .ZN(n924) );
  NAND2_X1 U844 ( .A1(n756), .A2(n924), .ZN(n758) );
  XNOR2_X1 U845 ( .A(n758), .B(n757), .ZN(n759) );
  NOR2_X1 U846 ( .A1(n814), .A2(n759), .ZN(n763) );
  NAND2_X1 U847 ( .A1(G1976), .A2(G288), .ZN(n925) );
  INV_X1 U848 ( .A(KEYINPUT33), .ZN(n765) );
  OR2_X1 U849 ( .A1(n814), .A2(n924), .ZN(n760) );
  NOR2_X1 U850 ( .A1(n765), .A2(n760), .ZN(n761) );
  XNOR2_X1 U851 ( .A(n761), .B(KEYINPUT101), .ZN(n764) );
  AND2_X1 U852 ( .A1(n925), .A2(n764), .ZN(n762) );
  NAND2_X1 U853 ( .A1(n763), .A2(n762), .ZN(n768) );
  INV_X1 U854 ( .A(n764), .ZN(n766) );
  OR2_X1 U855 ( .A1(n766), .A2(n765), .ZN(n767) );
  AND2_X1 U856 ( .A1(n768), .A2(n767), .ZN(n804) );
  XNOR2_X1 U857 ( .A(G1981), .B(G305), .ZN(n921) );
  XNOR2_X1 U858 ( .A(G1986), .B(G290), .ZN(n932) );
  NOR2_X1 U859 ( .A1(n691), .A2(n770), .ZN(n834) );
  AND2_X1 U860 ( .A1(n932), .A2(n834), .ZN(n802) );
  XNOR2_X1 U861 ( .A(KEYINPUT37), .B(G2067), .ZN(n823) );
  NAND2_X1 U862 ( .A1(G140), .A2(n887), .ZN(n772) );
  NAND2_X1 U863 ( .A1(G104), .A2(n889), .ZN(n771) );
  NAND2_X1 U864 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U865 ( .A(KEYINPUT34), .B(n773), .ZN(n778) );
  NAND2_X1 U866 ( .A1(n896), .A2(G116), .ZN(n775) );
  NAND2_X1 U867 ( .A1(G128), .A2(n893), .ZN(n774) );
  NAND2_X1 U868 ( .A1(n775), .A2(n774), .ZN(n776) );
  XOR2_X1 U869 ( .A(KEYINPUT35), .B(n776), .Z(n777) );
  NOR2_X1 U870 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U871 ( .A(KEYINPUT36), .B(n779), .ZN(n902) );
  NOR2_X1 U872 ( .A1(n823), .A2(n902), .ZN(n991) );
  NAND2_X1 U873 ( .A1(n834), .A2(n991), .ZN(n831) );
  NAND2_X1 U874 ( .A1(n889), .A2(G95), .ZN(n780) );
  XOR2_X1 U875 ( .A(KEYINPUT89), .B(n780), .Z(n782) );
  NAND2_X1 U876 ( .A1(n887), .A2(G131), .ZN(n781) );
  NAND2_X1 U877 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U878 ( .A(KEYINPUT90), .B(n783), .ZN(n787) );
  NAND2_X1 U879 ( .A1(n896), .A2(G107), .ZN(n785) );
  NAND2_X1 U880 ( .A1(G119), .A2(n893), .ZN(n784) );
  NAND2_X1 U881 ( .A1(n785), .A2(n784), .ZN(n786) );
  NOR2_X1 U882 ( .A1(n787), .A2(n786), .ZN(n886) );
  INV_X1 U883 ( .A(G1991), .ZN(n1008) );
  NOR2_X1 U884 ( .A1(n886), .A2(n1008), .ZN(n797) );
  NAND2_X1 U885 ( .A1(G141), .A2(n887), .ZN(n789) );
  NAND2_X1 U886 ( .A1(G129), .A2(n893), .ZN(n788) );
  NAND2_X1 U887 ( .A1(n789), .A2(n788), .ZN(n793) );
  NAND2_X1 U888 ( .A1(G105), .A2(n889), .ZN(n790) );
  XNOR2_X1 U889 ( .A(n790), .B(KEYINPUT91), .ZN(n791) );
  XNOR2_X1 U890 ( .A(n791), .B(KEYINPUT38), .ZN(n792) );
  NOR2_X1 U891 ( .A1(n793), .A2(n792), .ZN(n795) );
  NAND2_X1 U892 ( .A1(n896), .A2(G117), .ZN(n794) );
  NAND2_X1 U893 ( .A1(n795), .A2(n794), .ZN(n904) );
  AND2_X1 U894 ( .A1(n904), .A2(G1996), .ZN(n796) );
  NOR2_X1 U895 ( .A1(n797), .A2(n796), .ZN(n989) );
  INV_X1 U896 ( .A(n834), .ZN(n798) );
  NOR2_X1 U897 ( .A1(n989), .A2(n798), .ZN(n826) );
  INV_X1 U898 ( .A(n826), .ZN(n799) );
  NAND2_X1 U899 ( .A1(n831), .A2(n799), .ZN(n800) );
  XNOR2_X1 U900 ( .A(KEYINPUT92), .B(n800), .ZN(n801) );
  OR2_X1 U901 ( .A1(n802), .A2(n801), .ZN(n805) );
  OR2_X1 U902 ( .A1(n921), .A2(n805), .ZN(n803) );
  NOR2_X1 U903 ( .A1(n804), .A2(n803), .ZN(n822) );
  INV_X1 U904 ( .A(n805), .ZN(n820) );
  INV_X1 U905 ( .A(n806), .ZN(n809) );
  NOR2_X1 U906 ( .A1(G2090), .A2(G303), .ZN(n807) );
  NAND2_X1 U907 ( .A1(G8), .A2(n807), .ZN(n808) );
  NAND2_X1 U908 ( .A1(n809), .A2(n808), .ZN(n810) );
  XNOR2_X1 U909 ( .A(n810), .B(KEYINPUT102), .ZN(n811) );
  NAND2_X1 U910 ( .A1(n811), .A2(n814), .ZN(n818) );
  NOR2_X1 U911 ( .A1(G1981), .A2(G305), .ZN(n812) );
  XOR2_X1 U912 ( .A(n812), .B(KEYINPUT93), .Z(n813) );
  XNOR2_X1 U913 ( .A(KEYINPUT24), .B(n813), .ZN(n816) );
  INV_X1 U914 ( .A(n814), .ZN(n815) );
  NAND2_X1 U915 ( .A1(n816), .A2(n815), .ZN(n817) );
  NAND2_X1 U916 ( .A1(n818), .A2(n817), .ZN(n819) );
  AND2_X1 U917 ( .A1(n820), .A2(n819), .ZN(n821) );
  NOR2_X1 U918 ( .A1(n822), .A2(n821), .ZN(n837) );
  NAND2_X1 U919 ( .A1(n823), .A2(n902), .ZN(n993) );
  NOR2_X1 U920 ( .A1(G1996), .A2(n904), .ZN(n982) );
  NOR2_X1 U921 ( .A1(G1986), .A2(G290), .ZN(n824) );
  AND2_X1 U922 ( .A1(n1008), .A2(n886), .ZN(n978) );
  NOR2_X1 U923 ( .A1(n824), .A2(n978), .ZN(n825) );
  NOR2_X1 U924 ( .A1(n826), .A2(n825), .ZN(n827) );
  XOR2_X1 U925 ( .A(KEYINPUT103), .B(n827), .Z(n828) );
  NOR2_X1 U926 ( .A1(n982), .A2(n828), .ZN(n829) );
  XNOR2_X1 U927 ( .A(KEYINPUT104), .B(n829), .ZN(n830) );
  XNOR2_X1 U928 ( .A(n830), .B(KEYINPUT39), .ZN(n832) );
  NAND2_X1 U929 ( .A1(n832), .A2(n831), .ZN(n833) );
  NAND2_X1 U930 ( .A1(n993), .A2(n833), .ZN(n835) );
  NAND2_X1 U931 ( .A1(n835), .A2(n834), .ZN(n836) );
  NAND2_X1 U932 ( .A1(n837), .A2(n836), .ZN(n838) );
  XNOR2_X1 U933 ( .A(n838), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U934 ( .A1(G2106), .A2(n839), .ZN(G217) );
  AND2_X1 U935 ( .A1(G15), .A2(G2), .ZN(n840) );
  NAND2_X1 U936 ( .A1(G661), .A2(n840), .ZN(G259) );
  NAND2_X1 U937 ( .A1(G1), .A2(G3), .ZN(n842) );
  NAND2_X1 U938 ( .A1(n842), .A2(n841), .ZN(n843) );
  XNOR2_X1 U939 ( .A(n843), .B(KEYINPUT106), .ZN(G188) );
  XNOR2_X1 U940 ( .A(G120), .B(KEYINPUT107), .ZN(G236) );
  INV_X1 U942 ( .A(G132), .ZN(G219) );
  INV_X1 U943 ( .A(G108), .ZN(G238) );
  INV_X1 U944 ( .A(G96), .ZN(G221) );
  INV_X1 U945 ( .A(G82), .ZN(G220) );
  NOR2_X1 U946 ( .A1(n845), .A2(n844), .ZN(G325) );
  INV_X1 U947 ( .A(G325), .ZN(G261) );
  XOR2_X1 U948 ( .A(n846), .B(G286), .Z(n849) );
  XNOR2_X1 U949 ( .A(G171), .B(n847), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U951 ( .A(n935), .B(n850), .Z(n851) );
  NOR2_X1 U952 ( .A1(G37), .A2(n851), .ZN(G397) );
  XOR2_X1 U953 ( .A(G2100), .B(G2096), .Z(n853) );
  XNOR2_X1 U954 ( .A(KEYINPUT42), .B(G2678), .ZN(n852) );
  XNOR2_X1 U955 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U956 ( .A(KEYINPUT43), .B(G2090), .Z(n855) );
  XNOR2_X1 U957 ( .A(G2067), .B(G2072), .ZN(n854) );
  XNOR2_X1 U958 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U959 ( .A(n857), .B(n856), .Z(n859) );
  XNOR2_X1 U960 ( .A(G2078), .B(G2084), .ZN(n858) );
  XNOR2_X1 U961 ( .A(n859), .B(n858), .ZN(G227) );
  XOR2_X1 U962 ( .A(KEYINPUT41), .B(G1961), .Z(n861) );
  XNOR2_X1 U963 ( .A(G1996), .B(G1991), .ZN(n860) );
  XNOR2_X1 U964 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U965 ( .A(n862), .B(G2474), .Z(n864) );
  XNOR2_X1 U966 ( .A(G1956), .B(G1976), .ZN(n863) );
  XNOR2_X1 U967 ( .A(n864), .B(n863), .ZN(n868) );
  XOR2_X1 U968 ( .A(G1981), .B(G1971), .Z(n866) );
  XNOR2_X1 U969 ( .A(G1986), .B(G1966), .ZN(n865) );
  XNOR2_X1 U970 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U971 ( .A(n868), .B(n867), .Z(n870) );
  XNOR2_X1 U972 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n869) );
  XNOR2_X1 U973 ( .A(n870), .B(n869), .ZN(G229) );
  NAND2_X1 U974 ( .A1(G100), .A2(n889), .ZN(n872) );
  NAND2_X1 U975 ( .A1(G112), .A2(n896), .ZN(n871) );
  NAND2_X1 U976 ( .A1(n872), .A2(n871), .ZN(n877) );
  NAND2_X1 U977 ( .A1(n893), .A2(G124), .ZN(n873) );
  XNOR2_X1 U978 ( .A(n873), .B(KEYINPUT44), .ZN(n875) );
  NAND2_X1 U979 ( .A1(n887), .A2(G136), .ZN(n874) );
  NAND2_X1 U980 ( .A1(n875), .A2(n874), .ZN(n876) );
  NOR2_X1 U981 ( .A1(n877), .A2(n876), .ZN(G162) );
  NAND2_X1 U982 ( .A1(G139), .A2(n887), .ZN(n879) );
  NAND2_X1 U983 ( .A1(G103), .A2(n889), .ZN(n878) );
  NAND2_X1 U984 ( .A1(n879), .A2(n878), .ZN(n885) );
  NAND2_X1 U985 ( .A1(n896), .A2(G115), .ZN(n880) );
  XNOR2_X1 U986 ( .A(n880), .B(KEYINPUT112), .ZN(n882) );
  NAND2_X1 U987 ( .A1(G127), .A2(n893), .ZN(n881) );
  NAND2_X1 U988 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U989 ( .A(KEYINPUT47), .B(n883), .Z(n884) );
  NOR2_X1 U990 ( .A1(n885), .A2(n884), .ZN(n996) );
  XNOR2_X1 U991 ( .A(n886), .B(n996), .ZN(n911) );
  NAND2_X1 U992 ( .A1(n887), .A2(G142), .ZN(n888) );
  XOR2_X1 U993 ( .A(KEYINPUT111), .B(n888), .Z(n891) );
  NAND2_X1 U994 ( .A1(n889), .A2(G106), .ZN(n890) );
  NAND2_X1 U995 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U996 ( .A(n892), .B(KEYINPUT45), .ZN(n895) );
  NAND2_X1 U997 ( .A1(G130), .A2(n893), .ZN(n894) );
  NAND2_X1 U998 ( .A1(n895), .A2(n894), .ZN(n899) );
  NAND2_X1 U999 ( .A1(n896), .A2(G118), .ZN(n897) );
  XOR2_X1 U1000 ( .A(KEYINPUT110), .B(n897), .Z(n898) );
  NOR2_X1 U1001 ( .A1(n899), .A2(n898), .ZN(n909) );
  XOR2_X1 U1002 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n901) );
  XNOR2_X1 U1003 ( .A(G164), .B(G160), .ZN(n900) );
  XNOR2_X1 U1004 ( .A(n901), .B(n900), .ZN(n903) );
  XNOR2_X1 U1005 ( .A(n903), .B(n902), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(G162), .B(n980), .ZN(n905) );
  XNOR2_X1 U1007 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1008 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1009 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1010 ( .A(n911), .B(n910), .Z(n912) );
  NOR2_X1 U1011 ( .A1(G37), .A2(n912), .ZN(G395) );
  NOR2_X1 U1012 ( .A1(G227), .A2(G229), .ZN(n913) );
  XNOR2_X1 U1013 ( .A(KEYINPUT49), .B(n913), .ZN(n914) );
  NOR2_X1 U1014 ( .A1(G397), .A2(n914), .ZN(n918) );
  NOR2_X1 U1015 ( .A1(G401), .A2(n919), .ZN(n915) );
  XNOR2_X1 U1016 ( .A(KEYINPUT113), .B(n915), .ZN(n916) );
  NOR2_X1 U1017 ( .A1(G395), .A2(n916), .ZN(n917) );
  NAND2_X1 U1018 ( .A1(n918), .A2(n917), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(n919), .ZN(G319) );
  INV_X1 U1021 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1022 ( .A(G16), .B(KEYINPUT56), .ZN(n947) );
  XOR2_X1 U1023 ( .A(G168), .B(G1966), .Z(n920) );
  NOR2_X1 U1024 ( .A1(n921), .A2(n920), .ZN(n922) );
  XOR2_X1 U1025 ( .A(KEYINPUT57), .B(n922), .Z(n945) );
  XNOR2_X1 U1026 ( .A(G1971), .B(G303), .ZN(n923) );
  XNOR2_X1 U1027 ( .A(n923), .B(KEYINPUT123), .ZN(n928) );
  NAND2_X1 U1028 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1029 ( .A(KEYINPUT122), .B(n926), .Z(n927) );
  NAND2_X1 U1030 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1031 ( .A(n929), .B(KEYINPUT124), .ZN(n943) );
  XNOR2_X1 U1032 ( .A(G1348), .B(n930), .ZN(n931) );
  NOR2_X1 U1033 ( .A1(n932), .A2(n931), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(n933), .B(G1956), .ZN(n934) );
  XNOR2_X1 U1035 ( .A(n934), .B(KEYINPUT121), .ZN(n939) );
  XNOR2_X1 U1036 ( .A(G1341), .B(n935), .ZN(n937) );
  XNOR2_X1 U1037 ( .A(G171), .B(G1961), .ZN(n936) );
  NAND2_X1 U1038 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1039 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1040 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1041 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n975) );
  INV_X1 U1044 ( .A(G16), .ZN(n973) );
  XNOR2_X1 U1045 ( .A(KEYINPUT125), .B(G5), .ZN(n949) );
  XNOR2_X1 U1046 ( .A(n949), .B(n948), .ZN(n956) );
  XNOR2_X1 U1047 ( .A(G1971), .B(G22), .ZN(n951) );
  XNOR2_X1 U1048 ( .A(G23), .B(G1976), .ZN(n950) );
  NOR2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n953) );
  XOR2_X1 U1050 ( .A(G1986), .B(G24), .Z(n952) );
  NAND2_X1 U1051 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1052 ( .A(KEYINPUT58), .B(n954), .ZN(n955) );
  NOR2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n968) );
  XOR2_X1 U1054 ( .A(KEYINPUT126), .B(G4), .Z(n958) );
  XNOR2_X1 U1055 ( .A(G1348), .B(KEYINPUT59), .ZN(n957) );
  XNOR2_X1 U1056 ( .A(n958), .B(n957), .ZN(n965) );
  XNOR2_X1 U1057 ( .A(G19), .B(n959), .ZN(n963) );
  XNOR2_X1 U1058 ( .A(G1956), .B(G20), .ZN(n961) );
  XNOR2_X1 U1059 ( .A(G1981), .B(G6), .ZN(n960) );
  NOR2_X1 U1060 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1061 ( .A1(n963), .A2(n962), .ZN(n964) );
  NOR2_X1 U1062 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1063 ( .A(n966), .B(KEYINPUT60), .ZN(n967) );
  NAND2_X1 U1064 ( .A1(n968), .A2(n967), .ZN(n970) );
  XNOR2_X1 U1065 ( .A(G21), .B(G1966), .ZN(n969) );
  NOR2_X1 U1066 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1067 ( .A(KEYINPUT61), .B(n971), .ZN(n972) );
  NAND2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1070 ( .A(n976), .B(KEYINPUT127), .ZN(n1007) );
  XOR2_X1 U1071 ( .A(G160), .B(G2084), .Z(n977) );
  NOR2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n987) );
  XNOR2_X1 U1074 ( .A(KEYINPUT115), .B(KEYINPUT51), .ZN(n985) );
  XOR2_X1 U1075 ( .A(G2090), .B(G162), .Z(n981) );
  XNOR2_X1 U1076 ( .A(KEYINPUT114), .B(n981), .ZN(n983) );
  NOR2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1078 ( .A(n985), .B(n984), .Z(n986) );
  NOR2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1082 ( .A(n992), .B(KEYINPUT116), .ZN(n994) );
  NAND2_X1 U1083 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1084 ( .A(KEYINPUT117), .B(n995), .Z(n1001) );
  XOR2_X1 U1085 ( .A(G2072), .B(n996), .Z(n998) );
  XOR2_X1 U1086 ( .A(G164), .B(G2078), .Z(n997) );
  NOR2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1088 ( .A(KEYINPUT50), .B(n999), .Z(n1000) );
  NOR2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1090 ( .A(KEYINPUT52), .B(n1002), .ZN(n1004) );
  INV_X1 U1091 ( .A(KEYINPUT55), .ZN(n1003) );
  NAND2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1093 ( .A1(n1005), .A2(G29), .ZN(n1006) );
  NAND2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1033) );
  XNOR2_X1 U1095 ( .A(G29), .B(KEYINPUT119), .ZN(n1029) );
  XNOR2_X1 U1096 ( .A(G25), .B(n1008), .ZN(n1009) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(G28), .ZN(n1016) );
  XOR2_X1 U1098 ( .A(n1010), .B(G27), .Z(n1013) );
  XOR2_X1 U1099 ( .A(n1011), .B(G32), .Z(n1012) );
  NOR2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1101 ( .A(KEYINPUT118), .B(n1014), .Z(n1015) );
  NOR2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1020) );
  XNOR2_X1 U1103 ( .A(G2067), .B(G26), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(G33), .B(G2072), .ZN(n1017) );
  NOR2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1107 ( .A(n1021), .B(KEYINPUT53), .ZN(n1024) );
  XOR2_X1 U1108 ( .A(G2084), .B(G34), .Z(n1022) );
  XNOR2_X1 U1109 ( .A(KEYINPUT54), .B(n1022), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1026) );
  XNOR2_X1 U1111 ( .A(G35), .B(G2090), .ZN(n1025) );
  NOR2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1113 ( .A(KEYINPUT55), .B(n1027), .ZN(n1028) );
  NAND2_X1 U1114 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1115 ( .A1(G11), .A2(n1030), .ZN(n1031) );
  XNOR2_X1 U1116 ( .A(KEYINPUT120), .B(n1031), .ZN(n1032) );
  NOR2_X1 U1117 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XNOR2_X1 U1118 ( .A(KEYINPUT62), .B(n1034), .ZN(G311) );
  INV_X1 U1119 ( .A(G311), .ZN(G150) );
endmodule

