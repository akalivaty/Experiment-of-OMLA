

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781;

  INV_X1 U378 ( .A(G953), .ZN(n765) );
  XOR2_X1 U379 ( .A(n503), .B(KEYINPUT104), .Z(n356) );
  AND2_X2 U380 ( .A1(n398), .A2(n369), .ZN(n397) );
  NAND2_X2 U381 ( .A1(n413), .A2(n412), .ZN(n706) );
  AND2_X2 U382 ( .A1(n415), .A2(n414), .ZN(n413) );
  XNOR2_X2 U383 ( .A(n452), .B(G122), .ZN(n527) );
  XNOR2_X2 U384 ( .A(G113), .B(G104), .ZN(n452) );
  NOR2_X2 U385 ( .A1(n541), .A2(n706), .ZN(n504) );
  XNOR2_X1 U386 ( .A(n441), .B(n440), .ZN(n439) );
  BUF_X1 U387 ( .A(G143), .Z(n375) );
  NAND2_X1 U388 ( .A1(n633), .A2(n373), .ZN(n637) );
  NOR2_X1 U389 ( .A1(n635), .A2(n634), .ZN(n733) );
  NOR2_X1 U390 ( .A1(n774), .A2(n422), .ZN(n421) );
  XNOR2_X1 U391 ( .A(n556), .B(n555), .ZN(n775) );
  XNOR2_X1 U392 ( .A(n560), .B(n559), .ZN(n774) );
  AND2_X1 U393 ( .A1(n543), .A2(n716), .ZN(n677) );
  INV_X1 U394 ( .A(n597), .ZN(n688) );
  INV_X1 U395 ( .A(n576), .ZN(n357) );
  NAND2_X1 U396 ( .A1(n396), .A2(n395), .ZN(n394) );
  NAND2_X1 U397 ( .A1(n419), .A2(n418), .ZN(n417) );
  XNOR2_X1 U398 ( .A(n669), .B(n668), .ZN(n670) );
  INV_X1 U399 ( .A(n645), .ZN(n419) );
  OR2_X1 U400 ( .A1(n439), .A2(G902), .ZN(n404) );
  NAND2_X1 U401 ( .A1(n447), .A2(n446), .ZN(n360) );
  AND2_X1 U402 ( .A1(G217), .A2(n501), .ZN(n441) );
  XNOR2_X1 U403 ( .A(n428), .B(G110), .ZN(n488) );
  INV_X1 U404 ( .A(n631), .ZN(n570) );
  XNOR2_X1 U405 ( .A(n762), .B(G146), .ZN(n482) );
  XOR2_X1 U406 ( .A(G137), .B(G140), .Z(n494) );
  XOR2_X1 U407 ( .A(G902), .B(KEYINPUT15), .Z(n631) );
  NAND2_X1 U408 ( .A1(n357), .A2(n358), .ZN(n412) );
  NOR2_X1 U409 ( .A1(n356), .A2(n416), .ZN(n358) );
  BUF_X1 U410 ( .A(n753), .Z(n359) );
  XNOR2_X1 U411 ( .A(n393), .B(n426), .ZN(n753) );
  NAND2_X1 U412 ( .A1(n447), .A2(n446), .ZN(n469) );
  NAND2_X1 U413 ( .A1(n445), .A2(n444), .ZN(n361) );
  XNOR2_X1 U414 ( .A(n507), .B(KEYINPUT4), .ZN(n362) );
  INV_X1 U415 ( .A(n582), .ZN(n363) );
  XNOR2_X1 U416 ( .A(n417), .B(G469), .ZN(n591) );
  XNOR2_X1 U417 ( .A(n360), .B(n752), .ZN(n364) );
  XNOR2_X1 U418 ( .A(n469), .B(n752), .ZN(n486) );
  XNOR2_X1 U419 ( .A(n361), .B(KEYINPUT4), .ZN(n365) );
  BUF_X1 U420 ( .A(n600), .Z(n366) );
  XNOR2_X2 U421 ( .A(n600), .B(n459), .ZN(n613) );
  NOR2_X1 U422 ( .A1(G953), .A2(G237), .ZN(n518) );
  XNOR2_X1 U423 ( .A(G128), .B(KEYINPUT93), .ZN(n487) );
  XOR2_X1 U424 ( .A(KEYINPUT78), .B(KEYINPUT23), .Z(n490) );
  XNOR2_X1 U425 ( .A(n375), .B(G140), .ZN(n516) );
  INV_X1 U426 ( .A(KEYINPUT48), .ZN(n435) );
  XOR2_X1 U427 ( .A(KEYINPUT76), .B(KEYINPUT5), .Z(n484) );
  XNOR2_X1 U428 ( .A(n427), .B(G107), .ZN(n505) );
  INV_X1 U429 ( .A(G116), .ZN(n427) );
  INV_X1 U430 ( .A(G119), .ZN(n428) );
  XOR2_X1 U431 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n522) );
  XNOR2_X1 U432 ( .A(G131), .B(KEYINPUT11), .ZN(n521) );
  XOR2_X1 U433 ( .A(KEYINPUT97), .B(KEYINPUT12), .Z(n520) );
  INV_X1 U434 ( .A(KEYINPUT0), .ZN(n467) );
  NOR2_X1 U435 ( .A1(n710), .A2(n405), .ZN(n395) );
  NOR2_X1 U436 ( .A1(G902), .A2(n653), .ZN(n515) );
  INV_X1 U437 ( .A(KEYINPUT6), .ZN(n411) );
  XNOR2_X1 U438 ( .A(n432), .B(n454), .ZN(n391) );
  INV_X1 U439 ( .A(KEYINPUT66), .ZN(n422) );
  NOR2_X1 U440 ( .A1(n781), .A2(n780), .ZN(n431) );
  XNOR2_X1 U441 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n495) );
  INV_X1 U442 ( .A(KEYINPUT83), .ZN(n571) );
  NOR2_X1 U443 ( .A1(G902), .A2(G237), .ZN(n455) );
  XNOR2_X1 U444 ( .A(KEYINPUT24), .B(KEYINPUT92), .ZN(n489) );
  XNOR2_X1 U445 ( .A(n450), .B(n451), .ZN(n432) );
  XNOR2_X1 U446 ( .A(n493), .B(n449), .ZN(n450) );
  XOR2_X1 U447 ( .A(KEYINPUT17), .B(KEYINPUT88), .Z(n449) );
  AND2_X1 U448 ( .A1(n772), .A2(n434), .ZN(n433) );
  INV_X1 U449 ( .A(n693), .ZN(n434) );
  NAND2_X1 U450 ( .A1(G234), .A2(G237), .ZN(n460) );
  INV_X1 U451 ( .A(KEYINPUT25), .ZN(n440) );
  XNOR2_X1 U452 ( .A(n591), .B(KEYINPUT1), .ZN(n376) );
  XNOR2_X1 U453 ( .A(n485), .B(n367), .ZN(n429) );
  XNOR2_X1 U454 ( .A(n448), .B(KEYINPUT71), .ZN(n752) );
  XNOR2_X1 U455 ( .A(n488), .B(n505), .ZN(n426) );
  XOR2_X1 U456 ( .A(KEYINPUT77), .B(KEYINPUT16), .Z(n453) );
  XNOR2_X1 U457 ( .A(n528), .B(n388), .ZN(n638) );
  NAND2_X1 U458 ( .A1(n688), .A2(n386), .ZN(n599) );
  NOR2_X1 U459 ( .A1(n387), .A2(n596), .ZN(n386) );
  AND2_X1 U460 ( .A1(n581), .A2(n409), .ZN(n609) );
  NOR2_X1 U461 ( .A1(n582), .A2(n410), .ZN(n409) );
  INV_X1 U462 ( .A(n588), .ZN(n410) );
  NOR2_X1 U463 ( .A1(n596), .A2(n716), .ZN(n590) );
  NAND2_X1 U464 ( .A1(n586), .A2(n399), .ZN(n425) );
  OR2_X1 U465 ( .A1(n539), .A2(n540), .ZN(n597) );
  INV_X1 U466 ( .A(n376), .ZN(n622) );
  XNOR2_X1 U467 ( .A(n653), .B(KEYINPUT123), .ZN(n654) );
  XNOR2_X1 U468 ( .A(n638), .B(KEYINPUT59), .ZN(n639) );
  XNOR2_X1 U469 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U470 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U471 ( .A(n593), .B(n381), .ZN(n781) );
  XNOR2_X1 U472 ( .A(n382), .B(KEYINPUT111), .ZN(n381) );
  NOR2_X1 U473 ( .A1(n695), .A2(n614), .ZN(n593) );
  INV_X1 U474 ( .A(KEYINPUT42), .ZN(n382) );
  XNOR2_X1 U475 ( .A(n408), .B(KEYINPUT109), .ZN(n776) );
  NAND2_X1 U476 ( .A1(n608), .A2(n609), .ZN(n408) );
  AND2_X1 U477 ( .A1(n607), .A2(n627), .ZN(n608) );
  XNOR2_X1 U478 ( .A(KEYINPUT21), .B(n502), .ZN(n710) );
  XOR2_X1 U479 ( .A(n484), .B(n483), .Z(n367) );
  OR2_X1 U480 ( .A1(n712), .A2(n383), .ZN(n368) );
  OR2_X1 U481 ( .A1(n399), .A2(KEYINPUT67), .ZN(n369) );
  XOR2_X1 U482 ( .A(n620), .B(KEYINPUT74), .Z(n370) );
  XOR2_X1 U483 ( .A(KEYINPUT41), .B(KEYINPUT110), .Z(n371) );
  XNOR2_X1 U484 ( .A(n438), .B(n371), .ZN(n695) );
  XNOR2_X1 U485 ( .A(KEYINPUT30), .B(KEYINPUT108), .ZN(n372) );
  XOR2_X1 U486 ( .A(n632), .B(KEYINPUT65), .Z(n373) );
  INV_X1 U487 ( .A(n749), .ZN(n374) );
  OR2_X1 U488 ( .A1(n541), .A2(n425), .ZN(n424) );
  XNOR2_X1 U489 ( .A(n424), .B(KEYINPUT22), .ZN(n557) );
  INV_X1 U490 ( .A(n598), .ZN(n387) );
  NOR2_X1 U491 ( .A1(n557), .A2(n598), .ZN(n553) );
  AND2_X2 U492 ( .A1(n637), .A2(n636), .ZN(n377) );
  AND2_X2 U493 ( .A1(n637), .A2(n636), .ZN(n741) );
  XNOR2_X1 U494 ( .A(n761), .B(n497), .ZN(n378) );
  XNOR2_X1 U495 ( .A(n761), .B(n497), .ZN(n498) );
  OR2_X2 U496 ( .A1(n667), .A2(G902), .ZN(n407) );
  XNOR2_X1 U497 ( .A(n364), .B(n429), .ZN(n667) );
  NAND2_X1 U498 ( .A1(n709), .A2(n405), .ZN(n398) );
  BUF_X1 U499 ( .A(n574), .Z(n383) );
  BUF_X1 U500 ( .A(n659), .Z(n379) );
  XNOR2_X1 U501 ( .A(n378), .B(n499), .ZN(n380) );
  XNOR2_X1 U502 ( .A(n498), .B(n499), .ZN(n740) );
  XNOR2_X1 U503 ( .A(n486), .B(n753), .ZN(n392) );
  XNOR2_X1 U504 ( .A(n392), .B(n391), .ZN(n659) );
  NOR2_X1 U505 ( .A1(n540), .A2(n538), .ZN(n586) );
  NOR2_X1 U506 ( .A1(n700), .A2(n437), .ZN(n436) );
  XNOR2_X1 U507 ( .A(n385), .B(n435), .ZN(n384) );
  NAND2_X1 U508 ( .A1(n384), .A2(n433), .ZN(n635) );
  XNOR2_X1 U509 ( .A(n457), .B(n456), .ZN(n606) );
  XNOR2_X2 U510 ( .A(n525), .B(n494), .ZN(n761) );
  XNOR2_X2 U511 ( .A(n635), .B(KEYINPUT84), .ZN(n764) );
  NAND2_X1 U512 ( .A1(n621), .A2(n370), .ZN(n385) );
  NOR2_X1 U513 ( .A1(n638), .A2(G902), .ZN(n530) );
  XNOR2_X1 U514 ( .A(n389), .B(n526), .ZN(n388) );
  XNOR2_X1 U515 ( .A(n390), .B(n529), .ZN(n389) );
  INV_X1 U516 ( .A(n527), .ZN(n390) );
  XNOR2_X1 U517 ( .A(n527), .B(n453), .ZN(n393) );
  INV_X1 U518 ( .A(n710), .ZN(n399) );
  NAND2_X2 U519 ( .A1(n397), .A2(n394), .ZN(n576) );
  INV_X1 U520 ( .A(n709), .ZN(n396) );
  OR2_X2 U521 ( .A1(n403), .A2(n400), .ZN(n709) );
  NAND2_X1 U522 ( .A1(n402), .A2(n401), .ZN(n400) );
  NAND2_X1 U523 ( .A1(n439), .A2(G902), .ZN(n401) );
  NAND2_X1 U524 ( .A1(n740), .A2(n439), .ZN(n402) );
  NOR2_X1 U525 ( .A1(n380), .A2(n404), .ZN(n403) );
  INV_X1 U526 ( .A(KEYINPUT67), .ZN(n405) );
  XNOR2_X1 U527 ( .A(n406), .B(n372), .ZN(n575) );
  NAND2_X1 U528 ( .A1(n574), .A2(n697), .ZN(n406) );
  XNOR2_X2 U529 ( .A(n407), .B(G472), .ZN(n574) );
  INV_X1 U530 ( .A(n383), .ZN(n716) );
  XNOR2_X2 U531 ( .A(n574), .B(n411), .ZN(n598) );
  NAND2_X1 U532 ( .A1(n576), .A2(n356), .ZN(n414) );
  NAND2_X1 U533 ( .A1(n416), .A2(n356), .ZN(n415) );
  NAND2_X1 U534 ( .A1(n376), .A2(n598), .ZN(n416) );
  INV_X1 U535 ( .A(n591), .ZN(n582) );
  INV_X1 U536 ( .A(G902), .ZN(n418) );
  INV_X1 U537 ( .A(n775), .ZN(n420) );
  NOR2_X1 U538 ( .A1(n774), .A2(n775), .ZN(n563) );
  NAND2_X1 U539 ( .A1(n421), .A2(n420), .ZN(n423) );
  NAND2_X1 U540 ( .A1(n423), .A2(KEYINPUT44), .ZN(n566) );
  AND2_X1 U541 ( .A1(n430), .A2(n778), .ZN(n621) );
  XNOR2_X1 U542 ( .A(n431), .B(KEYINPUT46), .ZN(n430) );
  NAND2_X1 U543 ( .A1(n698), .A2(n697), .ZN(n703) );
  NAND2_X1 U544 ( .A1(n698), .A2(n436), .ZN(n438) );
  INV_X1 U545 ( .A(n697), .ZN(n437) );
  XNOR2_X2 U546 ( .A(G131), .B(G134), .ZN(n762) );
  NAND2_X1 U547 ( .A1(n606), .A2(n697), .ZN(n600) );
  XNOR2_X1 U548 ( .A(KEYINPUT77), .B(G110), .ZN(n470) );
  NOR2_X1 U549 ( .A1(n702), .A2(n547), .ZN(n548) );
  XNOR2_X1 U550 ( .A(n488), .B(n487), .ZN(n492) );
  INV_X1 U551 ( .A(KEYINPUT38), .ZN(n573) );
  INV_X1 U552 ( .A(KEYINPUT36), .ZN(n601) );
  XNOR2_X1 U553 ( .A(n601), .B(KEYINPUT87), .ZN(n602) );
  INV_X1 U554 ( .A(KEYINPUT19), .ZN(n459) );
  XNOR2_X1 U555 ( .A(n603), .B(n602), .ZN(n604) );
  XNOR2_X1 U556 ( .A(n554), .B(KEYINPUT64), .ZN(n555) );
  INV_X1 U557 ( .A(KEYINPUT124), .ZN(n657) );
  INV_X1 U558 ( .A(G128), .ZN(n442) );
  NAND2_X1 U559 ( .A1(n442), .A2(G143), .ZN(n445) );
  INV_X1 U560 ( .A(G143), .ZN(n443) );
  NAND2_X1 U561 ( .A1(n443), .A2(G128), .ZN(n444) );
  NAND2_X1 U562 ( .A1(n445), .A2(n444), .ZN(n506) );
  XNOR2_X1 U563 ( .A(n506), .B(KEYINPUT4), .ZN(n760) );
  OR2_X2 U564 ( .A1(n760), .A2(G101), .ZN(n447) );
  NAND2_X1 U565 ( .A1(G101), .A2(n365), .ZN(n446) );
  XOR2_X1 U566 ( .A(KEYINPUT70), .B(KEYINPUT3), .Z(n448) );
  XOR2_X2 U567 ( .A(G146), .B(G125), .Z(n493) );
  INV_X1 U568 ( .A(KEYINPUT18), .ZN(n451) );
  NAND2_X1 U569 ( .A1(G224), .A2(n765), .ZN(n454) );
  NOR2_X1 U570 ( .A1(n659), .A2(n631), .ZN(n457) );
  XNOR2_X1 U571 ( .A(n455), .B(KEYINPUT75), .ZN(n458) );
  NAND2_X1 U572 ( .A1(G210), .A2(n458), .ZN(n456) );
  NAND2_X1 U573 ( .A1(G214), .A2(n458), .ZN(n697) );
  XNOR2_X1 U574 ( .A(n460), .B(KEYINPUT14), .ZN(n462) );
  NAND2_X1 U575 ( .A1(G952), .A2(n462), .ZN(n726) );
  NOR2_X1 U576 ( .A1(G953), .A2(n726), .ZN(n461) );
  XOR2_X1 U577 ( .A(KEYINPUT90), .B(n461), .Z(n580) );
  INV_X1 U578 ( .A(n580), .ZN(n465) );
  NAND2_X1 U579 ( .A1(G902), .A2(n462), .ZN(n577) );
  NOR2_X1 U580 ( .A1(G898), .A2(n765), .ZN(n463) );
  XNOR2_X1 U581 ( .A(KEYINPUT91), .B(n463), .ZN(n757) );
  NOR2_X1 U582 ( .A1(n577), .A2(n757), .ZN(n464) );
  NOR2_X1 U583 ( .A1(n465), .A2(n464), .ZN(n466) );
  NOR2_X2 U584 ( .A1(n613), .A2(n466), .ZN(n468) );
  XNOR2_X2 U585 ( .A(n468), .B(n467), .ZN(n541) );
  XNOR2_X1 U586 ( .A(n360), .B(n482), .ZN(n478) );
  INV_X1 U587 ( .A(n470), .ZN(n472) );
  XNOR2_X1 U588 ( .A(G104), .B(G107), .ZN(n471) );
  XNOR2_X1 U589 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U590 ( .A(n494), .B(n473), .ZN(n474) );
  INV_X1 U591 ( .A(n474), .ZN(n476) );
  NAND2_X1 U592 ( .A1(G227), .A2(n765), .ZN(n475) );
  XNOR2_X1 U593 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U594 ( .A(n478), .B(n477), .ZN(n645) );
  XOR2_X1 U595 ( .A(G119), .B(G116), .Z(n480) );
  XNOR2_X1 U596 ( .A(G137), .B(G113), .ZN(n479) );
  XNOR2_X1 U597 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U598 ( .A(n482), .B(n481), .ZN(n485) );
  NAND2_X1 U599 ( .A1(n518), .A2(G210), .ZN(n483) );
  XNOR2_X1 U600 ( .A(n490), .B(n489), .ZN(n491) );
  XOR2_X1 U601 ( .A(n492), .B(n491), .Z(n499) );
  XNOR2_X2 U602 ( .A(n493), .B(KEYINPUT10), .ZN(n525) );
  NAND2_X1 U603 ( .A1(n765), .A2(G234), .ZN(n496) );
  XNOR2_X1 U604 ( .A(n496), .B(n495), .ZN(n510) );
  NAND2_X1 U605 ( .A1(G221), .A2(n510), .ZN(n497) );
  NAND2_X1 U606 ( .A1(n570), .A2(G234), .ZN(n500) );
  XNOR2_X1 U607 ( .A(n500), .B(KEYINPUT20), .ZN(n501) );
  NAND2_X1 U608 ( .A1(G221), .A2(n501), .ZN(n502) );
  XNOR2_X1 U609 ( .A(KEYINPUT33), .B(KEYINPUT72), .ZN(n503) );
  XNOR2_X1 U610 ( .A(n504), .B(KEYINPUT34), .ZN(n533) );
  XOR2_X1 U611 ( .A(KEYINPUT9), .B(n505), .Z(n509) );
  BUF_X1 U612 ( .A(n361), .Z(n507) );
  XNOR2_X1 U613 ( .A(n507), .B(G134), .ZN(n508) );
  XNOR2_X1 U614 ( .A(n509), .B(n508), .ZN(n514) );
  XOR2_X1 U615 ( .A(G122), .B(KEYINPUT7), .Z(n512) );
  NAND2_X1 U616 ( .A1(G217), .A2(n510), .ZN(n511) );
  XNOR2_X1 U617 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U618 ( .A(n514), .B(n513), .ZN(n653) );
  XOR2_X1 U619 ( .A(G478), .B(n515), .Z(n540) );
  XNOR2_X1 U620 ( .A(KEYINPUT13), .B(G475), .ZN(n531) );
  XOR2_X1 U621 ( .A(KEYINPUT98), .B(KEYINPUT96), .Z(n517) );
  XNOR2_X1 U622 ( .A(n517), .B(n516), .ZN(n529) );
  NAND2_X1 U623 ( .A1(G214), .A2(n518), .ZN(n519) );
  XNOR2_X1 U624 ( .A(n520), .B(n519), .ZN(n524) );
  XNOR2_X1 U625 ( .A(n522), .B(n521), .ZN(n523) );
  XOR2_X1 U626 ( .A(n524), .B(n523), .Z(n528) );
  INV_X1 U627 ( .A(n525), .ZN(n526) );
  XNOR2_X1 U628 ( .A(n531), .B(n530), .ZN(n538) );
  NAND2_X1 U629 ( .A1(n540), .A2(n538), .ZN(n532) );
  XNOR2_X1 U630 ( .A(KEYINPUT105), .B(n532), .ZN(n607) );
  NAND2_X1 U631 ( .A1(n533), .A2(n607), .ZN(n534) );
  XNOR2_X1 U632 ( .A(n534), .B(KEYINPUT35), .ZN(n561) );
  NAND2_X1 U633 ( .A1(n561), .A2(KEYINPUT44), .ZN(n535) );
  XNOR2_X1 U634 ( .A(n535), .B(KEYINPUT86), .ZN(n537) );
  INV_X1 U635 ( .A(n709), .ZN(n587) );
  AND2_X1 U636 ( .A1(n587), .A2(n553), .ZN(n536) );
  NAND2_X1 U637 ( .A1(n622), .A2(n536), .ZN(n674) );
  NAND2_X1 U638 ( .A1(n537), .A2(n674), .ZN(n549) );
  XNOR2_X1 U639 ( .A(n538), .B(KEYINPUT101), .ZN(n539) );
  NAND2_X1 U640 ( .A1(n540), .A2(n539), .ZN(n585) );
  INV_X1 U641 ( .A(n585), .ZN(n690) );
  NOR2_X1 U642 ( .A1(n688), .A2(n690), .ZN(n702) );
  NOR2_X1 U643 ( .A1(n541), .A2(n576), .ZN(n544) );
  AND2_X1 U644 ( .A1(n363), .A2(n544), .ZN(n542) );
  XNOR2_X1 U645 ( .A(n542), .B(KEYINPUT94), .ZN(n543) );
  XOR2_X1 U646 ( .A(KEYINPUT31), .B(KEYINPUT95), .Z(n546) );
  NOR2_X1 U647 ( .A1(n622), .A2(n716), .ZN(n708) );
  NAND2_X1 U648 ( .A1(n544), .A2(n708), .ZN(n545) );
  XNOR2_X1 U649 ( .A(n546), .B(n545), .ZN(n691) );
  NOR2_X1 U650 ( .A1(n677), .A2(n691), .ZN(n547) );
  NOR2_X2 U651 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U652 ( .A(n550), .B(KEYINPUT85), .ZN(n568) );
  NOR2_X1 U653 ( .A1(n622), .A2(n587), .ZN(n551) );
  XNOR2_X1 U654 ( .A(KEYINPUT102), .B(n551), .ZN(n552) );
  NAND2_X1 U655 ( .A1(n553), .A2(n552), .ZN(n556) );
  INV_X1 U656 ( .A(KEYINPUT32), .ZN(n554) );
  INV_X1 U657 ( .A(n622), .ZN(n712) );
  NOR2_X1 U658 ( .A1(n557), .A2(n368), .ZN(n558) );
  AND2_X1 U659 ( .A1(n558), .A2(n709), .ZN(n560) );
  INV_X1 U660 ( .A(KEYINPUT103), .ZN(n559) );
  BUF_X1 U661 ( .A(n561), .Z(n773) );
  XNOR2_X1 U662 ( .A(n773), .B(KEYINPUT66), .ZN(n562) );
  NOR2_X1 U663 ( .A1(KEYINPUT44), .A2(n562), .ZN(n564) );
  NAND2_X1 U664 ( .A1(n564), .A2(n563), .ZN(n565) );
  NAND2_X1 U665 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U666 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U667 ( .A(n569), .B(KEYINPUT45), .ZN(n727) );
  NOR2_X1 U668 ( .A1(n727), .A2(n570), .ZN(n572) );
  XNOR2_X1 U669 ( .A(n572), .B(n571), .ZN(n630) );
  XNOR2_X1 U670 ( .A(KEYINPUT73), .B(KEYINPUT39), .ZN(n584) );
  XNOR2_X1 U671 ( .A(n627), .B(n573), .ZN(n698) );
  NOR2_X1 U672 ( .A1(n576), .A2(n575), .ZN(n581) );
  NOR2_X1 U673 ( .A1(G900), .A2(n577), .ZN(n578) );
  NAND2_X1 U674 ( .A1(G953), .A2(n578), .ZN(n579) );
  NAND2_X1 U675 ( .A1(n580), .A2(n579), .ZN(n588) );
  NAND2_X1 U676 ( .A1(n698), .A2(n609), .ZN(n583) );
  XNOR2_X1 U677 ( .A(n584), .B(n583), .ZN(n594) );
  NOR2_X1 U678 ( .A1(n594), .A2(n585), .ZN(n693) );
  INV_X1 U679 ( .A(n586), .ZN(n700) );
  NOR2_X1 U680 ( .A1(n710), .A2(n587), .ZN(n589) );
  NAND2_X1 U681 ( .A1(n589), .A2(n588), .ZN(n596) );
  XNOR2_X1 U682 ( .A(KEYINPUT28), .B(n590), .ZN(n592) );
  NAND2_X1 U683 ( .A1(n592), .A2(n363), .ZN(n614) );
  NOR2_X1 U684 ( .A1(n597), .A2(n594), .ZN(n595) );
  XNOR2_X1 U685 ( .A(KEYINPUT40), .B(n595), .ZN(n780) );
  XNOR2_X1 U686 ( .A(KEYINPUT106), .B(n599), .ZN(n624) );
  NOR2_X1 U687 ( .A1(n624), .A2(n366), .ZN(n603) );
  NAND2_X1 U688 ( .A1(n604), .A2(n712), .ZN(n605) );
  XNOR2_X1 U689 ( .A(n605), .B(KEYINPUT112), .ZN(n778) );
  BUF_X1 U690 ( .A(n606), .Z(n627) );
  XNOR2_X1 U691 ( .A(n776), .B(KEYINPUT81), .ZN(n611) );
  NAND2_X1 U692 ( .A1(KEYINPUT47), .A2(n702), .ZN(n610) );
  NAND2_X1 U693 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U694 ( .A(KEYINPUT79), .B(n612), .ZN(n619) );
  NOR2_X1 U695 ( .A1(n614), .A2(n613), .ZN(n685) );
  NAND2_X1 U696 ( .A1(KEYINPUT68), .A2(n685), .ZN(n615) );
  XNOR2_X1 U697 ( .A(n615), .B(KEYINPUT47), .ZN(n617) );
  NAND2_X1 U698 ( .A1(n702), .A2(n685), .ZN(n616) );
  NAND2_X1 U699 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U700 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U701 ( .A1(n622), .A2(n697), .ZN(n623) );
  NOR2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U703 ( .A(n625), .B(KEYINPUT43), .ZN(n626) );
  NOR2_X1 U704 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U705 ( .A(KEYINPUT107), .B(n628), .ZN(n772) );
  INV_X1 U706 ( .A(n764), .ZN(n629) );
  NAND2_X1 U707 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U708 ( .A1(n631), .A2(KEYINPUT2), .ZN(n632) );
  INV_X1 U709 ( .A(n727), .ZN(n749) );
  NAND2_X1 U710 ( .A1(n749), .A2(KEYINPUT2), .ZN(n634) );
  INV_X1 U711 ( .A(n733), .ZN(n636) );
  NAND2_X1 U712 ( .A1(n377), .A2(G475), .ZN(n640) );
  XNOR2_X1 U713 ( .A(n640), .B(n639), .ZN(n642) );
  NOR2_X1 U714 ( .A1(G952), .A2(n765), .ZN(n641) );
  XNOR2_X1 U715 ( .A(KEYINPUT89), .B(n641), .ZN(n739) );
  NAND2_X1 U716 ( .A1(n642), .A2(n739), .ZN(n644) );
  INV_X1 U717 ( .A(KEYINPUT60), .ZN(n643) );
  XNOR2_X1 U718 ( .A(n644), .B(n643), .ZN(G60) );
  NAND2_X1 U719 ( .A1(n377), .A2(G469), .ZN(n649) );
  XOR2_X1 U720 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n647) );
  XNOR2_X1 U721 ( .A(n645), .B(KEYINPUT121), .ZN(n646) );
  XNOR2_X1 U722 ( .A(n649), .B(n648), .ZN(n650) );
  NAND2_X1 U723 ( .A1(n650), .A2(n739), .ZN(n652) );
  INV_X1 U724 ( .A(KEYINPUT122), .ZN(n651) );
  XNOR2_X1 U725 ( .A(n652), .B(n651), .ZN(G54) );
  NAND2_X1 U726 ( .A1(n741), .A2(G478), .ZN(n655) );
  XNOR2_X1 U727 ( .A(n655), .B(n654), .ZN(n656) );
  NAND2_X1 U728 ( .A1(n656), .A2(n739), .ZN(n658) );
  XNOR2_X1 U729 ( .A(n658), .B(n657), .ZN(G63) );
  NAND2_X1 U730 ( .A1(n741), .A2(G210), .ZN(n663) );
  XOR2_X1 U731 ( .A(n379), .B(KEYINPUT80), .Z(n661) );
  XOR2_X1 U732 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n660) );
  XNOR2_X1 U733 ( .A(n663), .B(n662), .ZN(n664) );
  NAND2_X1 U734 ( .A1(n664), .A2(n739), .ZN(n666) );
  INV_X1 U735 ( .A(KEYINPUT56), .ZN(n665) );
  XNOR2_X1 U736 ( .A(n666), .B(n665), .ZN(G51) );
  NAND2_X1 U737 ( .A1(n741), .A2(G472), .ZN(n671) );
  INV_X1 U738 ( .A(n667), .ZN(n669) );
  XOR2_X1 U739 ( .A(KEYINPUT62), .B(KEYINPUT113), .Z(n668) );
  XNOR2_X1 U740 ( .A(n671), .B(n670), .ZN(n672) );
  NAND2_X1 U741 ( .A1(n672), .A2(n739), .ZN(n673) );
  XNOR2_X1 U742 ( .A(n673), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U743 ( .A(G101), .B(KEYINPUT114), .ZN(n675) );
  XNOR2_X1 U744 ( .A(n675), .B(n674), .ZN(G3) );
  NAND2_X1 U745 ( .A1(n677), .A2(n688), .ZN(n676) );
  XNOR2_X1 U746 ( .A(n676), .B(G104), .ZN(G6) );
  XOR2_X1 U747 ( .A(KEYINPUT115), .B(KEYINPUT27), .Z(n679) );
  NAND2_X1 U748 ( .A1(n677), .A2(n690), .ZN(n678) );
  XNOR2_X1 U749 ( .A(n679), .B(n678), .ZN(n681) );
  XOR2_X1 U750 ( .A(G107), .B(KEYINPUT26), .Z(n680) );
  XNOR2_X1 U751 ( .A(n681), .B(n680), .ZN(G9) );
  XOR2_X1 U752 ( .A(KEYINPUT29), .B(KEYINPUT116), .Z(n683) );
  NAND2_X1 U753 ( .A1(n685), .A2(n690), .ZN(n682) );
  XNOR2_X1 U754 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U755 ( .A(G128), .B(n684), .ZN(G30) );
  NAND2_X1 U756 ( .A1(n685), .A2(n688), .ZN(n686) );
  XNOR2_X1 U757 ( .A(n686), .B(KEYINPUT118), .ZN(n687) );
  XNOR2_X1 U758 ( .A(G146), .B(n687), .ZN(G48) );
  NAND2_X1 U759 ( .A1(n691), .A2(n688), .ZN(n689) );
  XNOR2_X1 U760 ( .A(n689), .B(G113), .ZN(G15) );
  NAND2_X1 U761 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U762 ( .A(n692), .B(G116), .ZN(G18) );
  XNOR2_X1 U763 ( .A(G134), .B(n693), .ZN(n694) );
  XNOR2_X1 U764 ( .A(n694), .B(KEYINPUT119), .ZN(G36) );
  NOR2_X1 U765 ( .A1(n695), .A2(n706), .ZN(n696) );
  NOR2_X1 U766 ( .A1(G953), .A2(n696), .ZN(n737) );
  NOR2_X1 U767 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U768 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U769 ( .A(n701), .B(KEYINPUT120), .ZN(n705) );
  NOR2_X1 U770 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U771 ( .A1(n705), .A2(n704), .ZN(n707) );
  NOR2_X1 U772 ( .A1(n707), .A2(n706), .ZN(n723) );
  NAND2_X1 U773 ( .A1(n708), .A2(n357), .ZN(n719) );
  NAND2_X1 U774 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U775 ( .A(n711), .B(KEYINPUT49), .ZN(n715) );
  NOR2_X1 U776 ( .A1(n357), .A2(n712), .ZN(n713) );
  XNOR2_X1 U777 ( .A(n713), .B(KEYINPUT50), .ZN(n714) );
  NOR2_X1 U778 ( .A1(n715), .A2(n714), .ZN(n717) );
  NAND2_X1 U779 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U780 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U781 ( .A(KEYINPUT51), .B(n720), .ZN(n721) );
  NOR2_X1 U782 ( .A1(n695), .A2(n721), .ZN(n722) );
  NOR2_X1 U783 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U784 ( .A(n724), .B(KEYINPUT52), .ZN(n725) );
  NOR2_X1 U785 ( .A1(n726), .A2(n725), .ZN(n735) );
  INV_X1 U786 ( .A(KEYINPUT2), .ZN(n729) );
  NAND2_X1 U787 ( .A1(n374), .A2(n729), .ZN(n728) );
  XNOR2_X1 U788 ( .A(n728), .B(KEYINPUT82), .ZN(n731) );
  NAND2_X1 U789 ( .A1(n764), .A2(n729), .ZN(n730) );
  NAND2_X1 U790 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U791 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X1 U792 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U793 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U794 ( .A(KEYINPUT53), .B(n738), .Z(G75) );
  INV_X1 U795 ( .A(n739), .ZN(n745) );
  XNOR2_X1 U796 ( .A(KEYINPUT125), .B(n380), .ZN(n743) );
  NAND2_X1 U797 ( .A1(n377), .A2(G217), .ZN(n742) );
  XOR2_X1 U798 ( .A(n743), .B(n742), .Z(n744) );
  NOR2_X1 U799 ( .A1(n745), .A2(n744), .ZN(G66) );
  NAND2_X1 U800 ( .A1(G224), .A2(G953), .ZN(n746) );
  XNOR2_X1 U801 ( .A(n746), .B(KEYINPUT126), .ZN(n747) );
  XNOR2_X1 U802 ( .A(KEYINPUT61), .B(n747), .ZN(n748) );
  NAND2_X1 U803 ( .A1(G898), .A2(n748), .ZN(n751) );
  NAND2_X1 U804 ( .A1(n749), .A2(n765), .ZN(n750) );
  NAND2_X1 U805 ( .A1(n751), .A2(n750), .ZN(n759) );
  XNOR2_X1 U806 ( .A(KEYINPUT127), .B(n752), .ZN(n754) );
  XNOR2_X1 U807 ( .A(n754), .B(n359), .ZN(n755) );
  XNOR2_X1 U808 ( .A(G101), .B(n755), .ZN(n756) );
  NAND2_X1 U809 ( .A1(n757), .A2(n756), .ZN(n758) );
  XOR2_X1 U810 ( .A(n759), .B(n758), .Z(G69) );
  XNOR2_X1 U811 ( .A(n761), .B(n362), .ZN(n763) );
  XNOR2_X1 U812 ( .A(n763), .B(n762), .ZN(n767) );
  XNOR2_X1 U813 ( .A(n767), .B(n764), .ZN(n766) );
  NAND2_X1 U814 ( .A1(n766), .A2(n765), .ZN(n771) );
  XNOR2_X1 U815 ( .A(G227), .B(n767), .ZN(n768) );
  NAND2_X1 U816 ( .A1(n768), .A2(G900), .ZN(n769) );
  NAND2_X1 U817 ( .A1(n769), .A2(G953), .ZN(n770) );
  NAND2_X1 U818 ( .A1(n771), .A2(n770), .ZN(G72) );
  XNOR2_X1 U819 ( .A(G140), .B(n772), .ZN(G42) );
  XOR2_X1 U820 ( .A(G122), .B(n773), .Z(G24) );
  XOR2_X1 U821 ( .A(n774), .B(G110), .Z(G12) );
  XOR2_X1 U822 ( .A(n775), .B(G119), .Z(G21) );
  XNOR2_X1 U823 ( .A(n776), .B(n375), .ZN(n777) );
  XNOR2_X1 U824 ( .A(n777), .B(KEYINPUT117), .ZN(G45) );
  XOR2_X1 U825 ( .A(G125), .B(n778), .Z(n779) );
  XNOR2_X1 U826 ( .A(KEYINPUT37), .B(n779), .ZN(G27) );
  XOR2_X1 U827 ( .A(G131), .B(n780), .Z(G33) );
  XOR2_X1 U828 ( .A(n781), .B(G137), .Z(G39) );
endmodule

