//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 0 0 0 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 1 0 1 1 1 1 1 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n210, new_n211, new_n212, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1261, new_n1262, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1344, new_n1345, new_n1346;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  INV_X1    g0009(.A(G97), .ZN(new_n210));
  INV_X1    g0010(.A(G107), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G87), .ZN(G355));
  INV_X1    g0013(.A(G1), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT66), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n217), .B1(new_n219), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  INV_X1    g0025(.A(KEYINPUT65), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n226), .B1(new_n217), .B2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(G13), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n216), .A2(KEYINPUT65), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n230), .B(G250), .C1(G257), .C2(G264), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT0), .Z(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n233), .A2(new_n215), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n206), .A2(new_n207), .ZN(new_n235));
  AOI211_X1 g0035(.A(new_n225), .B(new_n232), .C1(new_n234), .C2(new_n235), .ZN(G361));
  XOR2_X1   g0036(.A(G238), .B(G244), .Z(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G226), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  NAND2_X1  g0045(.A1(new_n207), .A2(G68), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n203), .A2(G50), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G87), .B(G97), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(new_n250), .B(new_n253), .Z(G351));
  NAND2_X1  g0054(.A1(G33), .A2(G283), .ZN(new_n255));
  OAI211_X1 g0055(.A(new_n255), .B(new_n215), .C1(G33), .C2(new_n210), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n233), .ZN(new_n258));
  INV_X1    g0058(.A(G116), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G20), .ZN(new_n260));
  AND3_X1   g0060(.A1(new_n258), .A2(KEYINPUT81), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(KEYINPUT81), .B1(new_n258), .B2(new_n260), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n256), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT20), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI211_X1 g0065(.A(KEYINPUT20), .B(new_n256), .C1(new_n261), .C2(new_n262), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n214), .A2(G13), .A3(G20), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(new_n258), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n269), .B1(G1), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G116), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n267), .A2(new_n259), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n265), .A2(new_n266), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G41), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(G1), .A3(G13), .ZN(new_n276));
  NOR2_X1   g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n278), .A2(G303), .A3(new_n279), .ZN(new_n280));
  AND2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  OAI211_X1 g0081(.A(G264), .B(G1698), .C1(new_n281), .C2(new_n277), .ZN(new_n282));
  AND2_X1   g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  AND2_X1   g0083(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n284));
  NOR2_X1   g0084(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT3), .B(G33), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n286), .A2(new_n287), .A3(G257), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n276), .B1(new_n283), .B2(new_n288), .ZN(new_n289));
  AND2_X1   g0089(.A1(new_n276), .A2(G274), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n214), .A2(G45), .ZN(new_n291));
  OR2_X1    g0091(.A1(KEYINPUT5), .A2(G41), .ZN(new_n292));
  NAND2_X1  g0092(.A1(KEYINPUT5), .A2(G41), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n290), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G45), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(G1), .ZN(new_n297));
  AND2_X1   g0097(.A1(KEYINPUT5), .A2(G41), .ZN(new_n298));
  NOR2_X1   g0098(.A1(KEYINPUT5), .A2(G41), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n276), .ZN(new_n301));
  INV_X1    g0101(.A(G270), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n295), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(G169), .B1(new_n289), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT82), .B1(new_n274), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n274), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n233), .B1(G33), .B2(G41), .ZN(new_n307));
  INV_X1    g0107(.A(new_n288), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n280), .A2(new_n282), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n292), .A2(new_n293), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n307), .B1(new_n297), .B2(new_n311), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n312), .A2(G270), .B1(new_n294), .B2(new_n290), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n310), .A2(new_n313), .A3(G179), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n305), .A2(KEYINPUT21), .B1(new_n306), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT21), .ZN(new_n317));
  OAI211_X1 g0117(.A(KEYINPUT82), .B(new_n317), .C1(new_n274), .C2(new_n304), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n289), .A2(new_n303), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G190), .ZN(new_n320));
  INV_X1    g0120(.A(G200), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n320), .B(new_n274), .C1(new_n321), .C2(new_n319), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n316), .A2(new_n318), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n258), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n208), .A2(G20), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT8), .B(G58), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n215), .A2(G33), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  NOR2_X1   g0129(.A1(G20), .A2(G33), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n327), .A2(new_n329), .B1(G150), .B2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n324), .B1(new_n325), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n269), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n214), .A2(G20), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G50), .ZN(new_n335));
  OAI22_X1  g0135(.A1(new_n333), .A2(new_n335), .B1(G50), .B2(new_n267), .ZN(new_n336));
  OR2_X1    g0136(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n214), .B1(G41), .B2(G45), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n339), .A2(new_n276), .A3(G274), .ZN(new_n340));
  INV_X1    g0140(.A(G226), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n276), .A2(new_n338), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n286), .A2(new_n287), .A3(G222), .ZN(new_n344));
  INV_X1    g0144(.A(G77), .ZN(new_n345));
  INV_X1    g0145(.A(G223), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n287), .A2(G1698), .ZN(new_n347));
  OAI221_X1 g0147(.A(new_n344), .B1(new_n345), .B2(new_n287), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n343), .B1(new_n348), .B2(new_n307), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n337), .B1(G169), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(G179), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  OR3_X1    g0153(.A1(new_n349), .A2(KEYINPUT72), .A3(new_n321), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT9), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n337), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(KEYINPUT72), .B1(new_n349), .B2(new_n321), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n349), .A2(G190), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n354), .A2(new_n356), .A3(new_n357), .A4(new_n358), .ZN(new_n359));
  OR3_X1    g0159(.A1(new_n332), .A2(new_n355), .A3(new_n336), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n360), .B(KEYINPUT71), .ZN(new_n361));
  OR3_X1    g0161(.A1(new_n359), .A2(new_n361), .A3(KEYINPUT10), .ZN(new_n362));
  OAI21_X1  g0162(.A(KEYINPUT10), .B1(new_n361), .B2(new_n359), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n353), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(G33), .A2(G97), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT68), .ZN(new_n366));
  INV_X1    g0166(.A(G1698), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n368), .B(new_n369), .C1(new_n281), .C2(new_n277), .ZN(new_n370));
  INV_X1    g0170(.A(G232), .ZN(new_n371));
  OAI221_X1 g0171(.A(new_n365), .B1(new_n370), .B2(new_n341), .C1(new_n371), .C2(new_n347), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n307), .ZN(new_n373));
  INV_X1    g0173(.A(G238), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n340), .B1(new_n374), .B2(new_n342), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT13), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT13), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n373), .A2(new_n379), .A3(new_n376), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n378), .A2(G190), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n379), .B1(new_n373), .B2(new_n376), .ZN(new_n382));
  AOI211_X1 g0182(.A(KEYINPUT13), .B(new_n375), .C1(new_n372), .C2(new_n307), .ZN(new_n383));
  OAI21_X1  g0183(.A(G200), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n268), .A2(new_n203), .ZN(new_n385));
  XNOR2_X1  g0185(.A(new_n385), .B(KEYINPUT12), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n269), .A2(G68), .A3(new_n334), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT11), .ZN(new_n388));
  INV_X1    g0188(.A(new_n330), .ZN(new_n389));
  OAI22_X1  g0189(.A1(new_n389), .A2(new_n207), .B1(new_n215), .B2(G68), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n328), .A2(new_n345), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n258), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n386), .B(new_n387), .C1(new_n388), .C2(new_n392), .ZN(new_n393));
  AND2_X1   g0193(.A1(new_n392), .A2(new_n388), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AND3_X1   g0195(.A1(new_n381), .A2(new_n384), .A3(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(G169), .B1(new_n382), .B2(new_n383), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT14), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n378), .A2(G179), .A3(new_n380), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT14), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n400), .B(G169), .C1(new_n382), .C2(new_n383), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n398), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n395), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n396), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n327), .A2(new_n334), .ZN(new_n405));
  OAI22_X1  g0205(.A1(new_n333), .A2(new_n405), .B1(new_n267), .B2(new_n327), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n204), .B(new_n205), .C1(new_n202), .C2(new_n203), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n407), .A2(G20), .B1(G159), .B2(new_n330), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT7), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n287), .B2(G20), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n281), .A2(new_n277), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n411), .A2(KEYINPUT7), .A3(new_n215), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n408), .B1(new_n413), .B2(new_n203), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT16), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n324), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n412), .A2(KEYINPUT73), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT73), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n411), .A2(new_n418), .A3(KEYINPUT7), .A4(new_n215), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n417), .A2(new_n410), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(G68), .ZN(new_n421));
  AND2_X1   g0221(.A1(new_n408), .A2(KEYINPUT16), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n406), .B1(new_n416), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n340), .B1(new_n371), .B2(new_n342), .ZN(new_n425));
  XNOR2_X1  g0225(.A(new_n425), .B(KEYINPUT74), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n287), .A2(G226), .A3(G1698), .ZN(new_n427));
  NAND2_X1  g0227(.A1(G33), .A2(G87), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n427), .B(new_n428), .C1(new_n346), .C2(new_n370), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n307), .ZN(new_n430));
  INV_X1    g0230(.A(G190), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n425), .B1(new_n429), .B2(new_n307), .ZN(new_n433));
  OAI22_X1  g0233(.A1(new_n426), .A2(new_n432), .B1(G200), .B2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT17), .B1(new_n424), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n430), .A2(new_n351), .ZN(new_n437));
  OAI22_X1  g0237(.A1(new_n426), .A2(new_n437), .B1(G169), .B2(new_n433), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT18), .B1(new_n424), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n408), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n203), .B1(new_n410), .B2(new_n412), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n415), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n423), .A2(new_n258), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n406), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT18), .ZN(new_n446));
  INV_X1    g0246(.A(new_n438), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n424), .A2(KEYINPUT17), .A3(new_n434), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n436), .A2(new_n439), .A3(new_n448), .A4(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT69), .ZN(new_n452));
  XNOR2_X1  g0252(.A(new_n326), .B(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n330), .ZN(new_n454));
  XNOR2_X1  g0254(.A(KEYINPUT15), .B(G87), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n456), .A2(new_n329), .B1(G20), .B2(G77), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n324), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n269), .A2(G77), .A3(new_n334), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n459), .B1(G77), .B2(new_n267), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n411), .A2(G107), .ZN(new_n462));
  OAI221_X1 g0262(.A(new_n462), .B1(new_n370), .B2(new_n371), .C1(new_n374), .C2(new_n347), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n307), .ZN(new_n464));
  INV_X1    g0264(.A(new_n342), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n465), .A2(G244), .B1(new_n290), .B2(new_n339), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n461), .A2(KEYINPUT70), .B1(G200), .B2(new_n467), .ZN(new_n468));
  OAI221_X1 g0268(.A(new_n468), .B1(KEYINPUT70), .B2(new_n461), .C1(new_n431), .C2(new_n467), .ZN(new_n469));
  INV_X1    g0269(.A(G169), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n461), .B1(new_n470), .B2(new_n467), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n464), .A2(new_n351), .A3(new_n466), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  AND4_X1   g0274(.A1(new_n364), .A2(new_n404), .A3(new_n451), .A4(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT77), .ZN(new_n476));
  OAI211_X1 g0276(.A(G250), .B(G1698), .C1(new_n281), .C2(new_n277), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n255), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n286), .A2(new_n287), .A3(G244), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n478), .B1(new_n479), .B2(KEYINPUT4), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT4), .ZN(new_n481));
  INV_X1    g0281(.A(G244), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n481), .B1(new_n370), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT76), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n286), .A2(new_n287), .A3(G244), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT76), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n485), .A2(new_n486), .A3(new_n481), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n480), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n307), .ZN(new_n489));
  INV_X1    g0289(.A(G257), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n295), .B1(new_n301), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n476), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  AOI211_X1 g0293(.A(KEYINPUT77), .B(new_n491), .C1(new_n488), .C2(new_n307), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n470), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n491), .B1(new_n488), .B2(new_n307), .ZN(new_n496));
  INV_X1    g0296(.A(new_n271), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G97), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n268), .A2(new_n210), .ZN(new_n499));
  OR2_X1    g0299(.A1(new_n499), .A2(KEYINPUT75), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(KEYINPUT75), .ZN(new_n501));
  AND2_X1   g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT6), .ZN(new_n504));
  NOR3_X1   g0304(.A1(new_n504), .A2(new_n210), .A3(G107), .ZN(new_n505));
  XNOR2_X1  g0305(.A(G97), .B(G107), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n505), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  OAI22_X1  g0307(.A1(new_n507), .A2(new_n215), .B1(new_n345), .B2(new_n389), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n211), .B1(new_n410), .B2(new_n412), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n258), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n496), .A2(new_n351), .B1(new_n503), .B2(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n286), .A2(new_n287), .A3(KEYINPUT4), .A4(G244), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n512), .A2(new_n255), .A3(new_n477), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n486), .B1(new_n485), .B2(new_n481), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n276), .B1(new_n515), .B2(new_n487), .ZN(new_n516));
  OAI21_X1  g0316(.A(KEYINPUT77), .B1(new_n516), .B2(new_n491), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n489), .A2(new_n476), .A3(new_n492), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n517), .A2(G190), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n510), .A2(new_n498), .A3(new_n502), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n489), .A2(new_n492), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n520), .B1(new_n521), .B2(G200), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n495), .A2(new_n511), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  OAI211_X1 g0323(.A(G257), .B(G1698), .C1(new_n281), .C2(new_n277), .ZN(new_n524));
  INV_X1    g0324(.A(G294), .ZN(new_n525));
  INV_X1    g0325(.A(G250), .ZN(new_n526));
  OAI221_X1 g0326(.A(new_n524), .B1(new_n270), .B2(new_n525), .C1(new_n370), .C2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(G264), .ZN(new_n528));
  OAI21_X1  g0328(.A(KEYINPUT84), .B1(new_n301), .B2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT84), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n300), .A2(new_n530), .A3(G264), .A4(new_n276), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n307), .A2(new_n527), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n532), .A2(new_n351), .A3(new_n295), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n529), .A2(new_n531), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n524), .B1(new_n270), .B2(new_n525), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n370), .A2(new_n526), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n307), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n534), .A2(new_n295), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n470), .ZN(new_n539));
  NAND2_X1  g0339(.A1(G33), .A2(G116), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n540), .A2(G20), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT23), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n542), .B1(new_n215), .B2(G107), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n211), .A2(KEYINPUT23), .A3(G20), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n541), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n215), .B(G87), .C1(new_n281), .C2(new_n277), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n546), .A2(KEYINPUT22), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n546), .A2(KEYINPUT22), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n545), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(KEYINPUT24), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT24), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n551), .B(new_n545), .C1(new_n547), .C2(new_n548), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n324), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT83), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT25), .ZN(new_n555));
  AOI211_X1 g0355(.A(G107), .B(new_n267), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n554), .A2(new_n555), .ZN(new_n557));
  XNOR2_X1  g0357(.A(new_n556), .B(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n211), .B2(new_n271), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n533), .B(new_n539), .C1(new_n553), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n538), .A2(new_n321), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n561), .B1(G190), .B2(new_n538), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n553), .A2(new_n559), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n287), .A2(new_n215), .A3(G68), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT19), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n215), .B1(new_n365), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(G87), .B2(new_n212), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n566), .B1(new_n328), .B2(new_n210), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n565), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  OR2_X1    g0370(.A1(new_n570), .A2(KEYINPUT79), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n324), .B1(new_n570), .B2(KEYINPUT79), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n571), .A2(new_n572), .B1(new_n268), .B2(new_n455), .ZN(new_n573));
  XNOR2_X1  g0373(.A(new_n455), .B(KEYINPUT80), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n497), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n287), .A2(G244), .A3(G1698), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n577), .B(new_n540), .C1(new_n374), .C2(new_n370), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n307), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n526), .B1(new_n214), .B2(G45), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT78), .B1(new_n580), .B2(new_n276), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(new_n276), .A3(KEYINPUT78), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n582), .A2(new_n583), .B1(new_n297), .B2(new_n290), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n470), .ZN(new_n586));
  INV_X1    g0386(.A(new_n583), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n276), .A2(G274), .ZN(new_n588));
  OAI22_X1  g0388(.A1(new_n587), .A2(new_n581), .B1(new_n291), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n589), .B1(new_n307), .B2(new_n578), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n351), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n576), .A2(new_n586), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(G190), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n585), .A2(G200), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n497), .A2(G87), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n593), .A2(new_n573), .A3(new_n594), .A4(new_n595), .ZN(new_n596));
  AND4_X1   g0396(.A1(new_n560), .A2(new_n564), .A3(new_n592), .A4(new_n596), .ZN(new_n597));
  AND4_X1   g0397(.A1(new_n323), .A2(new_n475), .A3(new_n523), .A4(new_n597), .ZN(G372));
  NAND2_X1  g0398(.A1(new_n362), .A2(new_n363), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n436), .A2(new_n449), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n402), .A2(new_n403), .ZN(new_n601));
  INV_X1    g0401(.A(new_n473), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n381), .A2(new_n384), .A3(new_n395), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n600), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n448), .A2(new_n439), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n599), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n353), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(KEYINPUT86), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT86), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n607), .A2(new_n611), .A3(new_n608), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n475), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n316), .A2(new_n318), .A3(new_n560), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n495), .A2(new_n511), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n573), .A2(new_n595), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n593), .A2(new_n594), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n617), .A2(new_n618), .B1(new_n562), .B2(new_n563), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n519), .A2(new_n522), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n615), .A2(new_n616), .A3(new_n619), .A4(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n592), .ZN(new_n622));
  AOI21_X1  g0422(.A(G169), .B1(new_n517), .B2(new_n518), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n520), .B1(new_n521), .B2(G179), .ZN(new_n624));
  OAI21_X1  g0424(.A(KEYINPUT85), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT85), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n495), .A2(new_n626), .A3(new_n511), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n592), .A2(new_n596), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n625), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT26), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n517), .A2(new_n518), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n624), .B1(new_n632), .B2(new_n470), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n633), .A2(new_n628), .A3(KEYINPUT26), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n622), .B1(new_n631), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n613), .B1(new_n614), .B2(new_n636), .ZN(G369));
  NAND2_X1  g0437(.A1(new_n305), .A2(KEYINPUT21), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n306), .A2(new_n315), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n638), .A2(new_n318), .A3(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n214), .A2(new_n215), .A3(G13), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n641), .A2(KEYINPUT27), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(KEYINPUT27), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(new_n643), .A3(G213), .ZN(new_n644));
  INV_X1    g0444(.A(G343), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n274), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n640), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n648), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n316), .A2(new_n318), .A3(new_n322), .A4(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT87), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n649), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n652), .B1(new_n649), .B2(new_n651), .ZN(new_n654));
  OAI21_X1  g0454(.A(G330), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n564), .B(new_n560), .C1(new_n563), .C2(new_n647), .ZN(new_n657));
  INV_X1    g0457(.A(new_n560), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n646), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n640), .A2(new_n560), .A3(new_n564), .A4(new_n647), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n658), .A2(new_n647), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n661), .A2(new_n665), .ZN(G399));
  INV_X1    g0466(.A(new_n230), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(G41), .ZN(new_n668));
  NOR3_X1   g0468(.A1(new_n212), .A2(G87), .A3(G116), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NOR3_X1   g0470(.A1(new_n668), .A2(new_n214), .A3(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n671), .B1(new_n235), .B2(new_n668), .ZN(new_n672));
  XOR2_X1   g0472(.A(new_n672), .B(KEYINPUT28), .Z(new_n673));
  INV_X1    g0473(.A(G330), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n351), .B1(new_n289), .B2(new_n303), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(new_n590), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT88), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n521), .A2(new_n676), .A3(new_n677), .A4(new_n538), .ZN(new_n678));
  AOI21_X1  g0478(.A(G179), .B1(new_n310), .B2(new_n313), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n538), .A2(new_n679), .A3(new_n585), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT88), .B1(new_n680), .B2(new_n496), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n534), .A2(new_n579), .A3(new_n537), .A4(new_n584), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT30), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n683), .A2(new_n684), .A3(new_n314), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n517), .A2(new_n685), .A3(new_n518), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n493), .A2(new_n494), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n315), .A2(new_n532), .A3(new_n590), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(KEYINPUT30), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n646), .B1(new_n687), .B2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT31), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n684), .B1(new_n632), .B2(new_n689), .ZN(new_n694));
  OAI211_X1 g0494(.A(new_n694), .B(new_n686), .C1(new_n496), .C2(new_n680), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n647), .A2(new_n693), .ZN(new_n696));
  AOI22_X1  g0496(.A1(new_n692), .A2(new_n693), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n597), .A2(new_n523), .A3(new_n323), .A4(new_n647), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n674), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT29), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n636), .B2(new_n646), .ZN(new_n701));
  INV_X1    g0501(.A(new_n622), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n633), .A2(new_n628), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n630), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n625), .A2(new_n627), .A3(KEYINPUT26), .A4(new_n628), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n646), .B1(new_n702), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(KEYINPUT29), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n699), .B1(new_n701), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n673), .B1(new_n709), .B2(G1), .ZN(G364));
  NOR2_X1   g0510(.A1(new_n228), .A2(G20), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n214), .B1(new_n711), .B2(G45), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n668), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n233), .B1(G20), .B2(new_n470), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(G20), .A2(G179), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT92), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n719), .A2(G190), .A3(G200), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(G190), .A2(G200), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  AOI22_X1  g0523(.A1(new_n721), .A2(G50), .B1(new_n723), .B2(G77), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n719), .A2(G190), .A3(new_n321), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n724), .B1(new_n202), .B2(new_n725), .ZN(new_n726));
  XOR2_X1   g0526(.A(new_n726), .B(KEYINPUT93), .Z(new_n727));
  NOR2_X1   g0527(.A1(new_n215), .A2(G179), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(new_n722), .ZN(new_n729));
  INV_X1    g0529(.A(G159), .ZN(new_n730));
  OR3_X1    g0530(.A1(new_n729), .A2(KEYINPUT32), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(KEYINPUT32), .B1(new_n729), .B2(new_n730), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n728), .A2(G190), .A3(G200), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G87), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n321), .A2(G190), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n728), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n736), .B(new_n287), .C1(new_n211), .C2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(G179), .A2(G200), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n215), .B1(new_n740), .B2(G190), .ZN(new_n741));
  OR2_X1    g0541(.A1(new_n741), .A2(KEYINPUT95), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(KEYINPUT95), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI211_X1 g0544(.A(new_n733), .B(new_n739), .C1(G97), .C2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT94), .ZN(new_n746));
  AND3_X1   g0546(.A1(new_n719), .A2(new_n746), .A3(new_n737), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n746), .B1(new_n719), .B2(new_n737), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n727), .B(new_n745), .C1(new_n203), .C2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n738), .ZN(new_n751));
  INV_X1    g0551(.A(new_n729), .ZN(new_n752));
  AOI22_X1  g0552(.A1(G283), .A2(new_n751), .B1(new_n752), .B2(G329), .ZN(new_n753));
  INV_X1    g0553(.A(G303), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n753), .B(new_n411), .C1(new_n754), .C2(new_n734), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n755), .B1(G311), .B2(new_n723), .ZN(new_n756));
  INV_X1    g0556(.A(new_n749), .ZN(new_n757));
  XNOR2_X1  g0557(.A(KEYINPUT33), .B(G317), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n725), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G322), .ZN(new_n761));
  XOR2_X1   g0561(.A(KEYINPUT96), .B(G326), .Z(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI22_X1  g0563(.A1(new_n744), .A2(G294), .B1(new_n721), .B2(new_n763), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n756), .A2(new_n759), .A3(new_n761), .A4(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n717), .B1(new_n750), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G13), .A2(G33), .ZN(new_n767));
  XOR2_X1   g0567(.A(new_n767), .B(KEYINPUT90), .Z(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(new_n215), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT91), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n716), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n667), .A2(new_n411), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n773), .A2(G355), .B1(new_n259), .B2(new_n667), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n667), .A2(new_n287), .ZN(new_n775));
  INV_X1    g0575(.A(new_n235), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n775), .B1(G45), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n250), .A2(new_n296), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n774), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  AOI211_X1 g0579(.A(new_n715), .B(new_n766), .C1(new_n772), .C2(new_n779), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n780), .B(KEYINPUT97), .Z(new_n781));
  OR2_X1    g0581(.A1(new_n653), .A2(new_n654), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n781), .B1(new_n783), .B2(new_n771), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n674), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT89), .ZN(new_n786));
  AND3_X1   g0586(.A1(new_n786), .A2(new_n655), .A3(new_n715), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(G396));
  NAND2_X1  g0589(.A1(new_n602), .A2(new_n647), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n469), .B1(new_n461), .B2(new_n647), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n791), .B1(new_n473), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(new_n636), .B2(new_n646), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n474), .A2(new_n647), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n634), .B1(new_n630), .B2(new_n629), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n796), .B1(new_n797), .B2(new_n622), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n699), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n714), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n801), .B1(new_n800), .B2(new_n799), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n716), .A2(new_n767), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n715), .B1(new_n345), .B2(new_n803), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n525), .A2(new_n725), .B1(new_n720), .B2(new_n754), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n751), .A2(G87), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(G311), .B2(new_n752), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n287), .B1(new_n735), .B2(G107), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n723), .ZN(new_n810));
  INV_X1    g0610(.A(new_n744), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n809), .B1(new_n259), .B2(new_n810), .C1(new_n210), .C2(new_n811), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n805), .B(new_n812), .C1(G283), .C2(new_n757), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n721), .A2(G137), .B1(new_n723), .B2(G159), .ZN(new_n814));
  INV_X1    g0614(.A(G143), .ZN(new_n815));
  INV_X1    g0615(.A(G150), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n814), .B1(new_n815), .B2(new_n725), .C1(new_n816), .C2(new_n749), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT34), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n411), .B1(new_n735), .B2(G50), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n751), .A2(G68), .ZN(new_n820));
  INV_X1    g0620(.A(G132), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n819), .B(new_n820), .C1(new_n821), .C2(new_n729), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(G58), .B2(new_n744), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n813), .B1(new_n818), .B2(new_n823), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n804), .B1(new_n824), .B2(new_n717), .C1(new_n793), .C2(new_n768), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n802), .A2(new_n825), .ZN(G384));
  NOR2_X1   g0626(.A1(new_n711), .A2(new_n214), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT40), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n395), .A2(new_n647), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n402), .B2(new_n396), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(KEYINPUT99), .ZN(new_n831));
  INV_X1    g0631(.A(new_n829), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n601), .A2(new_n603), .A3(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT99), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n834), .B(new_n829), .C1(new_n402), .C2(new_n396), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n831), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n793), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n688), .A2(new_n685), .B1(new_n678), .B2(new_n681), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n693), .B(new_n647), .C1(new_n839), .C2(new_n694), .ZN(new_n840));
  NOR3_X1   g0640(.A1(new_n493), .A2(new_n494), .A3(new_n689), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n682), .B(new_n686), .C1(new_n841), .C2(KEYINPUT30), .ZN(new_n842));
  AOI21_X1  g0642(.A(KEYINPUT31), .B1(new_n842), .B2(new_n646), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(KEYINPUT103), .B1(new_n844), .B2(new_n698), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n692), .A2(new_n693), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n842), .A2(KEYINPUT31), .A3(new_n646), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n846), .A2(new_n698), .A3(KEYINPUT103), .A4(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n838), .B1(new_n845), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT38), .ZN(new_n851));
  INV_X1    g0651(.A(new_n644), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n423), .A2(new_n258), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n440), .B1(new_n420), .B2(G68), .ZN(new_n854));
  AOI21_X1  g0654(.A(KEYINPUT16), .B1(new_n854), .B2(KEYINPUT100), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n421), .A2(new_n408), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT100), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n853), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n852), .B1(new_n859), .B2(new_n406), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n851), .B1(new_n450), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n447), .B1(new_n859), .B2(new_n406), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n424), .A2(new_n434), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n863), .A2(new_n860), .A3(new_n864), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n865), .A2(KEYINPUT37), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n445), .A2(new_n447), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n445), .A2(new_n852), .ZN(new_n868));
  XNOR2_X1  g0668(.A(KEYINPUT101), .B(KEYINPUT37), .ZN(new_n869));
  AND4_X1   g0669(.A1(new_n867), .A2(new_n868), .A3(new_n864), .A4(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n862), .B1(new_n866), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n870), .B1(new_n865), .B2(KEYINPUT37), .ZN(new_n872));
  INV_X1    g0672(.A(new_n606), .ZN(new_n873));
  AND4_X1   g0673(.A1(KEYINPUT17), .A2(new_n434), .A3(new_n443), .A4(new_n444), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n874), .A2(new_n435), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n860), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n851), .B1(new_n872), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n871), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n828), .B1(new_n850), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT102), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n436), .A2(new_n881), .A3(new_n449), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT102), .B1(new_n874), .B2(new_n435), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n882), .A2(new_n873), .A3(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n868), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n867), .A2(new_n868), .A3(new_n864), .ZN(new_n887));
  INV_X1    g0687(.A(new_n869), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n887), .B(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT38), .B1(new_n886), .B2(new_n889), .ZN(new_n890));
  NOR3_X1   g0690(.A1(new_n872), .A2(new_n876), .A3(new_n851), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT40), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n880), .B1(new_n850), .B2(new_n892), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n893), .B(KEYINPUT104), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n846), .A2(new_n698), .A3(new_n847), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT103), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n614), .B1(new_n897), .B2(new_n848), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n674), .B1(new_n894), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n894), .B2(new_n898), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT39), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n890), .B2(new_n891), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n402), .A2(new_n403), .A3(new_n647), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n871), .A2(new_n877), .A3(KEYINPUT39), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n902), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n831), .A2(new_n833), .A3(new_n835), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n798), .B2(new_n790), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n878), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n606), .A2(new_n644), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n906), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n701), .A2(new_n708), .A3(new_n475), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n613), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n911), .B(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n827), .B1(new_n900), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n914), .B2(new_n900), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT35), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n507), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n918), .A2(G116), .A3(new_n234), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT98), .ZN(new_n920));
  OAI22_X1  g0720(.A1(new_n919), .A2(new_n920), .B1(new_n917), .B2(new_n507), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(new_n920), .B2(new_n919), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n922), .B(KEYINPUT36), .Z(new_n923));
  OAI21_X1  g0723(.A(G77), .B1(new_n202), .B2(new_n203), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n246), .B1(new_n776), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n925), .A2(G1), .A3(new_n228), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n916), .A2(new_n923), .A3(new_n926), .ZN(G367));
  AOI22_X1  g0727(.A1(new_n775), .A2(new_n244), .B1(new_n667), .B2(new_n456), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n715), .B1(new_n772), .B2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n771), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n617), .A2(new_n647), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n931), .A2(new_n592), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n628), .A2(new_n931), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(G317), .ZN(new_n935));
  OAI221_X1 g0735(.A(new_n411), .B1(new_n729), .B2(new_n935), .C1(new_n210), .C2(new_n738), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n734), .A2(new_n259), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT46), .ZN(new_n938));
  AOI211_X1 g0738(.A(new_n936), .B(new_n938), .C1(G283), .C2(new_n723), .ZN(new_n939));
  INV_X1    g0739(.A(G311), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n754), .A2(new_n725), .B1(new_n720), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n744), .B2(G107), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n939), .B(new_n942), .C1(new_n525), .C2(new_n749), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n811), .A2(new_n203), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  OAI221_X1 g0745(.A(new_n945), .B1(new_n815), .B2(new_n720), .C1(new_n816), .C2(new_n725), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n287), .B1(new_n345), .B2(new_n738), .C1(new_n810), .C2(new_n207), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n749), .A2(new_n730), .ZN(new_n948));
  INV_X1    g0748(.A(G137), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n734), .A2(new_n202), .B1(new_n729), .B2(new_n949), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT109), .ZN(new_n951));
  OR3_X1    g0751(.A1(new_n947), .A2(new_n948), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n943), .B1(new_n946), .B2(new_n952), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n953), .B(KEYINPUT47), .Z(new_n954));
  OAI221_X1 g0754(.A(new_n929), .B1(new_n930), .B2(new_n934), .C1(new_n954), .C2(new_n717), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT44), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT108), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n495), .A2(new_n511), .A3(new_n646), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT105), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n495), .A2(KEYINPUT105), .A3(new_n511), .A4(new_n646), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n520), .A2(new_n646), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n523), .A2(new_n963), .ZN(new_n964));
  AND4_X1   g0764(.A1(new_n957), .A2(new_n962), .A3(new_n664), .A4(new_n964), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n960), .A2(new_n961), .B1(new_n523), .B2(new_n963), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n957), .B1(new_n966), .B2(new_n664), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n956), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(KEYINPUT105), .B1(new_n633), .B2(new_n646), .ZN(new_n969));
  INV_X1    g0769(.A(new_n961), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n964), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n971), .A2(new_n665), .A3(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n972), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n966), .B2(new_n664), .ZN(new_n975));
  AND2_X1   g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(KEYINPUT108), .B1(new_n971), .B2(new_n665), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n966), .A2(new_n957), .A3(new_n664), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n977), .A2(KEYINPUT44), .A3(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n968), .A2(new_n976), .A3(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n661), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n646), .B1(new_n316), .B2(new_n318), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n662), .B1(new_n660), .B2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(new_n655), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n968), .A2(new_n976), .A3(new_n979), .A4(new_n661), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n982), .A2(new_n709), .A3(new_n986), .A4(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n709), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n668), .B(KEYINPUT41), .Z(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n713), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n966), .A2(new_n662), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT42), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n616), .B1(new_n966), .B2(new_n560), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT106), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI211_X1 g0797(.A(KEYINPUT106), .B(new_n616), .C1(new_n966), .C2(new_n560), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n997), .A2(new_n647), .A3(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT43), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n934), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n994), .A2(new_n999), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n934), .A2(KEYINPUT43), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1001), .A2(new_n1000), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n1004), .B(new_n1005), .C1(new_n994), .C2(new_n999), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n1003), .A2(new_n1006), .B1(new_n661), .B2(new_n966), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1005), .B1(new_n994), .B2(new_n999), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1004), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n661), .A2(new_n966), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1010), .A2(new_n1011), .A3(new_n1002), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1007), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n955), .B1(new_n992), .B2(new_n1013), .ZN(G387));
  NAND2_X1  g0814(.A1(new_n986), .A2(new_n713), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT110), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n660), .A2(new_n930), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n773), .A2(new_n670), .B1(new_n211), .B2(new_n667), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n241), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n775), .B1(new_n1019), .B2(new_n296), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n453), .A2(new_n207), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT50), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n296), .B1(new_n203), .B2(new_n345), .ZN(new_n1023));
  NOR3_X1   g0823(.A1(new_n1022), .A2(new_n670), .A3(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1018), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n772), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n714), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n757), .A2(new_n327), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n760), .A2(G50), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n287), .B1(new_n738), .B2(new_n210), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n734), .A2(new_n345), .B1(new_n729), .B2(new_n816), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n1030), .B(new_n1031), .C1(new_n723), .C2(G68), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n744), .A2(new_n574), .B1(new_n721), .B2(G159), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1028), .A2(new_n1029), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n287), .B1(new_n751), .B2(G116), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n744), .A2(G283), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n525), .B2(new_n734), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n810), .A2(new_n754), .B1(new_n935), .B2(new_n725), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(G322), .B2(new_n721), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n940), .B2(new_n749), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT48), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1037), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n1041), .B2(new_n1040), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT49), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1035), .B1(new_n729), .B2(new_n762), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1034), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n1017), .B(new_n1027), .C1(new_n1047), .C2(new_n716), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1016), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n668), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n709), .B2(new_n986), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n709), .B2(new_n986), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1049), .A2(new_n1052), .ZN(G393));
  AOI22_X1  g0853(.A1(new_n775), .A2(new_n253), .B1(G97), .B2(new_n667), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n772), .A2(new_n1054), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT113), .Z(new_n1056));
  AOI22_X1  g0856(.A1(new_n735), .A2(G283), .B1(new_n752), .B2(G322), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1057), .B(new_n411), .C1(new_n211), .C2(new_n738), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G294), .B2(new_n723), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1059), .B1(new_n259), .B2(new_n811), .C1(new_n754), .C2(new_n749), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n940), .A2(new_n725), .B1(new_n720), .B2(new_n935), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT52), .Z(new_n1062));
  NOR2_X1   g0862(.A1(new_n811), .A2(new_n345), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n735), .A2(G68), .B1(new_n752), .B2(G143), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1065), .A2(KEYINPUT114), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n453), .B2(new_n723), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n757), .A2(G50), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n411), .B(new_n806), .C1(new_n1065), .C2(KEYINPUT114), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1064), .A2(new_n1067), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n816), .A2(new_n720), .B1(new_n725), .B2(new_n730), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1071), .B(KEYINPUT51), .Z(new_n1072));
  OAI22_X1  g0872(.A1(new_n1060), .A2(new_n1062), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n715), .B(new_n1056), .C1(new_n716), .C2(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT115), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT112), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n971), .B2(new_n930), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n966), .A2(KEYINPUT112), .A3(new_n771), .ZN(new_n1078));
  AND3_X1   g0878(.A1(new_n1075), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n973), .A2(new_n975), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n965), .A2(new_n967), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1081), .B1(new_n1082), .B2(KEYINPUT44), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n661), .B1(new_n1083), .B2(new_n968), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n987), .ZN(new_n1085));
  OAI21_X1  g0885(.A(KEYINPUT111), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT111), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n987), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1080), .B1(new_n1089), .B2(new_n712), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n709), .A2(new_n986), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1087), .B1(new_n982), .B2(new_n987), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1088), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1091), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(KEYINPUT116), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT116), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1096), .B(new_n1091), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n988), .A2(new_n668), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1090), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(G390));
  AOI21_X1  g0902(.A(new_n606), .B1(new_n875), .B2(new_n881), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n868), .B1(new_n1103), .B2(new_n883), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n887), .B(new_n869), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n851), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(KEYINPUT39), .B1(new_n1106), .B2(new_n871), .ZN(new_n1107));
  AND3_X1   g0907(.A1(new_n871), .A2(new_n877), .A3(KEYINPUT39), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n904), .A2(new_n908), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n904), .B1(new_n1106), .B2(new_n871), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n792), .A2(new_n473), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n791), .B1(new_n707), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1110), .B1(new_n1112), .B2(new_n907), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n695), .A2(new_n696), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n846), .A2(new_n1114), .A3(new_n698), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1115), .A2(new_n836), .A3(G330), .A4(new_n793), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1109), .A2(new_n1113), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n798), .A2(new_n790), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n836), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n903), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n902), .A2(new_n905), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n702), .A2(new_n706), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1122), .A2(new_n647), .A3(new_n1111), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n790), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n836), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n1120), .A2(new_n1121), .B1(new_n1125), .B2(new_n1110), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n838), .B(G330), .C1(new_n845), .C2(new_n849), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1117), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  OAI211_X1 g0928(.A(G330), .B(new_n475), .C1(new_n845), .C2(new_n849), .ZN(new_n1129));
  AND3_X1   g0929(.A1(new_n912), .A2(new_n1129), .A3(new_n613), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n836), .B1(new_n699), .B2(new_n793), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n1132), .A2(new_n1127), .B1(new_n798), .B2(new_n790), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1123), .A2(new_n1116), .A3(new_n790), .ZN(new_n1134));
  OAI211_X1 g0934(.A(G330), .B(new_n793), .C1(new_n845), .C2(new_n849), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1134), .B1(new_n1135), .B2(new_n907), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1130), .B1(new_n1133), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1128), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1109), .A2(new_n1113), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n674), .B(new_n837), .C1(new_n897), .C2(new_n848), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1118), .B1(new_n1140), .B2(new_n1131), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n674), .B(new_n794), .C1(new_n897), .C2(new_n848), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1112), .B(new_n1116), .C1(new_n1143), .C2(new_n836), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1141), .A2(new_n1145), .A3(new_n1117), .A4(new_n1130), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1138), .A2(new_n668), .A3(new_n1146), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1109), .A2(new_n1113), .A3(new_n1116), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1127), .B1(new_n1109), .B2(new_n1113), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n713), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1121), .A2(new_n769), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n803), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n714), .B1(new_n327), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n752), .A2(G294), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n736), .A2(new_n820), .A3(new_n1155), .A4(new_n411), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n1156), .B(new_n1063), .C1(G97), .C2(new_n723), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(G116), .A2(new_n760), .B1(new_n721), .B2(G283), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1157), .B(new_n1158), .C1(new_n211), .C2(new_n749), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1159), .B(KEYINPUT119), .ZN(new_n1160));
  XOR2_X1   g0960(.A(KEYINPUT54), .B(G143), .Z(new_n1161));
  AOI22_X1  g0961(.A1(new_n744), .A2(G159), .B1(new_n723), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n949), .B2(new_n749), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT117), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(G128), .A2(new_n721), .B1(new_n760), .B2(G132), .ZN(new_n1165));
  XOR2_X1   g0965(.A(new_n1165), .B(KEYINPUT118), .Z(new_n1166));
  NOR2_X1   g0966(.A1(new_n734), .A2(new_n816), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT53), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n752), .A2(G125), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n411), .B1(new_n751), .B2(G50), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  OR2_X1    g0971(.A1(new_n1166), .A2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1160), .B1(new_n1164), .B2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1154), .B1(new_n1173), .B2(new_n716), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1152), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1147), .A2(new_n1151), .A3(new_n1175), .ZN(G378));
  NAND2_X1  g0976(.A1(new_n337), .A2(new_n852), .ZN(new_n1177));
  AND2_X1   g0977(.A1(new_n364), .A2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n364), .A2(new_n1177), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  OR3_X1    g0981(.A1(new_n1178), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1181), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(G330), .B1(new_n850), .B2(new_n892), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n837), .B1(new_n897), .B2(new_n848), .ZN(new_n1187));
  AOI21_X1  g0987(.A(KEYINPUT40), .B1(new_n1187), .B2(new_n878), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1185), .B1(new_n1186), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n911), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n828), .B1(new_n1106), .B2(new_n871), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n674), .B1(new_n1187), .B2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n880), .A2(new_n1192), .A3(new_n1184), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n1189), .A2(new_n1190), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1190), .B1(new_n1189), .B2(new_n1193), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n713), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n714), .B1(G50), .B2(new_n1153), .ZN(new_n1197));
  OR2_X1    g0997(.A1(new_n287), .A2(G41), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(G283), .B2(new_n752), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n735), .A2(G77), .B1(new_n751), .B2(G58), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1201), .B(new_n944), .C1(new_n574), .C2(new_n723), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(G107), .A2(new_n760), .B1(new_n721), .B2(G116), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1202), .B(new_n1203), .C1(new_n210), .C2(new_n749), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n1205));
  INV_X1    g1005(.A(G41), .ZN(new_n1206));
  AOI21_X1  g1006(.A(G50), .B1(new_n270), .B2(new_n1206), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n1204), .A2(new_n1205), .B1(new_n1198), .B2(new_n1207), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n744), .A2(G150), .B1(new_n760), .B2(G128), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n721), .A2(G125), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n723), .A2(G137), .B1(new_n735), .B2(new_n1161), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(G132), .B2(new_n757), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1214), .A2(KEYINPUT59), .ZN(new_n1215));
  AOI211_X1 g1015(.A(G33), .B(G41), .C1(new_n751), .C2(G159), .ZN(new_n1216));
  INV_X1    g1016(.A(G124), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1216), .B1(new_n1217), .B2(new_n729), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT121), .Z(new_n1219));
  INV_X1    g1019(.A(KEYINPUT59), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1219), .B1(new_n1213), .B2(new_n1220), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n1208), .B1(new_n1215), .B2(new_n1221), .C1(new_n1205), .C2(new_n1204), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1197), .B1(new_n1222), .B2(new_n716), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n1184), .B2(new_n768), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n1196), .A2(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(KEYINPUT57), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n912), .A2(new_n1129), .A3(new_n613), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n1150), .B2(new_n1145), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n668), .B1(new_n1226), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1189), .A2(new_n1193), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(new_n911), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1189), .A2(new_n1190), .A3(new_n1193), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1130), .B1(new_n1128), .B2(new_n1137), .ZN(new_n1234));
  AOI21_X1  g1034(.A(KEYINPUT57), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1225), .B1(new_n1229), .B2(new_n1235), .ZN(G375));
  NOR2_X1   g1036(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n1227), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1238), .A2(new_n1137), .A3(new_n991), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n907), .A2(new_n767), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT122), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n744), .A2(new_n574), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n287), .B1(new_n751), .B2(G77), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n735), .A2(G97), .B1(new_n752), .B2(G303), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n721), .A2(G294), .B1(new_n723), .B2(G107), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n259), .B2(new_n749), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(KEYINPUT123), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1245), .B(new_n1248), .C1(G283), .C2(new_n760), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n811), .A2(new_n207), .B1(new_n821), .B2(new_n720), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n734), .A2(new_n730), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n287), .B1(new_n738), .B2(new_n202), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n1251), .B(new_n1252), .C1(G128), .C2(new_n752), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n1253), .B1(new_n949), .B2(new_n725), .C1(new_n816), .C2(new_n810), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n1250), .B(new_n1254), .C1(new_n757), .C2(new_n1161), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n716), .B1(new_n1249), .B2(new_n1255), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1256), .B(new_n714), .C1(G68), .C2(new_n1153), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1241), .A2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(new_n1145), .B2(new_n713), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1239), .A2(new_n1259), .ZN(G381));
  OR4_X1    g1060(.A1(G396), .A2(G381), .A3(G384), .A4(G393), .ZN(new_n1261));
  NOR4_X1   g1061(.A1(new_n1261), .A2(G387), .A3(G390), .A4(G378), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1262), .B(new_n1225), .C1(new_n1235), .C2(new_n1229), .ZN(G407));
  OAI21_X1  g1063(.A(new_n1175), .B1(new_n1128), .B2(new_n712), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1050), .B1(new_n1128), .B2(new_n1137), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1264), .B1(new_n1146), .B2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n645), .A2(G213), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1269));
  OAI211_X1 g1069(.A(G407), .B(G213), .C1(G375), .C2(new_n1269), .ZN(G409));
  INV_X1    g1070(.A(KEYINPUT126), .ZN(new_n1271));
  OAI21_X1  g1071(.A(KEYINPUT125), .B1(new_n1101), .B2(G387), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(G393), .B(new_n788), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n990), .B1(new_n988), .B2(new_n709), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1012), .B(new_n1007), .C1(new_n1274), .C2(new_n713), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1099), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1275), .B(new_n955), .C1(new_n1276), .C2(new_n1090), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1096), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1097), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1100), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1090), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1280), .A2(G387), .A3(new_n1281), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n1272), .A2(new_n1273), .B1(new_n1277), .B2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT125), .ZN(new_n1284));
  AND4_X1   g1084(.A1(new_n1284), .A2(new_n1277), .A3(new_n1282), .A4(new_n1273), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1271), .B1(new_n1283), .B2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(G387), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1273), .B1(new_n1287), .B2(new_n1284), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1277), .A2(new_n1282), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1277), .A2(new_n1282), .A3(new_n1284), .A4(new_n1273), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1290), .A2(KEYINPUT126), .A3(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1286), .A2(new_n1292), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1225), .B(G378), .C1(new_n1229), .C2(new_n1235), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1233), .A2(new_n1234), .A3(new_n991), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1196), .A2(new_n1224), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1266), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1294), .A2(new_n1297), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1142), .A2(new_n1144), .A3(KEYINPUT60), .A4(new_n1227), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1299), .A2(new_n668), .A3(new_n1137), .ZN(new_n1300));
  AOI21_X1  g1100(.A(KEYINPUT60), .B1(new_n1237), .B2(new_n1227), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1259), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(G384), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  OAI211_X1 g1104(.A(G384), .B(new_n1259), .C1(new_n1300), .C2(new_n1301), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1298), .A2(new_n1267), .A3(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT62), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1268), .B1(new_n1294), .B2(new_n1297), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1311), .A2(KEYINPUT62), .A3(new_n1307), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1310), .A2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1298), .A2(new_n1267), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1268), .A2(G2897), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1304), .A2(KEYINPUT124), .A3(new_n1305), .A4(new_n1316), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1304), .A2(KEYINPUT124), .A3(new_n1305), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(new_n1315), .ZN(new_n1319));
  AOI21_X1  g1119(.A(KEYINPUT124), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1317), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1121(.A(KEYINPUT61), .B1(new_n1314), .B2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1293), .B1(new_n1313), .B2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1314), .A2(new_n1321), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT61), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1311), .A2(KEYINPUT63), .A3(new_n1307), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1324), .A2(new_n1325), .A3(new_n1326), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1283), .A2(new_n1285), .ZN(new_n1328));
  AOI211_X1 g1128(.A(new_n1268), .B(new_n1306), .C1(new_n1294), .C2(new_n1297), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1328), .B1(new_n1329), .B2(KEYINPUT63), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1327), .A2(new_n1330), .ZN(new_n1331));
  OAI21_X1  g1131(.A(KEYINPUT127), .B1(new_n1323), .B2(new_n1331), .ZN(new_n1332));
  AND3_X1   g1132(.A1(new_n1311), .A2(KEYINPUT62), .A3(new_n1307), .ZN(new_n1333));
  AOI21_X1  g1133(.A(KEYINPUT62), .B1(new_n1311), .B2(new_n1307), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1322), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  AND2_X1   g1135(.A1(new_n1286), .A2(new_n1292), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT127), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT63), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1308), .A2(new_n1339), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1322), .A2(new_n1340), .A3(new_n1328), .A4(new_n1326), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1337), .A2(new_n1338), .A3(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1332), .A2(new_n1342), .ZN(G405));
  NAND2_X1  g1143(.A1(G375), .A2(new_n1266), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1344), .A2(new_n1294), .ZN(new_n1345));
  XNOR2_X1  g1145(.A(new_n1345), .B(new_n1306), .ZN(new_n1346));
  XNOR2_X1  g1146(.A(new_n1346), .B(new_n1328), .ZN(G402));
endmodule


