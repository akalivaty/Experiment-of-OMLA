//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 1 0 0 1 1 0 0 0 1 0 0 0 0 0 1 0 0 0 1 0 0 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 1 1 0 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n794, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n816, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G122), .ZN(new_n189));
  OR2_X1    g003(.A1(KEYINPUT69), .A2(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(KEYINPUT69), .A2(G119), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(G116), .A3(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G116), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G119), .ZN(new_n194));
  INV_X1    g008(.A(G113), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT2), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT2), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G113), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n192), .A2(new_n194), .A3(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT70), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT70), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n192), .A2(new_n199), .A3(new_n202), .A4(new_n194), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n192), .A2(new_n194), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(new_n196), .A3(new_n198), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT4), .ZN(new_n207));
  INV_X1    g021(.A(G101), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT79), .ZN(new_n209));
  INV_X1    g023(.A(G107), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n209), .B1(new_n210), .B2(G104), .ZN(new_n211));
  INV_X1    g025(.A(G104), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(KEYINPUT79), .A3(G107), .ZN(new_n213));
  AND2_X1   g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n215), .B1(new_n212), .B2(G107), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n210), .A2(KEYINPUT3), .A3(G104), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n208), .B1(new_n214), .B2(new_n218), .ZN(new_n219));
  AOI22_X1  g033(.A1(new_n204), .A2(new_n206), .B1(new_n207), .B2(new_n219), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n218), .A2(new_n208), .A3(new_n211), .A4(new_n213), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT80), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n214), .A2(KEYINPUT80), .A3(new_n208), .A4(new_n218), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n219), .A2(new_n207), .ZN(new_n226));
  AND3_X1   g040(.A1(new_n225), .A2(KEYINPUT81), .A3(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(KEYINPUT81), .B1(new_n225), .B2(new_n226), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n220), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n210), .A2(G104), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n212), .A2(G107), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n208), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n232), .B1(new_n223), .B2(new_n224), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT5), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n190), .A2(new_n234), .A3(G116), .A4(new_n191), .ZN(new_n235));
  AND2_X1   g049(.A1(new_n235), .A2(G113), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n192), .A2(KEYINPUT5), .A3(new_n194), .ZN(new_n237));
  AOI22_X1  g051(.A1(new_n201), .A2(new_n203), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n233), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n189), .B1(new_n229), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT6), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT6), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n229), .A2(new_n239), .A3(new_n189), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT85), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT85), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n229), .A2(new_n245), .A3(new_n239), .A4(new_n189), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n242), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n241), .B1(new_n247), .B2(new_n240), .ZN(new_n248));
  INV_X1    g062(.A(G125), .ZN(new_n249));
  INV_X1    g063(.A(G146), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G143), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT1), .ZN(new_n252));
  INV_X1    g066(.A(G143), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G146), .ZN(new_n254));
  AOI22_X1  g068(.A1(new_n252), .A2(G128), .B1(new_n251), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT1), .ZN(new_n256));
  AND4_X1   g070(.A1(new_n256), .A2(new_n251), .A3(new_n254), .A4(G128), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n249), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(G143), .B(G146), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT0), .ZN(new_n260));
  INV_X1    g074(.A(G128), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n251), .A2(new_n254), .ZN(new_n264));
  NOR2_X1   g078(.A1(KEYINPUT0), .A2(G128), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT64), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(KEYINPUT0), .A2(G128), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n269), .B1(new_n265), .B2(new_n266), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n263), .B(G125), .C1(new_n268), .C2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n258), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G224), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n273), .A2(G953), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n274), .B(KEYINPUT86), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n272), .B(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n248), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n244), .A2(new_n246), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT88), .ZN(new_n279));
  XOR2_X1   g093(.A(new_n189), .B(KEYINPUT8), .Z(new_n280));
  INV_X1    g094(.A(new_n232), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n225), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n236), .A2(new_n237), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n204), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n280), .B1(new_n285), .B2(new_n239), .ZN(new_n286));
  OAI21_X1  g100(.A(KEYINPUT7), .B1(new_n273), .B2(G953), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT87), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n272), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n287), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT87), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n272), .A2(new_n291), .A3(new_n290), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n279), .B1(new_n286), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n280), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n233), .A2(new_n238), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n233), .A2(new_n238), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n292), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n301), .B1(new_n272), .B2(new_n288), .ZN(new_n302));
  AOI211_X1 g116(.A(KEYINPUT87), .B(new_n287), .C1(new_n258), .C2(new_n271), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n300), .A2(KEYINPUT88), .A3(new_n304), .ZN(new_n305));
  AND2_X1   g119(.A1(new_n296), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n278), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G902), .ZN(new_n308));
  AOI21_X1  g122(.A(KEYINPUT89), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT89), .ZN(new_n310));
  AOI211_X1 g124(.A(new_n310), .B(G902), .C1(new_n278), .C2(new_n306), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n277), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(G210), .B1(G237), .B2(G902), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n296), .A2(new_n305), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n316), .B1(new_n246), .B2(new_n244), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n310), .B1(new_n317), .B2(G902), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n307), .A2(KEYINPUT89), .A3(new_n308), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(new_n313), .A3(new_n277), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n188), .B1(new_n315), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G217), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n323), .B1(G234), .B2(new_n308), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT69), .B(G119), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G128), .ZN(new_n327));
  OR2_X1    g141(.A1(G119), .A2(G128), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT24), .B(G110), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  OR2_X1    g144(.A1(new_n330), .A2(KEYINPUT78), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(KEYINPUT78), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n326), .A2(new_n261), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT23), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n327), .A2(new_n328), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n335), .B1(new_n336), .B2(new_n334), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n331), .B(new_n332), .C1(new_n337), .C2(G110), .ZN(new_n338));
  NOR3_X1   g152(.A1(new_n249), .A2(KEYINPUT16), .A3(G140), .ZN(new_n339));
  XNOR2_X1  g153(.A(G125), .B(G140), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n339), .B1(new_n340), .B2(KEYINPUT16), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G146), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n250), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n338), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n337), .A2(G110), .ZN(new_n346));
  OR2_X1    g160(.A1(new_n341), .A2(G146), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n342), .ZN(new_n348));
  INV_X1    g162(.A(new_n336), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n346), .B(new_n348), .C1(new_n349), .C2(new_n329), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n345), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(KEYINPUT22), .B(G137), .ZN(new_n352));
  INV_X1    g166(.A(G953), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n353), .A2(G221), .A3(G234), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n352), .B(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n355), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n345), .A2(new_n350), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n356), .A2(new_n308), .A3(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT25), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n356), .A2(KEYINPUT25), .A3(new_n308), .A4(new_n358), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n325), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n345), .A2(new_n350), .A3(new_n357), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n357), .B1(new_n345), .B2(new_n350), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n324), .A2(G902), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(G472), .A2(G902), .ZN(new_n371));
  NOR2_X1   g185(.A1(G237), .A2(G953), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G210), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n373), .B(KEYINPUT27), .ZN(new_n374));
  XNOR2_X1  g188(.A(KEYINPUT26), .B(G101), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n374), .B(new_n375), .ZN(new_n376));
  XOR2_X1   g190(.A(new_n376), .B(KEYINPUT73), .Z(new_n377));
  INV_X1    g191(.A(KEYINPUT66), .ZN(new_n378));
  INV_X1    g192(.A(G137), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n378), .B1(new_n379), .B2(G134), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(G134), .ZN(new_n381));
  INV_X1    g195(.A(G134), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(KEYINPUT66), .A3(G137), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n380), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT67), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n385), .A3(G131), .ZN(new_n386));
  INV_X1    g200(.A(G131), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n382), .A2(G137), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT11), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n389), .B1(G134), .B2(new_n379), .ZN(new_n390));
  NOR3_X1   g204(.A1(new_n382), .A2(KEYINPUT11), .A3(G137), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n387), .B(new_n388), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n386), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n385), .B1(new_n384), .B2(G131), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT68), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n384), .A2(G131), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT67), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT68), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n397), .A2(new_n398), .A3(new_n392), .A4(new_n386), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n259), .A2(new_n256), .A3(G128), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n261), .B1(new_n251), .B2(KEYINPUT1), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n400), .B1(new_n401), .B2(new_n259), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n395), .A2(new_n399), .A3(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n388), .B1(new_n390), .B2(new_n391), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G131), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT65), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n406), .A3(new_n392), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n268), .A2(new_n270), .ZN(new_n408));
  INV_X1    g222(.A(new_n263), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n404), .A2(KEYINPUT65), .A3(G131), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n407), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n403), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n204), .A2(new_n206), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(KEYINPUT74), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n414), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n397), .A2(new_n392), .A3(new_n386), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT71), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n418), .B1(new_n255), .B2(new_n257), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n400), .B(KEYINPUT71), .C1(new_n401), .C2(new_n259), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n416), .B(new_n412), .C1(new_n417), .C2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n415), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n416), .B1(new_n403), .B2(new_n412), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n424), .A2(KEYINPUT74), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT28), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT28), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n377), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  OR2_X1    g243(.A1(KEYINPUT72), .A2(KEYINPUT31), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n407), .A2(new_n410), .A3(new_n411), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n421), .A2(new_n417), .ZN(new_n432));
  OAI21_X1  g246(.A(KEYINPUT30), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT30), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n403), .A2(new_n434), .A3(new_n412), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n416), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n422), .A2(new_n376), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n430), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n433), .A2(new_n435), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n414), .ZN(new_n440));
  INV_X1    g254(.A(new_n437), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  XOR2_X1   g256(.A(KEYINPUT72), .B(KEYINPUT31), .Z(new_n443));
  OAI21_X1  g257(.A(new_n438), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n371), .B1(new_n429), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(KEYINPUT32), .ZN(new_n446));
  NOR3_X1   g260(.A1(new_n436), .A2(new_n437), .A3(new_n443), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n447), .B1(new_n442), .B2(new_n430), .ZN(new_n448));
  INV_X1    g262(.A(new_n377), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n431), .A2(new_n432), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n424), .A2(KEYINPUT74), .B1(new_n450), .B2(new_n416), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n413), .A2(new_n414), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT74), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n427), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n428), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n449), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n448), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT32), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(new_n459), .A3(new_n371), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n446), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n414), .B1(new_n431), .B2(new_n432), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT76), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n462), .A2(new_n422), .A3(new_n463), .ZN(new_n464));
  OAI211_X1 g278(.A(KEYINPUT76), .B(new_n414), .C1(new_n431), .C2(new_n432), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n464), .A2(KEYINPUT28), .A3(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT77), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n466), .A2(new_n467), .A3(new_n428), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n464), .A2(KEYINPUT77), .A3(KEYINPUT28), .A4(new_n465), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n376), .A2(KEYINPUT29), .ZN(new_n471));
  AOI21_X1  g285(.A(G902), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n426), .A2(KEYINPUT75), .A3(new_n428), .A4(new_n377), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT75), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n428), .A2(new_n377), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n474), .B1(new_n455), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n440), .A2(new_n422), .ZN(new_n477));
  INV_X1    g291(.A(new_n376), .ZN(new_n478));
  AOI21_X1  g292(.A(KEYINPUT29), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n473), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n472), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(G472), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n370), .B1(new_n461), .B2(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT9), .B(G234), .ZN(new_n484));
  OAI21_X1  g298(.A(G221), .B1(new_n484), .B2(G902), .ZN(new_n485));
  INV_X1    g299(.A(G469), .ZN(new_n486));
  XNOR2_X1  g300(.A(G110), .B(G140), .ZN(new_n487));
  INV_X1    g301(.A(G227), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n488), .A2(G953), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n487), .B(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT12), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n407), .A2(new_n411), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT82), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n251), .A2(new_n495), .A3(KEYINPUT1), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(G128), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n495), .B1(new_n251), .B2(KEYINPUT1), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n264), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n400), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n225), .A2(new_n281), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n402), .B1(new_n225), .B2(new_n281), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n492), .B(new_n494), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n225), .A2(new_n281), .A3(new_n500), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n505), .B1(new_n402), .B2(new_n233), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n492), .B1(new_n506), .B2(new_n494), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n219), .A2(new_n207), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n410), .B(new_n509), .C1(new_n227), .C2(new_n228), .ZN(new_n510));
  XOR2_X1   g324(.A(KEYINPUT83), .B(KEYINPUT10), .Z(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n419), .A2(new_n420), .A3(KEYINPUT10), .ZN(new_n513));
  AOI22_X1  g327(.A1(new_n505), .A2(new_n512), .B1(new_n513), .B2(new_n233), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n510), .A2(new_n493), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n491), .B1(new_n508), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n410), .A2(new_n509), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n225), .A2(new_n226), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT81), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n225), .A2(new_n226), .A3(KEYINPUT81), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n517), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n513), .A2(new_n233), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n523), .B1(new_n501), .B2(new_n511), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n494), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n525), .A2(new_n515), .A3(new_n491), .ZN(new_n526));
  OAI21_X1  g340(.A(KEYINPUT84), .B1(new_n516), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n506), .A2(new_n494), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(KEYINPUT12), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n515), .A2(new_n529), .A3(new_n503), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n490), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT84), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n525), .A2(new_n515), .A3(new_n491), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n486), .B1(new_n527), .B2(new_n534), .ZN(new_n535));
  AND4_X1   g349(.A1(new_n515), .A2(new_n529), .A3(new_n503), .A4(new_n491), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n491), .B1(new_n525), .B2(new_n515), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n486), .B(new_n308), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(G469), .A2(G902), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n485), .B1(new_n535), .B2(new_n540), .ZN(new_n541));
  OR2_X1    g355(.A1(KEYINPUT96), .A2(KEYINPUT13), .ZN(new_n542));
  NAND2_X1  g356(.A1(KEYINPUT96), .A2(KEYINPUT13), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n253), .A2(G128), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n544), .A2(KEYINPUT97), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n261), .A2(G143), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n542), .A2(new_n545), .A3(new_n543), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(KEYINPUT97), .B1(new_n544), .B2(new_n546), .ZN(new_n551));
  OAI21_X1  g365(.A(G134), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n545), .A2(new_n548), .A3(new_n382), .ZN(new_n553));
  INV_X1    g367(.A(G122), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(G116), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n193), .A2(G122), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(G107), .ZN(new_n558));
  XNOR2_X1  g372(.A(G116), .B(G122), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n210), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n552), .A2(new_n553), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n545), .A2(new_n548), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(G134), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n553), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT98), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n560), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n193), .A2(KEYINPUT14), .A3(G122), .ZN(new_n568));
  OAI211_X1 g382(.A(G107), .B(new_n568), .C1(new_n557), .C2(KEYINPUT14), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n559), .A2(KEYINPUT98), .A3(new_n210), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n565), .A2(new_n567), .A3(new_n569), .A4(new_n570), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n484), .A2(new_n323), .A3(G953), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n562), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n572), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n561), .A2(new_n553), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n544), .A2(new_n546), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT97), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n578), .A2(new_n547), .A3(new_n548), .A4(new_n549), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n575), .B1(new_n579), .B2(G134), .ZN(new_n580));
  INV_X1    g394(.A(new_n571), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n574), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n573), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n308), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT100), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n584), .B(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(G478), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT15), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n587), .B1(KEYINPUT99), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n589), .B1(KEYINPUT99), .B2(new_n588), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n586), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n584), .A2(new_n585), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n590), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT95), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n372), .A2(G143), .A3(G214), .ZN(new_n597));
  AOI21_X1  g411(.A(G143), .B1(new_n372), .B2(G214), .ZN(new_n598));
  OAI21_X1  g412(.A(G131), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n372), .A2(G214), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n253), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n372), .A2(G143), .A3(G214), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n601), .A2(new_n387), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT17), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n599), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  OAI211_X1 g419(.A(KEYINPUT17), .B(G131), .C1(new_n597), .C2(new_n598), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n605), .A2(new_n347), .A3(new_n342), .A4(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(G113), .B(G122), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(new_n212), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n597), .A2(new_n598), .ZN(new_n610));
  NAND2_X1  g424(.A1(KEYINPUT18), .A2(G131), .ZN(new_n611));
  OR2_X1    g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(G140), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(G125), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n249), .A2(G140), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(G146), .ZN(new_n617));
  AOI22_X1  g431(.A1(new_n610), .A2(new_n611), .B1(new_n617), .B2(new_n343), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n612), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n607), .A2(new_n609), .A3(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n609), .B1(new_n607), .B2(new_n619), .ZN(new_n622));
  OAI211_X1 g436(.A(KEYINPUT94), .B(new_n308), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(G475), .ZN(new_n624));
  INV_X1    g438(.A(new_n622), .ZN(new_n625));
  AOI21_X1  g439(.A(G902), .B1(new_n625), .B2(new_n620), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n626), .A2(KEYINPUT94), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT91), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n628), .B1(new_n616), .B2(KEYINPUT19), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT19), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n340), .A2(KEYINPUT91), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT90), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n633), .B1(new_n340), .B2(new_n630), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n616), .A2(KEYINPUT90), .A3(KEYINPUT19), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n632), .A2(new_n636), .A3(new_n250), .ZN(new_n637));
  AOI22_X1  g451(.A1(new_n599), .A2(new_n603), .B1(new_n341), .B2(G146), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n619), .ZN(new_n640));
  INV_X1    g454(.A(new_n609), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n640), .A2(KEYINPUT92), .A3(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT92), .ZN(new_n643));
  AOI22_X1  g457(.A1(new_n637), .A2(new_n638), .B1(new_n612), .B2(new_n618), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n643), .B1(new_n644), .B2(new_n609), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n642), .A2(new_n645), .A3(new_n620), .ZN(new_n646));
  NOR2_X1   g460(.A1(G475), .A2(G902), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT93), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n647), .B1(new_n648), .B2(KEYINPUT20), .ZN(new_n649));
  OAI21_X1  g463(.A(KEYINPUT93), .B1(G475), .B2(G902), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n646), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT20), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n654), .B1(new_n646), .B2(new_n647), .ZN(new_n655));
  OAI221_X1 g469(.A(new_n596), .B1(new_n624), .B2(new_n627), .C1(new_n653), .C2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n627), .A2(new_n624), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n646), .A2(new_n647), .ZN(new_n658));
  AOI22_X1  g472(.A1(new_n658), .A2(KEYINPUT20), .B1(new_n646), .B2(new_n651), .ZN(new_n659));
  OAI21_X1  g473(.A(KEYINPUT95), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(G952), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n661), .A2(G953), .ZN(new_n662));
  INV_X1    g476(.A(G234), .ZN(new_n663));
  INV_X1    g477(.A(G237), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  AOI211_X1 g480(.A(new_n308), .B(new_n353), .C1(G234), .C2(G237), .ZN(new_n667));
  XNOR2_X1  g481(.A(KEYINPUT21), .B(G898), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n595), .A2(new_n656), .A3(new_n660), .A4(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n541), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n322), .A2(new_n483), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G101), .ZN(G3));
  INV_X1    g488(.A(KEYINPUT101), .ZN(new_n675));
  AOI221_X4 g489(.A(new_n314), .B1(new_n248), .B2(new_n276), .C1(new_n318), .C2(new_n319), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n313), .B1(new_n320), .B2(new_n277), .ZN(new_n677));
  OAI211_X1 g491(.A(new_n187), .B(new_n670), .C1(new_n676), .C2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n584), .A2(G478), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n587), .A2(new_n308), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n583), .B(KEYINPUT33), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n681), .B1(new_n682), .B2(new_n587), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n683), .B1(new_n656), .B2(new_n660), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n675), .B1(new_n678), .B2(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n322), .A2(KEYINPUT101), .A3(new_n670), .A4(new_n684), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OAI211_X1 g502(.A(new_n369), .B(new_n485), .C1(new_n535), .C2(new_n540), .ZN(new_n689));
  AOI21_X1  g503(.A(G902), .B1(new_n448), .B2(new_n457), .ZN(new_n690));
  INV_X1    g504(.A(G472), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n445), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n688), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT34), .B(G104), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G6));
  INV_X1    g510(.A(KEYINPUT102), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n655), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n658), .A2(KEYINPUT20), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n592), .A2(new_n594), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n702), .A2(new_n657), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n322), .A2(new_n670), .A3(new_n703), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n704), .A2(new_n692), .A3(new_n689), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT35), .B(G107), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G9));
  NAND2_X1  g521(.A1(new_n315), .A2(new_n321), .ZN(new_n708));
  AOI21_X1  g522(.A(KEYINPUT25), .B1(new_n366), .B2(new_n308), .ZN(new_n709));
  INV_X1    g523(.A(new_n362), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n324), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n355), .A2(KEYINPUT36), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n345), .A2(new_n350), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n712), .B1(new_n345), .B2(new_n350), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT103), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n715), .A2(new_n716), .A3(new_n367), .ZN(new_n717));
  INV_X1    g531(.A(new_n712), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n351), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n345), .A2(new_n350), .A3(new_n712), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n719), .A2(new_n367), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(KEYINPUT103), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n717), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n711), .A2(new_n723), .ZN(new_n724));
  OAI211_X1 g538(.A(new_n724), .B(new_n445), .C1(new_n690), .C2(new_n691), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n708), .A2(new_n672), .A3(new_n187), .A4(new_n726), .ZN(new_n727));
  XOR2_X1   g541(.A(KEYINPUT37), .B(G110), .Z(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G12));
  INV_X1    g543(.A(G900), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n666), .B1(new_n667), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n657), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n700), .A2(new_n724), .A3(new_n701), .A4(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n541), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n461), .A2(new_n482), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n708), .A2(new_n734), .A3(new_n735), .A4(new_n187), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G128), .ZN(G30));
  XNOR2_X1  g551(.A(new_n708), .B(KEYINPUT38), .ZN(new_n738));
  XOR2_X1   g552(.A(new_n731), .B(KEYINPUT39), .Z(new_n739));
  OAI211_X1 g553(.A(new_n485), .B(new_n739), .C1(new_n535), .C2(new_n540), .ZN(new_n740));
  OR2_X1    g554(.A1(new_n740), .A2(KEYINPUT40), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n656), .A2(new_n660), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n743), .A2(new_n595), .ZN(new_n744));
  INV_X1    g558(.A(new_n724), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n744), .A2(new_n187), .A3(new_n745), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n746), .B1(new_n740), .B2(KEYINPUT40), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n449), .A2(new_n465), .A3(new_n464), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n442), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n691), .B1(new_n749), .B2(new_n308), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n750), .B1(new_n446), .B2(new_n460), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n738), .A2(new_n741), .A3(new_n747), .A4(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G143), .ZN(G45));
  OAI211_X1 g568(.A(new_n485), .B(new_n724), .C1(new_n535), .C2(new_n540), .ZN(new_n755));
  INV_X1    g569(.A(new_n731), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n684), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n758), .A2(new_n708), .A3(new_n735), .A4(new_n187), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G146), .ZN(G48));
  NOR3_X1   g574(.A1(new_n522), .A2(new_n524), .A3(new_n494), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n493), .B1(new_n510), .B2(new_n514), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n490), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n763), .B1(new_n530), .B2(new_n490), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n308), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(G469), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n766), .A2(new_n485), .A3(new_n538), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n483), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n768), .B1(new_n686), .B2(new_n687), .ZN(new_n769));
  XOR2_X1   g583(.A(KEYINPUT41), .B(G113), .Z(new_n770));
  XNOR2_X1  g584(.A(new_n769), .B(new_n770), .ZN(G15));
  NOR2_X1   g585(.A1(new_n704), .A2(new_n768), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(new_n193), .ZN(G18));
  INV_X1    g587(.A(new_n671), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n735), .A2(new_n774), .A3(new_n724), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n187), .B(new_n767), .C1(new_n676), .C2(new_n677), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT104), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n322), .A2(KEYINPUT104), .A3(new_n767), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n775), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  XOR2_X1   g594(.A(KEYINPUT105), .B(G119), .Z(new_n781));
  XNOR2_X1  g595(.A(new_n780), .B(new_n781), .ZN(G21));
  NAND2_X1  g596(.A1(new_n458), .A2(new_n308), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(G472), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n448), .B1(new_n470), .B2(new_n377), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n371), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n784), .A2(new_n369), .A3(new_n786), .ZN(new_n787));
  AND4_X1   g601(.A1(new_n670), .A2(new_n766), .A3(new_n485), .A4(new_n538), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n322), .A2(new_n744), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G122), .ZN(G24));
  NAND3_X1  g604(.A1(new_n784), .A2(new_n724), .A3(new_n786), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(new_n757), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n793), .B1(new_n778), .B2(new_n779), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(new_n249), .ZN(G27));
  AND3_X1   g609(.A1(new_n315), .A2(new_n187), .A3(new_n321), .ZN(new_n796));
  INV_X1    g610(.A(new_n757), .ZN(new_n797));
  INV_X1    g611(.A(new_n485), .ZN(new_n798));
  XOR2_X1   g612(.A(new_n539), .B(KEYINPUT106), .Z(new_n799));
  AND2_X1   g613(.A1(new_n538), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT107), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n801), .B1(new_n530), .B2(new_n490), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n530), .A2(new_n801), .A3(new_n490), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n803), .A2(G469), .A3(new_n533), .A4(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n798), .B1(new_n800), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n796), .A2(new_n483), .A3(new_n797), .A4(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT42), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n735), .A2(new_n369), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n315), .A2(new_n806), .A3(new_n187), .A4(new_n321), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n812), .A2(KEYINPUT42), .A3(new_n797), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G131), .ZN(G33));
  NOR3_X1   g629(.A1(new_n702), .A2(new_n657), .A3(new_n731), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n796), .A2(new_n483), .A3(new_n816), .A4(new_n806), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G134), .ZN(G36));
  INV_X1    g632(.A(new_n683), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n819), .A2(new_n660), .A3(new_n656), .ZN(new_n820));
  XOR2_X1   g634(.A(new_n820), .B(KEYINPUT43), .Z(new_n821));
  NAND3_X1  g635(.A1(new_n821), .A2(new_n692), .A3(new_n724), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT44), .ZN(new_n823));
  OR2_X1    g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n796), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n825), .B1(new_n822), .B2(new_n823), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT109), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT109), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n824), .A2(new_n829), .A3(new_n826), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT46), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n527), .A2(new_n534), .ZN(new_n833));
  OAI21_X1  g647(.A(G469), .B1(new_n833), .B2(KEYINPUT45), .ZN(new_n834));
  OR2_X1    g648(.A1(new_n834), .A2(KEYINPUT108), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n804), .A2(new_n533), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n836), .A2(new_n802), .ZN(new_n837));
  AOI22_X1  g651(.A1(new_n834), .A2(KEYINPUT108), .B1(KEYINPUT45), .B2(new_n837), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n799), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n832), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n538), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n839), .A2(new_n832), .A3(new_n840), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n485), .B(new_n739), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n831), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(new_n379), .ZN(G39));
  OAI21_X1  g660(.A(new_n485), .B1(new_n842), .B2(new_n843), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT47), .ZN(new_n848));
  OR2_X1    g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n847), .A2(new_n848), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n461), .A2(new_n482), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n825), .A2(new_n369), .A3(new_n757), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(G140), .ZN(G42));
  AND2_X1   g669(.A1(new_n766), .A2(new_n538), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(KEYINPUT49), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n820), .A2(new_n188), .A3(new_n798), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OR4_X1    g673(.A1(new_n370), .A2(new_n738), .A3(new_n859), .A4(new_n752), .ZN(new_n860));
  INV_X1    g674(.A(new_n767), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n825), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(KEYINPUT115), .ZN(new_n863));
  INV_X1    g677(.A(new_n791), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n821), .A2(new_n666), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT114), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n821), .A2(KEYINPUT114), .A3(new_n666), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n863), .A2(new_n864), .A3(new_n869), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n752), .A2(new_n370), .A3(new_n665), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n863), .A2(new_n743), .A3(new_n683), .A4(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n869), .A2(new_n787), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n738), .A2(new_n187), .A3(new_n861), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n874), .A2(new_n875), .A3(KEYINPUT50), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT50), .B1(new_n874), .B2(new_n875), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n870), .B(new_n872), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(KEYINPUT116), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n872), .A2(new_n870), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT116), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n881), .B(new_n882), .C1(new_n878), .C2(new_n877), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n856), .A2(new_n798), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n849), .A2(new_n850), .A3(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n873), .A2(new_n825), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n880), .A2(new_n883), .A3(KEYINPUT51), .A4(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT104), .B1(new_n322), .B2(new_n767), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n776), .A2(new_n777), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n874), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n863), .A2(new_n684), .A3(new_n871), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n891), .A2(new_n662), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n863), .A2(new_n869), .ZN(new_n894));
  OR3_X1    g708(.A1(new_n894), .A2(KEYINPUT48), .A3(new_n810), .ZN(new_n895));
  OAI21_X1  g709(.A(KEYINPUT48), .B1(new_n894), .B2(new_n810), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n893), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n879), .B1(new_n885), .B2(new_n886), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n888), .B(new_n897), .C1(KEYINPUT51), .C2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n796), .A2(new_n792), .A3(new_n806), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n817), .A2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n676), .A2(new_n677), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT110), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n595), .A2(new_n700), .A3(new_n732), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n903), .A2(new_n904), .A3(new_n187), .A4(new_n905), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n315), .A2(new_n905), .A3(new_n187), .A4(new_n321), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(KEYINPUT110), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n852), .A2(new_n755), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n906), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n701), .A2(new_n656), .A3(new_n660), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n669), .B1(new_n685), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n322), .A2(new_n693), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n673), .A2(new_n913), .A3(new_n727), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n814), .A2(new_n902), .A3(new_n910), .A4(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n768), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n688), .A2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n780), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n789), .B1(new_n704), .B2(new_n768), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n916), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n792), .B1(new_n890), .B2(new_n889), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n717), .A2(new_n722), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n363), .A2(new_n925), .A3(new_n731), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n836), .A2(new_n486), .A3(new_n802), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n538), .A2(new_n799), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n926), .B(new_n485), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n751), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n322), .A2(new_n930), .A3(new_n744), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n931), .A2(new_n759), .A3(new_n736), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT52), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n924), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n931), .A2(new_n759), .A3(new_n736), .ZN(new_n935));
  OAI21_X1  g749(.A(KEYINPUT52), .B1(new_n794), .B2(new_n935), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n934), .A2(new_n936), .A3(KEYINPUT53), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n923), .A2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT53), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n933), .B1(new_n924), .B2(new_n932), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n794), .A2(new_n935), .A3(KEYINPUT52), .ZN(new_n941));
  OAI21_X1  g755(.A(KEYINPUT112), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT112), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n934), .A2(new_n936), .A3(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n923), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n938), .B1(new_n939), .B2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT113), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT54), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n945), .A2(new_n939), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n923), .A2(new_n937), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n950), .A2(new_n948), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(KEYINPUT113), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n945), .A2(KEYINPUT53), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n923), .A2(KEYINPUT111), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n940), .A2(new_n941), .A3(KEYINPUT53), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(new_n923), .B2(KEYINPUT111), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n954), .B(KEYINPUT54), .C1(new_n956), .C2(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n949), .A2(new_n953), .A3(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n899), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g775(.A1(G952), .A2(G953), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n860), .B1(new_n961), .B2(new_n962), .ZN(G75));
  NAND2_X1  g777(.A1(new_n661), .A2(G953), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT117), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n950), .A2(new_n951), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n967), .A2(G210), .A3(G902), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n248), .B(new_n276), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT55), .Z(new_n970));
  OR3_X1    g784(.A1(new_n968), .A2(KEYINPUT56), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n970), .B1(new_n968), .B2(KEYINPUT56), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n966), .B1(new_n971), .B2(new_n972), .ZN(G51));
  NOR3_X1   g787(.A1(new_n769), .A2(new_n780), .A3(new_n920), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n906), .A2(new_n908), .A3(new_n909), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n975), .A2(new_n901), .A3(new_n914), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n974), .A2(new_n976), .A3(new_n814), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n943), .B1(new_n934), .B2(new_n936), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(KEYINPUT53), .B1(new_n979), .B2(new_n944), .ZN(new_n980));
  OAI21_X1  g794(.A(KEYINPUT54), .B1(new_n980), .B2(new_n938), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n952), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n799), .B(KEYINPUT57), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n764), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n946), .A2(new_n308), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(new_n839), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n966), .B1(new_n985), .B2(new_n987), .ZN(G54));
  NAND2_X1  g802(.A1(KEYINPUT58), .A2(G475), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT118), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n989), .B(new_n990), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n986), .A2(new_n646), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n646), .B1(new_n986), .B2(new_n991), .ZN(new_n993));
  NOR3_X1   g807(.A1(new_n992), .A2(new_n993), .A3(new_n966), .ZN(G60));
  XOR2_X1   g808(.A(new_n680), .B(KEYINPUT59), .Z(new_n995));
  NAND2_X1  g809(.A1(new_n682), .A2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(KEYINPUT119), .B1(new_n982), .B2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT119), .ZN(new_n999));
  AOI211_X1 g813(.A(new_n999), .B(new_n996), .C1(new_n981), .C2(new_n952), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n965), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n682), .B1(new_n960), .B2(new_n995), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n1001), .A2(new_n1002), .ZN(G63));
  NAND2_X1  g817(.A1(G217), .A2(G902), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1004), .B(KEYINPUT60), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n967), .A2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n366), .B(KEYINPUT122), .Z(new_n1008));
  AOI21_X1  g822(.A(new_n966), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n946), .A2(new_n1005), .ZN(new_n1010));
  AOI21_X1  g824(.A(KEYINPUT121), .B1(new_n1010), .B2(new_n715), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n967), .A2(new_n715), .A3(new_n1006), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT121), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g828(.A(KEYINPUT61), .B(new_n1009), .C1(new_n1011), .C2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1008), .B1(new_n946), .B2(new_n1005), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(new_n965), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1010), .A2(KEYINPUT121), .A3(new_n715), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g834(.A(KEYINPUT120), .B(KEYINPUT61), .Z(new_n1021));
  OAI21_X1  g835(.A(new_n1015), .B1(new_n1020), .B2(new_n1021), .ZN(G66));
  OAI21_X1  g836(.A(G953), .B1(new_n668), .B2(new_n273), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n922), .A2(new_n914), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1023), .B1(new_n1024), .B2(G953), .ZN(new_n1025));
  INV_X1    g839(.A(new_n248), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1026), .B1(G898), .B2(new_n353), .ZN(new_n1027));
  XNOR2_X1  g841(.A(new_n1025), .B(new_n1027), .ZN(G69));
  NAND2_X1  g842(.A1(new_n632), .A2(new_n636), .ZN(new_n1029));
  XNOR2_X1  g843(.A(new_n1029), .B(KEYINPUT123), .ZN(new_n1030));
  XNOR2_X1  g844(.A(new_n439), .B(new_n1030), .ZN(new_n1031));
  INV_X1    g845(.A(new_n1031), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n322), .A2(new_n483), .A3(new_n744), .ZN(new_n1033));
  OR2_X1    g847(.A1(new_n844), .A2(new_n1033), .ZN(new_n1034));
  AND3_X1   g848(.A1(new_n924), .A2(new_n736), .A3(new_n759), .ZN(new_n1035));
  OAI211_X1 g849(.A(new_n1034), .B(new_n1035), .C1(new_n844), .C2(new_n831), .ZN(new_n1036));
  INV_X1    g850(.A(new_n1036), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n814), .A2(new_n817), .ZN(new_n1038));
  XNOR2_X1  g852(.A(new_n1038), .B(KEYINPUT125), .ZN(new_n1039));
  NAND4_X1  g853(.A1(new_n1037), .A2(new_n353), .A3(new_n854), .A4(new_n1039), .ZN(new_n1040));
  NAND2_X1  g854(.A1(G900), .A2(G953), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n1032), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g856(.A(KEYINPUT62), .ZN(new_n1043));
  AOI21_X1  g857(.A(new_n1043), .B1(new_n1035), .B2(new_n753), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n684), .B1(new_n743), .B2(new_n701), .ZN(new_n1045));
  NOR4_X1   g859(.A1(new_n825), .A2(new_n810), .A3(new_n740), .A4(new_n1045), .ZN(new_n1046));
  NOR3_X1   g860(.A1(new_n845), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n1035), .A2(new_n1043), .A3(new_n753), .ZN(new_n1048));
  XNOR2_X1  g862(.A(new_n1048), .B(KEYINPUT124), .ZN(new_n1049));
  NAND3_X1  g863(.A1(new_n1047), .A2(new_n1049), .A3(new_n854), .ZN(new_n1050));
  NOR2_X1   g864(.A1(new_n1031), .A2(G953), .ZN(new_n1051));
  AND2_X1   g865(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g866(.A(new_n353), .B1(G227), .B2(G900), .ZN(new_n1053));
  XNOR2_X1  g867(.A(new_n1053), .B(KEYINPUT126), .ZN(new_n1054));
  OR3_X1    g868(.A1(new_n1042), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  OAI21_X1  g869(.A(new_n1054), .B1(new_n1042), .B2(new_n1052), .ZN(new_n1056));
  NAND2_X1  g870(.A1(new_n1055), .A2(new_n1056), .ZN(G72));
  NAND2_X1  g871(.A1(new_n477), .A2(new_n376), .ZN(new_n1058));
  NAND4_X1  g872(.A1(new_n1047), .A2(new_n854), .A3(new_n1024), .A4(new_n1049), .ZN(new_n1059));
  NAND2_X1  g873(.A1(G472), .A2(G902), .ZN(new_n1060));
  XOR2_X1   g874(.A(new_n1060), .B(KEYINPUT63), .Z(new_n1061));
  NAND2_X1  g875(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g876(.A1(new_n1062), .A2(KEYINPUT127), .ZN(new_n1063));
  INV_X1    g877(.A(KEYINPUT127), .ZN(new_n1064));
  NAND3_X1  g878(.A1(new_n1059), .A2(new_n1064), .A3(new_n1061), .ZN(new_n1065));
  AOI21_X1  g879(.A(new_n1058), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g880(.A(new_n1061), .ZN(new_n1067));
  NAND2_X1  g881(.A1(new_n477), .A2(new_n478), .ZN(new_n1068));
  AOI21_X1  g882(.A(new_n1067), .B1(new_n1068), .B2(new_n442), .ZN(new_n1069));
  OAI211_X1 g883(.A(new_n954), .B(new_n1069), .C1(new_n958), .C2(new_n956), .ZN(new_n1070));
  NAND4_X1  g884(.A1(new_n1037), .A2(new_n854), .A3(new_n1024), .A4(new_n1039), .ZN(new_n1071));
  AND2_X1   g885(.A1(new_n1071), .A2(new_n1061), .ZN(new_n1072));
  NAND3_X1  g886(.A1(new_n440), .A2(new_n422), .A3(new_n478), .ZN(new_n1073));
  OAI211_X1 g887(.A(new_n965), .B(new_n1070), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g888(.A1(new_n1066), .A2(new_n1074), .ZN(G57));
endmodule


