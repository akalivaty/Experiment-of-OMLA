//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 1 0 1 1 0 1 1 0 1 1 1 0 0 0 1 1 0 0 0 0 1 0 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 1 0 1 1 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:14 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(KEYINPUT1), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  AND3_X1   g006(.A1(new_n188), .A2(new_n190), .A3(new_n192), .ZN(new_n193));
  AOI21_X1  g007(.A(G128), .B1(new_n190), .B2(new_n192), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n189), .A2(KEYINPUT1), .A3(G146), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  NOR3_X1   g010(.A1(new_n193), .A2(new_n194), .A3(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G134), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G137), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n198), .A2(G137), .ZN(new_n201));
  OAI21_X1  g015(.A(G131), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT11), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n203), .B1(new_n198), .B2(G137), .ZN(new_n204));
  INV_X1    g018(.A(G137), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(KEYINPUT11), .A3(G134), .ZN(new_n206));
  INV_X1    g020(.A(G131), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n204), .A2(new_n206), .A3(new_n207), .A4(new_n199), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n202), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT66), .B1(new_n197), .B2(new_n209), .ZN(new_n210));
  AND2_X1   g024(.A1(new_n202), .A2(new_n208), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n188), .A2(new_n190), .A3(new_n192), .ZN(new_n213));
  XNOR2_X1  g027(.A(G143), .B(G146), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n213), .B(new_n195), .C1(G128), .C2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n211), .A2(new_n212), .A3(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n204), .A2(new_n199), .A3(new_n206), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G131), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(new_n208), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n190), .A2(new_n192), .ZN(new_n220));
  NAND2_X1  g034(.A1(KEYINPUT0), .A2(G128), .ZN(new_n221));
  NOR2_X1   g035(.A1(KEYINPUT0), .A2(G128), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT64), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n220), .A2(new_n221), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  AND2_X1   g040(.A1(KEYINPUT0), .A2(G128), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n190), .A2(new_n192), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT65), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n190), .A2(new_n192), .B1(new_n222), .B2(new_n223), .ZN(new_n231));
  AND2_X1   g045(.A1(new_n225), .A2(new_n221), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(KEYINPUT65), .A3(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n219), .A2(new_n230), .A3(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n210), .A2(new_n216), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT30), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n238));
  INV_X1    g052(.A(G116), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n238), .B1(new_n239), .B2(G119), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(G119), .ZN(new_n241));
  INV_X1    g055(.A(G119), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(KEYINPUT67), .A3(G116), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n240), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT2), .B(G113), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n247), .B(new_n248), .C1(new_n244), .C2(new_n245), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G113), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT2), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT2), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G113), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n255), .A2(new_n241), .A3(new_n240), .A4(new_n243), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n248), .B1(new_n256), .B2(new_n247), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n246), .B1(new_n250), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n247), .B1(new_n244), .B2(new_n245), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT69), .ZN(new_n260));
  INV_X1    g074(.A(new_n246), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(new_n261), .A3(new_n249), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  AND3_X1   g077(.A1(new_n231), .A2(KEYINPUT65), .A3(new_n232), .ZN(new_n264));
  AOI22_X1  g078(.A1(new_n231), .A2(new_n232), .B1(new_n228), .B2(KEYINPUT65), .ZN(new_n265));
  OAI21_X1  g079(.A(KEYINPUT70), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n230), .A2(new_n267), .A3(new_n233), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n266), .A2(new_n219), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT71), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n215), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n194), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n272), .A2(KEYINPUT71), .A3(new_n195), .A4(new_n213), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n211), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n269), .A2(new_n275), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n237), .B(new_n263), .C1(new_n276), .C2(new_n236), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n269), .A2(new_n262), .A3(new_n275), .A4(new_n258), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G237), .ZN(new_n280));
  INV_X1    g094(.A(G953), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n281), .A3(G210), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n282), .B(G101), .ZN(new_n283));
  XNOR2_X1  g097(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n283), .B(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT29), .B1(new_n279), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n276), .A2(KEYINPUT74), .ZN(new_n288));
  INV_X1    g102(.A(new_n263), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT74), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n269), .A2(new_n290), .A3(new_n275), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n288), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT28), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n263), .A2(KEYINPUT73), .A3(new_n235), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n278), .ZN(new_n296));
  AOI21_X1  g110(.A(KEYINPUT73), .B1(new_n263), .B2(new_n235), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT28), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n287), .B1(new_n299), .B2(new_n286), .ZN(new_n300));
  INV_X1    g114(.A(G902), .ZN(new_n301));
  INV_X1    g115(.A(new_n278), .ZN(new_n302));
  AOI22_X1  g116(.A1(new_n269), .A2(new_n275), .B1(new_n262), .B2(new_n258), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT28), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n294), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n285), .A2(KEYINPUT29), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n300), .B(new_n301), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G472), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT32), .ZN(new_n309));
  NOR2_X1   g123(.A1(G472), .A2(G902), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n278), .A2(new_n285), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT72), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT72), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n278), .A2(new_n313), .A3(new_n285), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n312), .A2(new_n277), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT31), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT31), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n312), .A2(new_n317), .A3(new_n277), .A4(new_n314), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n285), .B1(new_n294), .B2(new_n298), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n309), .B(new_n310), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n299), .A2(new_n286), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(new_n316), .A3(new_n318), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n309), .B1(new_n324), .B2(new_n310), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n308), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT79), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n187), .A2(KEYINPUT23), .A3(G119), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n328), .B(KEYINPUT75), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT23), .B1(new_n187), .B2(G119), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(KEYINPUT76), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n187), .A2(G119), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n242), .A2(G128), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(new_n334), .A3(KEYINPUT23), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n331), .A2(new_n332), .A3(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G110), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n329), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n332), .A2(new_n333), .ZN(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT24), .B(G110), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G125), .ZN(new_n343));
  NOR3_X1   g157(.A1(new_n343), .A2(KEYINPUT16), .A3(G140), .ZN(new_n344));
  XNOR2_X1  g158(.A(G125), .B(G140), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n344), .B1(new_n345), .B2(KEYINPUT16), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G146), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n191), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n342), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n329), .A2(new_n336), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G110), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT16), .ZN(new_n353));
  OR2_X1    g167(.A1(G125), .A2(G140), .ZN(new_n354));
  NAND2_X1  g168(.A1(G125), .A2(G140), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n191), .B1(new_n356), .B2(new_n344), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n347), .A2(new_n357), .ZN(new_n358));
  OR2_X1    g172(.A1(new_n339), .A2(new_n340), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n352), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(KEYINPUT22), .B(G137), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n281), .A2(G221), .A3(G234), .ZN(new_n362));
  OR2_X1    g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n362), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AND3_X1   g179(.A1(new_n350), .A2(new_n360), .A3(new_n365), .ZN(new_n366));
  AND3_X1   g180(.A1(new_n363), .A2(new_n364), .A3(KEYINPUT77), .ZN(new_n367));
  AOI21_X1  g181(.A(KEYINPUT77), .B1(new_n363), .B2(new_n364), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n369), .B1(new_n350), .B2(new_n360), .ZN(new_n370));
  OR2_X1    g184(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G217), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n372), .B1(G234), .B2(new_n301), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n373), .A2(G902), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n375), .A2(KEYINPUT78), .ZN(new_n376));
  AOI21_X1  g190(.A(KEYINPUT78), .B1(new_n371), .B2(new_n374), .ZN(new_n377));
  OR2_X1    g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n301), .B1(new_n366), .B2(new_n370), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT25), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT25), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n381), .B(new_n301), .C1(new_n366), .C2(new_n370), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n380), .A2(new_n373), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n327), .B1(new_n378), .B2(new_n384), .ZN(new_n385));
  OR4_X1    g199(.A1(new_n327), .A2(new_n376), .A3(new_n384), .A4(new_n377), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n326), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(G214), .B1(G237), .B2(G902), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT6), .ZN(new_n391));
  INV_X1    g205(.A(G104), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G107), .ZN(new_n393));
  INV_X1    g207(.A(G107), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G104), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G101), .ZN(new_n397));
  OAI21_X1  g211(.A(KEYINPUT3), .B1(new_n392), .B2(G107), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT3), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(new_n394), .A3(G104), .ZN(new_n400));
  INV_X1    g214(.A(G101), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n398), .A2(new_n400), .A3(new_n401), .A4(new_n393), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n402), .A2(KEYINPUT81), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n402), .A2(KEYINPUT81), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n397), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT5), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(new_n242), .A3(G116), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n407), .B1(new_n244), .B2(new_n406), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n256), .B1(new_n408), .B2(new_n251), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n398), .A2(new_n400), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT81), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n411), .A2(new_n412), .A3(new_n401), .A4(new_n393), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n402), .A2(KEYINPUT81), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n398), .A2(new_n400), .A3(new_n393), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G101), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n413), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT4), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT82), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n418), .B1(new_n416), .B2(new_n419), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n415), .A2(KEYINPUT82), .A3(KEYINPUT4), .A4(G101), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n417), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n410), .B1(new_n263), .B2(new_n422), .ZN(new_n423));
  XOR2_X1   g237(.A(G110), .B(G122), .Z(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n391), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NOR3_X1   g240(.A1(new_n250), .A2(new_n257), .A3(new_n246), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n261), .B1(new_n260), .B2(new_n249), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n422), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n410), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n424), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n426), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n230), .A2(G125), .A3(new_n233), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n215), .A2(new_n343), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G224), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n437), .A2(G953), .ZN(new_n438));
  XOR2_X1   g252(.A(new_n436), .B(new_n438), .Z(new_n439));
  INV_X1    g253(.A(KEYINPUT85), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n425), .B1(new_n429), .B2(new_n430), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n440), .B1(new_n441), .B2(new_n391), .ZN(new_n442));
  NOR4_X1   g256(.A1(new_n423), .A2(KEYINPUT85), .A3(KEYINPUT6), .A4(new_n425), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n433), .B(new_n439), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n424), .B(KEYINPUT8), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n405), .A2(new_n409), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n445), .B1(new_n430), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n447), .B1(new_n423), .B2(new_n425), .ZN(new_n448));
  INV_X1    g262(.A(new_n436), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n438), .B(KEYINPUT87), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n438), .B1(KEYINPUT86), .B2(KEYINPUT7), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n452), .B1(KEYINPUT86), .B2(KEYINPUT7), .ZN(new_n453));
  AOI22_X1  g267(.A1(new_n451), .A2(KEYINPUT7), .B1(new_n449), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(G902), .B1(new_n448), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n444), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(G210), .B1(G237), .B2(G902), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n444), .A2(new_n457), .A3(new_n455), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n390), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(G234), .A2(G237), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(G952), .A3(new_n281), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  XOR2_X1   g278(.A(KEYINPUT21), .B(G898), .Z(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n462), .A2(G902), .A3(G953), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n464), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n461), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(G478), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n472), .A2(KEYINPUT15), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT93), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n189), .A2(G128), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n187), .A2(G143), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT92), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(KEYINPUT92), .B1(new_n187), .B2(G143), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n475), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n478), .A2(new_n479), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n480), .B(G134), .C1(new_n481), .C2(KEYINPUT13), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n476), .B(new_n477), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT13), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n483), .B(new_n475), .C1(new_n484), .C2(new_n198), .ZN(new_n485));
  XNOR2_X1  g299(.A(G116), .B(G122), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(new_n394), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n482), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n483), .A2(G134), .A3(new_n475), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n480), .A2(new_n198), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n239), .A2(KEYINPUT14), .A3(G122), .ZN(new_n491));
  INV_X1    g305(.A(new_n486), .ZN(new_n492));
  OAI211_X1 g306(.A(G107), .B(new_n491), .C1(new_n492), .C2(KEYINPUT14), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n486), .A2(new_n394), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n489), .A2(new_n490), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n488), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(KEYINPUT9), .B(G234), .ZN(new_n497));
  NOR3_X1   g311(.A1(new_n497), .A2(new_n372), .A3(G953), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n488), .A2(new_n495), .A3(new_n498), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n474), .B1(new_n502), .B2(new_n301), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n488), .A2(new_n495), .A3(new_n498), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n498), .B1(new_n488), .B2(new_n495), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n474), .B(new_n301), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n473), .B1(new_n503), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n508), .B1(new_n473), .B2(new_n503), .ZN(new_n509));
  XNOR2_X1  g323(.A(G113), .B(G122), .ZN(new_n510));
  XNOR2_X1  g324(.A(KEYINPUT89), .B(G104), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n510), .B(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n280), .A2(new_n281), .A3(G214), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n189), .A2(KEYINPUT88), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n514), .B(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n207), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT17), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n514), .A2(KEYINPUT88), .A3(new_n189), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n515), .A2(G214), .A3(new_n280), .A4(new_n281), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(G131), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n517), .A2(new_n518), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n207), .B1(new_n519), .B2(new_n520), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT17), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n523), .A2(new_n357), .A3(new_n347), .A4(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT18), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n516), .B1(new_n527), .B2(new_n207), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n345), .B(new_n191), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n528), .B(new_n529), .C1(new_n527), .C2(new_n522), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n513), .B1(new_n526), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT91), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n526), .A2(new_n513), .A3(new_n530), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT91), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n532), .B(new_n301), .C1(new_n535), .C2(new_n531), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(G475), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT19), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n345), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n354), .A2(KEYINPUT19), .A3(new_n355), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n539), .A2(new_n191), .A3(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n521), .A2(G131), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n347), .B(new_n541), .C1(new_n542), .C2(new_n524), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n530), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n512), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n533), .ZN(new_n546));
  NOR2_X1   g360(.A1(G475), .A2(G902), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT20), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n546), .A2(KEYINPUT90), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT90), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n545), .A2(new_n533), .A3(new_n552), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n551), .A2(KEYINPUT20), .A3(new_n547), .A4(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n537), .A2(new_n550), .A3(new_n554), .ZN(new_n555));
  NOR3_X1   g369(.A1(new_n471), .A2(new_n509), .A3(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(G221), .B1(new_n497), .B2(G902), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n397), .B(new_n215), .C1(new_n403), .C2(new_n404), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n413), .A2(new_n414), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n215), .B1(new_n561), .B2(new_n397), .ZN(new_n562));
  OAI211_X1 g376(.A(KEYINPUT12), .B(new_n219), .C1(new_n560), .C2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT83), .ZN(new_n564));
  INV_X1    g378(.A(new_n219), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n405), .A2(new_n197), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n565), .B1(new_n566), .B2(new_n559), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT83), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n567), .A2(new_n568), .A3(KEYINPUT12), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n219), .B1(new_n560), .B2(new_n562), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT12), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n564), .A2(new_n569), .A3(new_n572), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n413), .A2(new_n414), .B1(G101), .B2(new_n396), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT10), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n575), .B1(new_n271), .B2(new_n273), .ZN(new_n576));
  AOI22_X1  g390(.A1(new_n574), .A2(new_n576), .B1(new_n559), .B2(new_n575), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n422), .A2(new_n266), .A3(new_n268), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(new_n578), .A3(new_n565), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n573), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n281), .A2(G227), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(G140), .ZN(new_n582));
  XNOR2_X1  g396(.A(KEYINPUT80), .B(G110), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n582), .B(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n577), .A2(new_n578), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT84), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n577), .A2(new_n578), .A3(KEYINPUT84), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n587), .A2(new_n219), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n584), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n579), .A2(new_n590), .ZN(new_n591));
  AOI22_X1  g405(.A1(new_n580), .A2(new_n584), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(G469), .B1(new_n592), .B2(G902), .ZN(new_n593));
  INV_X1    g407(.A(G469), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n590), .B1(new_n589), .B2(new_n579), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n573), .A2(new_n591), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n594), .B(new_n301), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n558), .B1(new_n593), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n388), .A2(new_n556), .A3(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(G101), .ZN(G3));
  INV_X1    g414(.A(new_n387), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n593), .A2(new_n597), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n557), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n324), .A2(new_n301), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(G472), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n310), .B1(new_n319), .B2(new_n320), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n601), .A2(new_n603), .A3(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n472), .A2(new_n301), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n502), .A2(new_n472), .A3(new_n301), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(KEYINPUT33), .B1(new_n498), .B2(KEYINPUT94), .ZN(new_n612));
  OR2_X1    g426(.A1(new_n502), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n502), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI211_X1 g429(.A(new_n609), .B(new_n611), .C1(new_n615), .C2(G478), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n555), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n471), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n608), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G104), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT95), .B(KEYINPUT34), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G6));
  AND3_X1   g436(.A1(new_n444), .A2(new_n457), .A3(new_n455), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n457), .B1(new_n444), .B2(new_n455), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n389), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n509), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n537), .A2(new_n554), .ZN(new_n627));
  AND2_X1   g441(.A1(new_n551), .A2(new_n553), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n628), .A2(new_n547), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n627), .B1(new_n629), .B2(KEYINPUT20), .ZN(new_n630));
  NOR4_X1   g444(.A1(new_n625), .A2(new_n626), .A3(new_n469), .A4(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n608), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT35), .B(G107), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  NOR2_X1   g448(.A1(new_n607), .A2(new_n603), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT97), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT96), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n350), .A2(new_n360), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n369), .A2(KEYINPUT36), .ZN(new_n639));
  OR2_X1    g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n640), .A2(new_n374), .A3(new_n641), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n383), .A2(new_n637), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n637), .B1(new_n383), .B2(new_n642), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n636), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n383), .A2(new_n642), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(KEYINPUT96), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n383), .A2(new_n637), .A3(new_n642), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n647), .A2(KEYINPUT97), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n645), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n556), .A2(new_n635), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT37), .B(G110), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G12));
  NOR2_X1   g468(.A1(new_n650), .A2(new_n625), .ZN(new_n655));
  OR3_X1    g469(.A1(new_n467), .A2(KEYINPUT98), .A3(G900), .ZN(new_n656));
  OAI21_X1  g470(.A(KEYINPUT98), .B1(new_n467), .B2(G900), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n656), .A2(new_n463), .A3(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n630), .A2(new_n626), .A3(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n655), .A2(new_n326), .A3(new_n598), .A4(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(KEYINPUT99), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n606), .A2(KEYINPUT32), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n321), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n603), .B1(new_n664), .B2(new_n308), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT99), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n665), .A2(new_n666), .A3(new_n660), .A4(new_n655), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n662), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G128), .ZN(G30));
  XOR2_X1   g483(.A(new_n658), .B(KEYINPUT39), .Z(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n598), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(KEYINPUT40), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n459), .A2(new_n460), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(new_n676));
  OR2_X1    g490(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n643), .A2(new_n644), .ZN(new_n678));
  AOI211_X1 g492(.A(new_n390), .B(new_n678), .C1(new_n672), .C2(KEYINPUT40), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n286), .B1(new_n302), .B2(new_n303), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n315), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g495(.A(G472), .B1(new_n681), .B2(G902), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n682), .B1(new_n322), .B2(new_n325), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n555), .ZN(new_n685));
  NOR4_X1   g499(.A1(new_n677), .A2(new_n684), .A3(new_n626), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT101), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(new_n189), .ZN(G45));
  NAND3_X1  g502(.A1(new_n616), .A2(new_n555), .A3(new_n658), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n655), .A2(new_n326), .A3(new_n598), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G146), .ZN(G48));
  OAI21_X1  g506(.A(new_n301), .B1(new_n595), .B2(new_n596), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(G469), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(new_n557), .A3(new_n597), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n618), .A2(new_n696), .A3(new_n387), .A4(new_n326), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT41), .B(G113), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G15));
  NAND4_X1  g513(.A1(new_n631), .A2(new_n696), .A3(new_n387), .A4(new_n326), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G116), .ZN(G18));
  NOR2_X1   g515(.A1(new_n695), .A2(new_n625), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n556), .A2(new_n326), .A3(new_n651), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G119), .ZN(G21));
  INV_X1    g518(.A(KEYINPUT103), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n294), .A2(KEYINPUT102), .A3(new_n304), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT102), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n285), .B1(new_n305), .B2(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n319), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n310), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n705), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n706), .ZN(new_n712));
  AOI21_X1  g526(.A(KEYINPUT102), .B1(new_n294), .B2(new_n304), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n712), .A2(new_n713), .A3(new_n285), .ZN(new_n714));
  OAI211_X1 g528(.A(KEYINPUT103), .B(new_n310), .C1(new_n714), .C2(new_n319), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n711), .A2(new_n605), .A3(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n378), .A2(new_n384), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n555), .A2(new_n509), .A3(KEYINPUT104), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n718), .B(new_n389), .C1(new_n623), .C2(new_n624), .ZN(new_n719));
  AOI21_X1  g533(.A(KEYINPUT104), .B1(new_n555), .B2(new_n509), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n719), .A2(new_n469), .A3(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n716), .A2(new_n717), .A3(new_n696), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G122), .ZN(G24));
  INV_X1    g537(.A(KEYINPUT105), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n695), .A2(new_n625), .A3(new_n689), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n716), .A2(new_n724), .A3(new_n678), .A4(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n711), .A2(new_n605), .A3(new_n715), .A4(new_n678), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n694), .A2(new_n597), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n728), .A2(new_n461), .A3(new_n557), .A4(new_n690), .ZN(new_n729));
  OAI21_X1  g543(.A(KEYINPUT105), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(KEYINPUT106), .B(G125), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n731), .B(new_n732), .ZN(G27));
  NOR2_X1   g547(.A1(new_n623), .A2(new_n624), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n690), .A2(new_n389), .A3(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n603), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n388), .A2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT42), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n664), .A2(KEYINPUT107), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT107), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n663), .A2(new_n741), .A3(new_n321), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n740), .A2(new_n308), .A3(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n743), .A2(KEYINPUT42), .A3(new_n717), .A4(new_n736), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n739), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G131), .ZN(G33));
  NAND4_X1  g560(.A1(new_n326), .A2(new_n387), .A3(new_n598), .A4(new_n660), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT108), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n734), .A2(new_n389), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n748), .B1(new_n747), .B2(new_n749), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n198), .ZN(G36));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n592), .B(new_n755), .ZN(new_n756));
  OAI21_X1  g570(.A(G469), .B1(new_n756), .B2(G902), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(KEYINPUT46), .ZN(new_n758));
  OR2_X1    g572(.A1(new_n758), .A2(KEYINPUT109), .ZN(new_n759));
  OR2_X1    g573(.A1(new_n757), .A2(KEYINPUT46), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n758), .A2(KEYINPUT109), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n759), .A2(new_n597), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n557), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n763), .A2(new_n670), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n685), .A2(new_n616), .ZN(new_n765));
  XOR2_X1   g579(.A(new_n765), .B(KEYINPUT43), .Z(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n607), .A3(new_n678), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(KEYINPUT44), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n749), .B(KEYINPUT110), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n764), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G137), .ZN(G39));
  NOR2_X1   g585(.A1(new_n326), .A2(new_n735), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n762), .A2(KEYINPUT47), .A3(new_n557), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT47), .B1(new_n762), .B2(new_n557), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n601), .B(new_n772), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G140), .ZN(G42));
  NOR2_X1   g590(.A1(new_n749), .A2(new_n695), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n766), .A2(new_n464), .A3(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n778), .A2(new_n717), .A3(new_n743), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT48), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n281), .A2(G952), .ZN(new_n782));
  AND4_X1   g596(.A1(new_n464), .A2(new_n716), .A3(new_n717), .A4(new_n766), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n782), .B1(new_n783), .B2(new_n702), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n786));
  INV_X1    g600(.A(new_n777), .ZN(new_n787));
  NOR4_X1   g601(.A1(new_n787), .A2(new_n601), .A3(new_n463), .A4(new_n683), .ZN(new_n788));
  INV_X1    g602(.A(new_n616), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n788), .A2(new_n685), .A3(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT117), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n727), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n778), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n790), .A2(new_n791), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n792), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n786), .B1(new_n796), .B2(KEYINPUT118), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n797), .B1(KEYINPUT118), .B2(new_n796), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n773), .A2(new_n774), .ZN(new_n799));
  INV_X1    g613(.A(new_n728), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n799), .B1(new_n557), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n801), .A2(new_n769), .A3(new_n783), .ZN(new_n802));
  NOR2_X1   g616(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n695), .A2(new_n389), .A3(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n783), .A2(new_n676), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n802), .A2(new_n807), .ZN(new_n808));
  OAI221_X1 g622(.A(new_n785), .B1(new_n780), .B2(new_n779), .C1(new_n798), .C2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n796), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n802), .A2(new_n807), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n809), .B1(new_n786), .B2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n788), .A2(new_n555), .A3(new_n616), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n814));
  AOI22_X1  g628(.A1(new_n751), .A2(new_n752), .B1(new_n739), .B2(new_n744), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n599), .A2(new_n652), .A3(new_n697), .A4(new_n700), .ZN(new_n816));
  INV_X1    g630(.A(new_n471), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n617), .B1(new_n626), .B2(new_n555), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n635), .A2(new_n817), .A3(new_n387), .A4(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n703), .A2(new_n722), .A3(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n749), .A2(new_n509), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n650), .A2(new_n630), .A3(new_n659), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n665), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  XOR2_X1   g638(.A(new_n824), .B(KEYINPUT112), .Z(new_n825));
  NAND2_X1  g639(.A1(new_n793), .A2(new_n736), .ZN(new_n826));
  AND4_X1   g640(.A1(new_n815), .A2(new_n821), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  AOI22_X1  g641(.A1(new_n667), .A2(new_n662), .B1(new_n726), .B2(new_n730), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(KEYINPUT113), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n719), .A2(new_n720), .ZN(new_n830));
  INV_X1    g644(.A(new_n646), .ZN(new_n831));
  AOI211_X1 g645(.A(new_n558), .B(new_n659), .C1(new_n593), .C2(new_n597), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n830), .A2(new_n683), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n691), .A2(new_n833), .A3(KEYINPUT52), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n829), .A2(new_n835), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n691), .A2(new_n833), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT52), .B1(new_n828), .B2(new_n837), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n814), .B(new_n827), .C1(new_n836), .C2(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n815), .A2(new_n821), .A3(new_n825), .A4(new_n826), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n668), .A2(new_n834), .A3(new_n731), .ZN(new_n841));
  OAI21_X1  g655(.A(KEYINPUT114), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n668), .A2(new_n731), .A3(new_n837), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT52), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT114), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n828), .A2(new_n834), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n840), .B1(new_n842), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n839), .B1(new_n814), .B2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n851));
  OR2_X1    g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT115), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n853), .B1(new_n849), .B2(KEYINPUT53), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n838), .A2(KEYINPUT114), .A3(new_n841), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n846), .B1(new_n845), .B2(new_n847), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n827), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n857), .A2(KEYINPUT115), .A3(new_n814), .ZN(new_n858));
  OAI211_X1 g672(.A(KEYINPUT53), .B(new_n827), .C1(new_n836), .C2(new_n838), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n854), .A2(new_n858), .A3(new_n851), .A4(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n812), .A2(new_n813), .A3(new_n852), .A4(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n861), .B1(G952), .B2(G953), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n717), .A2(new_n389), .A3(new_n557), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n863), .A2(KEYINPUT111), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(new_n765), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n683), .B1(KEYINPUT111), .B2(new_n863), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n728), .B(KEYINPUT49), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n865), .A2(new_n676), .A3(new_n866), .A4(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n862), .A2(new_n868), .ZN(G75));
  NAND3_X1  g683(.A1(new_n854), .A2(new_n858), .A3(new_n859), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n870), .A2(G210), .A3(G902), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT56), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n871), .A2(KEYINPUT119), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n433), .B1(new_n442), .B2(new_n443), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(new_n439), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n875), .B(KEYINPUT55), .Z(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  OR2_X1    g691(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n281), .A2(G952), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT119), .B1(new_n871), .B2(new_n872), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n877), .B1(new_n873), .B2(new_n881), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n878), .A2(new_n880), .A3(new_n882), .ZN(G51));
  NAND2_X1  g697(.A1(new_n870), .A2(KEYINPUT54), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n860), .ZN(new_n885));
  NAND2_X1  g699(.A1(G469), .A2(G902), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n886), .B(KEYINPUT57), .Z(new_n887));
  NAND2_X1  g701(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n595), .A2(new_n596), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n888), .A2(KEYINPUT120), .A3(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n870), .A2(G469), .A3(G902), .A4(new_n756), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT120), .ZN(new_n893));
  INV_X1    g707(.A(new_n887), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n894), .B1(new_n884), .B2(new_n860), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n893), .B1(new_n895), .B2(new_n889), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n891), .A2(new_n892), .A3(new_n896), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n897), .A2(new_n880), .ZN(G54));
  NAND4_X1  g712(.A1(new_n870), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n899));
  INV_X1    g713(.A(new_n628), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT121), .ZN(new_n902));
  OR3_X1    g716(.A1(new_n899), .A2(new_n902), .A3(new_n900), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n902), .B1(new_n899), .B2(new_n900), .ZN(new_n904));
  AOI211_X1 g718(.A(new_n879), .B(new_n901), .C1(new_n903), .C2(new_n904), .ZN(G60));
  XNOR2_X1  g719(.A(new_n609), .B(KEYINPUT59), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n906), .B1(new_n852), .B2(new_n860), .ZN(new_n907));
  INV_X1    g721(.A(new_n615), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n880), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n906), .B1(new_n884), .B2(new_n860), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n909), .B1(new_n908), .B2(new_n910), .ZN(G63));
  XNOR2_X1  g725(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n372), .A2(new_n301), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n912), .B(new_n913), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n870), .A2(new_n641), .A3(new_n640), .A4(new_n914), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n870), .A2(new_n914), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n880), .B(new_n915), .C1(new_n916), .C2(new_n371), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g732(.A(G953), .B1(new_n466), .B2(new_n437), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n919), .B1(new_n821), .B2(G953), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n874), .B1(G898), .B2(new_n281), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n920), .B(new_n921), .ZN(G69));
  NAND2_X1  g736(.A1(new_n775), .A2(new_n770), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n818), .A2(new_n598), .A3(new_n671), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n388), .A2(new_n389), .A3(new_n734), .A4(new_n925), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT123), .Z(new_n927));
  INV_X1    g741(.A(new_n691), .ZN(new_n928));
  OR2_X1    g742(.A1(new_n829), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n929), .A2(new_n687), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n930), .A2(KEYINPUT62), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n930), .A2(KEYINPUT62), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n924), .B(new_n927), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n237), .B1(new_n276), .B2(new_n236), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n539), .A2(new_n540), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n934), .B(new_n935), .Z(new_n936));
  NAND3_X1  g750(.A1(new_n933), .A2(new_n281), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n281), .B1(G227), .B2(G900), .ZN(new_n938));
  XOR2_X1   g752(.A(KEYINPUT124), .B(G900), .Z(new_n939));
  OAI21_X1  g753(.A(new_n938), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT125), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n936), .A2(new_n938), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n764), .A2(new_n717), .A3(new_n830), .A4(new_n743), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n815), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n929), .A2(new_n944), .A3(new_n923), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n942), .B1(new_n945), .B2(G953), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n937), .A2(new_n941), .A3(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT126), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n947), .B(new_n948), .ZN(G72));
  INV_X1    g763(.A(new_n279), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n945), .A2(new_n821), .ZN(new_n951));
  NAND2_X1  g765(.A1(G472), .A2(G902), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT63), .Z(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n286), .B(new_n950), .C1(new_n951), .C2(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n315), .B1(new_n950), .B2(new_n285), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n953), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT127), .Z(new_n958));
  OAI211_X1 g772(.A(new_n955), .B(new_n880), .C1(new_n850), .C2(new_n958), .ZN(new_n959));
  OR3_X1    g773(.A1(new_n933), .A2(new_n820), .A3(new_n816), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n950), .B1(new_n960), .B2(new_n953), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n959), .B1(new_n961), .B2(new_n285), .ZN(G57));
endmodule


