

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U555 ( .A(KEYINPUT32), .B(n676), .ZN(n684) );
  AND2_X2 U556 ( .A1(n675), .A2(n674), .ZN(n676) );
  OR2_X1 U557 ( .A1(n761), .A2(n760), .ZN(n762) );
  NOR2_X2 U558 ( .A1(G2105), .A2(n527), .ZN(n889) );
  NOR2_X1 U559 ( .A1(n532), .A2(n531), .ZN(G160) );
  OR2_X1 U560 ( .A1(n754), .A2(n690), .ZN(n521) );
  NAND2_X1 U561 ( .A1(n688), .A2(n754), .ZN(n522) );
  INV_X1 U562 ( .A(KEYINPUT69), .ZN(n606) );
  XNOR2_X1 U563 ( .A(n606), .B(KEYINPUT14), .ZN(n607) );
  XNOR2_X1 U564 ( .A(n608), .B(n607), .ZN(n610) );
  XOR2_X1 U565 ( .A(KEYINPUT1), .B(n541), .Z(n796) );
  NOR2_X1 U566 ( .A1(G2105), .A2(G2104), .ZN(n523) );
  XOR2_X2 U567 ( .A(KEYINPUT17), .B(n523), .Z(n888) );
  NAND2_X1 U568 ( .A1(n888), .A2(G137), .ZN(n526) );
  INV_X1 U569 ( .A(G2104), .ZN(n527) );
  NAND2_X1 U570 ( .A1(G101), .A2(n889), .ZN(n524) );
  XOR2_X1 U571 ( .A(KEYINPUT23), .B(n524), .Z(n525) );
  NAND2_X1 U572 ( .A1(n526), .A2(n525), .ZN(n532) );
  INV_X1 U573 ( .A(G2105), .ZN(n528) );
  NOR2_X1 U574 ( .A1(n528), .A2(n527), .ZN(n883) );
  NAND2_X1 U575 ( .A1(G113), .A2(n883), .ZN(n530) );
  NOR2_X1 U576 ( .A1(G2104), .A2(n528), .ZN(n884) );
  NAND2_X1 U577 ( .A1(G125), .A2(n884), .ZN(n529) );
  NAND2_X1 U578 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U579 ( .A1(G138), .A2(n888), .ZN(n534) );
  NAND2_X1 U580 ( .A1(G102), .A2(n889), .ZN(n533) );
  NAND2_X1 U581 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U582 ( .A(n535), .B(KEYINPUT93), .ZN(n537) );
  NAND2_X1 U583 ( .A1(G126), .A2(n884), .ZN(n536) );
  NAND2_X1 U584 ( .A1(n537), .A2(n536), .ZN(n540) );
  NAND2_X1 U585 ( .A1(G114), .A2(n883), .ZN(n538) );
  XOR2_X1 U586 ( .A(KEYINPUT92), .B(n538), .Z(n539) );
  NOR2_X2 U587 ( .A1(n540), .A2(n539), .ZN(G164) );
  XOR2_X1 U588 ( .A(G543), .B(KEYINPUT0), .Z(n599) );
  NOR2_X1 U589 ( .A1(G651), .A2(n599), .ZN(n795) );
  NAND2_X1 U590 ( .A1(n795), .A2(G52), .ZN(n543) );
  XNOR2_X1 U591 ( .A(KEYINPUT65), .B(G651), .ZN(n544) );
  NOR2_X1 U592 ( .A1(G543), .A2(n544), .ZN(n541) );
  NAND2_X1 U593 ( .A1(G64), .A2(n796), .ZN(n542) );
  NAND2_X1 U594 ( .A1(n543), .A2(n542), .ZN(n549) );
  NOR2_X1 U595 ( .A1(G651), .A2(G543), .ZN(n800) );
  NAND2_X1 U596 ( .A1(n800), .A2(G90), .ZN(n546) );
  NOR2_X1 U597 ( .A1(n599), .A2(n544), .ZN(n803) );
  NAND2_X1 U598 ( .A1(G77), .A2(n803), .ZN(n545) );
  NAND2_X1 U599 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U600 ( .A(KEYINPUT9), .B(n547), .Z(n548) );
  NOR2_X1 U601 ( .A1(n549), .A2(n548), .ZN(G171) );
  NAND2_X1 U602 ( .A1(n796), .A2(G65), .ZN(n550) );
  XNOR2_X1 U603 ( .A(n550), .B(KEYINPUT68), .ZN(n557) );
  NAND2_X1 U604 ( .A1(G91), .A2(n800), .ZN(n552) );
  NAND2_X1 U605 ( .A1(G53), .A2(n795), .ZN(n551) );
  NAND2_X1 U606 ( .A1(n552), .A2(n551), .ZN(n555) );
  NAND2_X1 U607 ( .A1(G78), .A2(n803), .ZN(n553) );
  XNOR2_X1 U608 ( .A(KEYINPUT67), .B(n553), .ZN(n554) );
  NOR2_X1 U609 ( .A1(n555), .A2(n554), .ZN(n556) );
  NAND2_X1 U610 ( .A1(n557), .A2(n556), .ZN(G299) );
  NAND2_X1 U611 ( .A1(n795), .A2(G51), .ZN(n559) );
  NAND2_X1 U612 ( .A1(G63), .A2(n796), .ZN(n558) );
  NAND2_X1 U613 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U614 ( .A(KEYINPUT6), .B(n560), .ZN(n566) );
  NAND2_X1 U615 ( .A1(n800), .A2(G89), .ZN(n561) );
  XNOR2_X1 U616 ( .A(n561), .B(KEYINPUT4), .ZN(n563) );
  NAND2_X1 U617 ( .A1(G76), .A2(n803), .ZN(n562) );
  NAND2_X1 U618 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U619 ( .A(n564), .B(KEYINPUT5), .Z(n565) );
  NOR2_X1 U620 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U621 ( .A(KEYINPUT77), .B(n567), .Z(n569) );
  XOR2_X1 U622 ( .A(KEYINPUT76), .B(KEYINPUT7), .Z(n568) );
  XNOR2_X1 U623 ( .A(n569), .B(n568), .ZN(G168) );
  XOR2_X1 U624 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U625 ( .A1(n803), .A2(G75), .ZN(n570) );
  XNOR2_X1 U626 ( .A(n570), .B(KEYINPUT86), .ZN(n577) );
  NAND2_X1 U627 ( .A1(G88), .A2(n800), .ZN(n572) );
  NAND2_X1 U628 ( .A1(G50), .A2(n795), .ZN(n571) );
  NAND2_X1 U629 ( .A1(n572), .A2(n571), .ZN(n575) );
  NAND2_X1 U630 ( .A1(G62), .A2(n796), .ZN(n573) );
  XNOR2_X1 U631 ( .A(KEYINPUT85), .B(n573), .ZN(n574) );
  NOR2_X1 U632 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U633 ( .A1(n577), .A2(n576), .ZN(G303) );
  NAND2_X1 U634 ( .A1(G73), .A2(n803), .ZN(n579) );
  XNOR2_X1 U635 ( .A(KEYINPUT2), .B(KEYINPUT84), .ZN(n578) );
  XNOR2_X1 U636 ( .A(n579), .B(n578), .ZN(n586) );
  NAND2_X1 U637 ( .A1(G86), .A2(n800), .ZN(n581) );
  NAND2_X1 U638 ( .A1(G48), .A2(n795), .ZN(n580) );
  NAND2_X1 U639 ( .A1(n581), .A2(n580), .ZN(n584) );
  NAND2_X1 U640 ( .A1(G61), .A2(n796), .ZN(n582) );
  XNOR2_X1 U641 ( .A(KEYINPUT83), .B(n582), .ZN(n583) );
  NOR2_X1 U642 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U643 ( .A1(n586), .A2(n585), .ZN(G305) );
  NAND2_X1 U644 ( .A1(G85), .A2(n800), .ZN(n587) );
  XNOR2_X1 U645 ( .A(n587), .B(KEYINPUT64), .ZN(n594) );
  NAND2_X1 U646 ( .A1(n795), .A2(G47), .ZN(n589) );
  NAND2_X1 U647 ( .A1(G60), .A2(n796), .ZN(n588) );
  NAND2_X1 U648 ( .A1(n589), .A2(n588), .ZN(n592) );
  NAND2_X1 U649 ( .A1(n803), .A2(G72), .ZN(n590) );
  XOR2_X1 U650 ( .A(KEYINPUT66), .B(n590), .Z(n591) );
  NOR2_X1 U651 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U652 ( .A1(n594), .A2(n593), .ZN(G290) );
  NAND2_X1 U653 ( .A1(G49), .A2(n795), .ZN(n596) );
  NAND2_X1 U654 ( .A1(G74), .A2(G651), .ZN(n595) );
  NAND2_X1 U655 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U656 ( .A(KEYINPUT82), .B(n597), .ZN(n598) );
  NOR2_X1 U657 ( .A1(n796), .A2(n598), .ZN(n601) );
  NAND2_X1 U658 ( .A1(n599), .A2(G87), .ZN(n600) );
  NAND2_X1 U659 ( .A1(n601), .A2(n600), .ZN(G288) );
  NOR2_X2 U660 ( .A1(G164), .A2(G1384), .ZN(n702) );
  NAND2_X1 U661 ( .A1(G160), .A2(G40), .ZN(n703) );
  INV_X1 U662 ( .A(n703), .ZN(n602) );
  NAND2_X1 U663 ( .A1(n702), .A2(n602), .ZN(n668) );
  NAND2_X1 U664 ( .A1(n668), .A2(G1961), .ZN(n604) );
  AND2_X2 U665 ( .A1(n702), .A2(n602), .ZN(n645) );
  XOR2_X1 U666 ( .A(G2078), .B(KEYINPUT25), .Z(n923) );
  NAND2_X1 U667 ( .A1(n645), .A2(n923), .ZN(n603) );
  NAND2_X1 U668 ( .A1(n604), .A2(n603), .ZN(n605) );
  XOR2_X1 U669 ( .A(n605), .B(KEYINPUT100), .Z(n662) );
  NAND2_X1 U670 ( .A1(n662), .A2(G171), .ZN(n657) );
  INV_X1 U671 ( .A(KEYINPUT71), .ZN(n619) );
  NAND2_X1 U672 ( .A1(n796), .A2(G56), .ZN(n608) );
  NAND2_X1 U673 ( .A1(G43), .A2(n795), .ZN(n609) );
  NAND2_X1 U674 ( .A1(n610), .A2(n609), .ZN(n617) );
  NAND2_X1 U675 ( .A1(n800), .A2(G81), .ZN(n611) );
  XNOR2_X1 U676 ( .A(n611), .B(KEYINPUT12), .ZN(n613) );
  NAND2_X1 U677 ( .A1(G68), .A2(n803), .ZN(n612) );
  NAND2_X1 U678 ( .A1(n613), .A2(n612), .ZN(n614) );
  XOR2_X1 U679 ( .A(KEYINPUT70), .B(n614), .Z(n615) );
  XNOR2_X1 U680 ( .A(KEYINPUT13), .B(n615), .ZN(n616) );
  NOR2_X1 U681 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X2 U682 ( .A(n619), .B(n618), .ZN(n997) );
  NAND2_X1 U683 ( .A1(G1996), .A2(n645), .ZN(n620) );
  XNOR2_X1 U684 ( .A(n620), .B(KEYINPUT26), .ZN(n622) );
  NAND2_X1 U685 ( .A1(G1341), .A2(n668), .ZN(n621) );
  NAND2_X1 U686 ( .A1(n622), .A2(n621), .ZN(n623) );
  XOR2_X1 U687 ( .A(n623), .B(KEYINPUT102), .Z(n624) );
  NAND2_X1 U688 ( .A1(n997), .A2(n624), .ZN(n640) );
  NAND2_X1 U689 ( .A1(G54), .A2(n795), .ZN(n625) );
  XNOR2_X1 U690 ( .A(n625), .B(KEYINPUT74), .ZN(n630) );
  NAND2_X1 U691 ( .A1(n800), .A2(G92), .ZN(n627) );
  NAND2_X1 U692 ( .A1(G66), .A2(n796), .ZN(n626) );
  NAND2_X1 U693 ( .A1(n627), .A2(n626), .ZN(n628) );
  XOR2_X1 U694 ( .A(KEYINPUT72), .B(n628), .Z(n629) );
  NAND2_X1 U695 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U696 ( .A1(G79), .A2(n803), .ZN(n631) );
  XNOR2_X1 U697 ( .A(KEYINPUT73), .B(n631), .ZN(n632) );
  NOR2_X1 U698 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U699 ( .A(KEYINPUT15), .B(n634), .ZN(n1017) );
  NOR2_X1 U700 ( .A1(n640), .A2(n1017), .ZN(n635) );
  XNOR2_X1 U701 ( .A(n635), .B(KEYINPUT103), .ZN(n639) );
  NOR2_X1 U702 ( .A1(n645), .A2(G1348), .ZN(n637) );
  NOR2_X1 U703 ( .A1(G2067), .A2(n668), .ZN(n636) );
  NOR2_X1 U704 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U705 ( .A1(n639), .A2(n638), .ZN(n642) );
  NAND2_X1 U706 ( .A1(n640), .A2(n1017), .ZN(n641) );
  NAND2_X1 U707 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U708 ( .A(n643), .B(KEYINPUT104), .ZN(n649) );
  NAND2_X1 U709 ( .A1(n645), .A2(G2072), .ZN(n644) );
  XNOR2_X1 U710 ( .A(n644), .B(KEYINPUT27), .ZN(n647) );
  INV_X1 U711 ( .A(G1956), .ZN(n970) );
  NOR2_X1 U712 ( .A1(n970), .A2(n645), .ZN(n646) );
  NOR2_X1 U713 ( .A1(n647), .A2(n646), .ZN(n650) );
  INV_X1 U714 ( .A(G299), .ZN(n1002) );
  NAND2_X1 U715 ( .A1(n650), .A2(n1002), .ZN(n648) );
  NAND2_X1 U716 ( .A1(n649), .A2(n648), .ZN(n654) );
  NOR2_X1 U717 ( .A1(n650), .A2(n1002), .ZN(n652) );
  XNOR2_X1 U718 ( .A(KEYINPUT28), .B(KEYINPUT101), .ZN(n651) );
  XNOR2_X1 U719 ( .A(n652), .B(n651), .ZN(n653) );
  NAND2_X1 U720 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U721 ( .A(KEYINPUT29), .B(n655), .Z(n656) );
  NAND2_X1 U722 ( .A1(n657), .A2(n656), .ZN(n667) );
  NAND2_X1 U723 ( .A1(G8), .A2(n668), .ZN(n754) );
  NOR2_X1 U724 ( .A1(G1966), .A2(n754), .ZN(n680) );
  NOR2_X1 U725 ( .A1(G2084), .A2(n668), .ZN(n677) );
  NOR2_X1 U726 ( .A1(n680), .A2(n677), .ZN(n658) );
  NAND2_X1 U727 ( .A1(G8), .A2(n658), .ZN(n659) );
  XNOR2_X1 U728 ( .A(KEYINPUT30), .B(n659), .ZN(n660) );
  NOR2_X1 U729 ( .A1(G168), .A2(n660), .ZN(n661) );
  XNOR2_X1 U730 ( .A(n661), .B(KEYINPUT105), .ZN(n664) );
  OR2_X1 U731 ( .A1(n662), .A2(G171), .ZN(n663) );
  NAND2_X1 U732 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U733 ( .A(KEYINPUT31), .B(n665), .ZN(n666) );
  NAND2_X1 U734 ( .A1(n667), .A2(n666), .ZN(n678) );
  NAND2_X1 U735 ( .A1(n678), .A2(G286), .ZN(n675) );
  INV_X1 U736 ( .A(G8), .ZN(n673) );
  NOR2_X1 U737 ( .A1(G1971), .A2(n754), .ZN(n670) );
  NOR2_X1 U738 ( .A1(G2090), .A2(n668), .ZN(n669) );
  NOR2_X1 U739 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U740 ( .A1(n671), .A2(G303), .ZN(n672) );
  OR2_X1 U741 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U742 ( .A1(G8), .A2(n677), .ZN(n682) );
  INV_X1 U743 ( .A(n678), .ZN(n679) );
  NOR2_X1 U744 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U745 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U746 ( .A1(n684), .A2(n683), .ZN(n746) );
  NOR2_X1 U747 ( .A1(G2090), .A2(G303), .ZN(n685) );
  XNOR2_X1 U748 ( .A(n685), .B(KEYINPUT110), .ZN(n686) );
  NAND2_X1 U749 ( .A1(n686), .A2(G8), .ZN(n687) );
  NAND2_X1 U750 ( .A1(n746), .A2(n687), .ZN(n688) );
  NOR2_X1 U751 ( .A1(G1981), .A2(G305), .ZN(n689) );
  XOR2_X1 U752 ( .A(n689), .B(KEYINPUT24), .Z(n690) );
  NAND2_X1 U753 ( .A1(n522), .A2(n521), .ZN(n727) );
  NAND2_X1 U754 ( .A1(G140), .A2(n888), .ZN(n692) );
  NAND2_X1 U755 ( .A1(G104), .A2(n889), .ZN(n691) );
  NAND2_X1 U756 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U757 ( .A(KEYINPUT34), .B(n693), .ZN(n699) );
  NAND2_X1 U758 ( .A1(n883), .A2(G116), .ZN(n694) );
  XOR2_X1 U759 ( .A(KEYINPUT95), .B(n694), .Z(n696) );
  NAND2_X1 U760 ( .A1(n884), .A2(G128), .ZN(n695) );
  NAND2_X1 U761 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U762 ( .A(n697), .B(KEYINPUT35), .Z(n698) );
  NOR2_X1 U763 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U764 ( .A(KEYINPUT36), .B(n700), .Z(n701) );
  XOR2_X1 U765 ( .A(KEYINPUT96), .B(n701), .Z(n901) );
  XNOR2_X1 U766 ( .A(G2067), .B(KEYINPUT37), .ZN(n736) );
  NOR2_X1 U767 ( .A1(n901), .A2(n736), .ZN(n950) );
  NOR2_X1 U768 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U769 ( .A(n704), .B(KEYINPUT94), .ZN(n738) );
  NAND2_X1 U770 ( .A1(n950), .A2(n738), .ZN(n734) );
  INV_X1 U771 ( .A(n738), .ZN(n722) );
  NAND2_X1 U772 ( .A1(G117), .A2(n883), .ZN(n706) );
  NAND2_X1 U773 ( .A1(G129), .A2(n884), .ZN(n705) );
  NAND2_X1 U774 ( .A1(n706), .A2(n705), .ZN(n709) );
  NAND2_X1 U775 ( .A1(n889), .A2(G105), .ZN(n707) );
  XOR2_X1 U776 ( .A(KEYINPUT38), .B(n707), .Z(n708) );
  NOR2_X1 U777 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U778 ( .A(n710), .B(KEYINPUT98), .ZN(n712) );
  NAND2_X1 U779 ( .A1(G141), .A2(n888), .ZN(n711) );
  NAND2_X1 U780 ( .A1(n712), .A2(n711), .ZN(n904) );
  NAND2_X1 U781 ( .A1(G1996), .A2(n904), .ZN(n713) );
  XNOR2_X1 U782 ( .A(n713), .B(KEYINPUT99), .ZN(n721) );
  XNOR2_X1 U783 ( .A(KEYINPUT97), .B(G1991), .ZN(n922) );
  NAND2_X1 U784 ( .A1(G131), .A2(n888), .ZN(n715) );
  NAND2_X1 U785 ( .A1(G119), .A2(n884), .ZN(n714) );
  NAND2_X1 U786 ( .A1(n715), .A2(n714), .ZN(n719) );
  NAND2_X1 U787 ( .A1(G95), .A2(n889), .ZN(n717) );
  NAND2_X1 U788 ( .A1(G107), .A2(n883), .ZN(n716) );
  NAND2_X1 U789 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U790 ( .A1(n719), .A2(n718), .ZN(n900) );
  NOR2_X1 U791 ( .A1(n922), .A2(n900), .ZN(n720) );
  NOR2_X1 U792 ( .A1(n721), .A2(n720), .ZN(n952) );
  NOR2_X1 U793 ( .A1(n722), .A2(n952), .ZN(n730) );
  INV_X1 U794 ( .A(n730), .ZN(n723) );
  NAND2_X1 U795 ( .A1(n734), .A2(n723), .ZN(n725) );
  XNOR2_X1 U796 ( .A(G1986), .B(G290), .ZN(n1006) );
  AND2_X1 U797 ( .A1(n1006), .A2(n738), .ZN(n724) );
  OR2_X1 U798 ( .A1(n725), .A2(n724), .ZN(n758) );
  INV_X1 U799 ( .A(n758), .ZN(n726) );
  NAND2_X1 U800 ( .A1(n727), .A2(n726), .ZN(n741) );
  NOR2_X1 U801 ( .A1(G1996), .A2(n904), .ZN(n940) );
  NOR2_X1 U802 ( .A1(G1986), .A2(G290), .ZN(n728) );
  AND2_X1 U803 ( .A1(n922), .A2(n900), .ZN(n943) );
  NOR2_X1 U804 ( .A1(n728), .A2(n943), .ZN(n729) );
  NOR2_X1 U805 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U806 ( .A(KEYINPUT111), .B(n731), .Z(n732) );
  NOR2_X1 U807 ( .A1(n940), .A2(n732), .ZN(n733) );
  XNOR2_X1 U808 ( .A(n733), .B(KEYINPUT39), .ZN(n735) );
  NAND2_X1 U809 ( .A1(n735), .A2(n734), .ZN(n737) );
  NAND2_X1 U810 ( .A1(n901), .A2(n736), .ZN(n954) );
  NAND2_X1 U811 ( .A1(n737), .A2(n954), .ZN(n739) );
  NAND2_X1 U812 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U813 ( .A1(n741), .A2(n740), .ZN(n763) );
  OR2_X1 U814 ( .A1(G1971), .A2(G303), .ZN(n745) );
  NOR2_X1 U815 ( .A1(G1976), .A2(G288), .ZN(n742) );
  XOR2_X1 U816 ( .A(KEYINPUT106), .B(n742), .Z(n1008) );
  INV_X1 U817 ( .A(KEYINPUT33), .ZN(n743) );
  AND2_X1 U818 ( .A1(n1008), .A2(n743), .ZN(n744) );
  AND2_X1 U819 ( .A1(n745), .A2(n744), .ZN(n747) );
  NAND2_X1 U820 ( .A1(n747), .A2(n746), .ZN(n752) );
  INV_X1 U821 ( .A(n754), .ZN(n749) );
  NAND2_X1 U822 ( .A1(G288), .A2(G1976), .ZN(n748) );
  XOR2_X1 U823 ( .A(KEYINPUT107), .B(n748), .Z(n1003) );
  AND2_X1 U824 ( .A1(n749), .A2(n1003), .ZN(n750) );
  OR2_X1 U825 ( .A1(KEYINPUT33), .A2(n750), .ZN(n751) );
  NAND2_X1 U826 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U827 ( .A(n753), .B(KEYINPUT108), .ZN(n761) );
  XOR2_X1 U828 ( .A(G1981), .B(G305), .Z(n1009) );
  NOR2_X1 U829 ( .A1(n754), .A2(n1008), .ZN(n755) );
  NAND2_X1 U830 ( .A1(KEYINPUT33), .A2(n755), .ZN(n756) );
  XOR2_X1 U831 ( .A(KEYINPUT109), .B(n756), .Z(n757) );
  NAND2_X1 U832 ( .A1(n1009), .A2(n757), .ZN(n759) );
  OR2_X1 U833 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U834 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U835 ( .A(n764), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U836 ( .A(G2443), .B(G2446), .Z(n766) );
  XNOR2_X1 U837 ( .A(G2427), .B(G2451), .ZN(n765) );
  XNOR2_X1 U838 ( .A(n766), .B(n765), .ZN(n772) );
  XOR2_X1 U839 ( .A(G2430), .B(G2454), .Z(n768) );
  XNOR2_X1 U840 ( .A(G1341), .B(G1348), .ZN(n767) );
  XNOR2_X1 U841 ( .A(n768), .B(n767), .ZN(n770) );
  XOR2_X1 U842 ( .A(G2435), .B(G2438), .Z(n769) );
  XNOR2_X1 U843 ( .A(n770), .B(n769), .ZN(n771) );
  XOR2_X1 U844 ( .A(n772), .B(n771), .Z(n773) );
  AND2_X1 U845 ( .A1(G14), .A2(n773), .ZN(G401) );
  AND2_X1 U846 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U847 ( .A(G132), .ZN(G219) );
  INV_X1 U848 ( .A(G82), .ZN(G220) );
  INV_X1 U849 ( .A(G120), .ZN(G236) );
  INV_X1 U850 ( .A(G69), .ZN(G235) );
  INV_X1 U851 ( .A(G57), .ZN(G237) );
  NAND2_X1 U852 ( .A1(G7), .A2(G661), .ZN(n774) );
  XNOR2_X1 U853 ( .A(n774), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U854 ( .A(G223), .ZN(n840) );
  NAND2_X1 U855 ( .A1(n840), .A2(G567), .ZN(n775) );
  XOR2_X1 U856 ( .A(KEYINPUT11), .B(n775), .Z(G234) );
  NAND2_X1 U857 ( .A1(n997), .A2(G860), .ZN(G153) );
  INV_X1 U858 ( .A(G171), .ZN(G301) );
  INV_X1 U859 ( .A(n1017), .ZN(n807) );
  NOR2_X1 U860 ( .A1(n807), .A2(G868), .ZN(n776) );
  XNOR2_X1 U861 ( .A(n776), .B(KEYINPUT75), .ZN(n778) );
  NAND2_X1 U862 ( .A1(G868), .A2(G301), .ZN(n777) );
  NAND2_X1 U863 ( .A1(n778), .A2(n777), .ZN(G284) );
  NAND2_X1 U864 ( .A1(G868), .A2(G286), .ZN(n780) );
  INV_X1 U865 ( .A(G868), .ZN(n820) );
  NAND2_X1 U866 ( .A1(G299), .A2(n820), .ZN(n779) );
  NAND2_X1 U867 ( .A1(n780), .A2(n779), .ZN(G297) );
  INV_X1 U868 ( .A(G860), .ZN(n809) );
  NAND2_X1 U869 ( .A1(n809), .A2(G559), .ZN(n781) );
  NAND2_X1 U870 ( .A1(n781), .A2(n807), .ZN(n782) );
  XNOR2_X1 U871 ( .A(n782), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U872 ( .A1(G559), .A2(n1017), .ZN(n783) );
  NOR2_X1 U873 ( .A1(n820), .A2(n783), .ZN(n785) );
  NOR2_X1 U874 ( .A1(n997), .A2(G868), .ZN(n784) );
  OR2_X1 U875 ( .A1(n785), .A2(n784), .ZN(G282) );
  NAND2_X1 U876 ( .A1(G123), .A2(n884), .ZN(n786) );
  XNOR2_X1 U877 ( .A(n786), .B(KEYINPUT18), .ZN(n788) );
  NAND2_X1 U878 ( .A1(n889), .A2(G99), .ZN(n787) );
  NAND2_X1 U879 ( .A1(n788), .A2(n787), .ZN(n792) );
  NAND2_X1 U880 ( .A1(G135), .A2(n888), .ZN(n790) );
  NAND2_X1 U881 ( .A1(G111), .A2(n883), .ZN(n789) );
  NAND2_X1 U882 ( .A1(n790), .A2(n789), .ZN(n791) );
  NOR2_X1 U883 ( .A1(n792), .A2(n791), .ZN(n942) );
  XOR2_X1 U884 ( .A(n942), .B(G2096), .Z(n793) );
  NOR2_X1 U885 ( .A1(G2100), .A2(n793), .ZN(n794) );
  XOR2_X1 U886 ( .A(KEYINPUT78), .B(n794), .Z(G156) );
  NAND2_X1 U887 ( .A1(n795), .A2(G55), .ZN(n798) );
  NAND2_X1 U888 ( .A1(G67), .A2(n796), .ZN(n797) );
  NAND2_X1 U889 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U890 ( .A(n799), .B(KEYINPUT81), .ZN(n802) );
  NAND2_X1 U891 ( .A1(G93), .A2(n800), .ZN(n801) );
  NAND2_X1 U892 ( .A1(n802), .A2(n801), .ZN(n806) );
  NAND2_X1 U893 ( .A1(n803), .A2(G80), .ZN(n804) );
  XOR2_X1 U894 ( .A(KEYINPUT80), .B(n804), .Z(n805) );
  OR2_X1 U895 ( .A1(n806), .A2(n805), .ZN(n819) );
  NAND2_X1 U896 ( .A1(G559), .A2(n807), .ZN(n808) );
  XNOR2_X1 U897 ( .A(n808), .B(n997), .ZN(n817) );
  NAND2_X1 U898 ( .A1(n809), .A2(n817), .ZN(n810) );
  XNOR2_X1 U899 ( .A(n810), .B(KEYINPUT79), .ZN(n811) );
  XOR2_X1 U900 ( .A(n819), .B(n811), .Z(G145) );
  INV_X1 U901 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U902 ( .A(KEYINPUT19), .B(G288), .ZN(n816) );
  XNOR2_X1 U903 ( .A(n819), .B(n1002), .ZN(n812) );
  XNOR2_X1 U904 ( .A(n812), .B(G305), .ZN(n813) );
  XNOR2_X1 U905 ( .A(G166), .B(n813), .ZN(n814) );
  XNOR2_X1 U906 ( .A(n814), .B(G290), .ZN(n815) );
  XNOR2_X1 U907 ( .A(n816), .B(n815), .ZN(n908) );
  XNOR2_X1 U908 ( .A(n817), .B(n908), .ZN(n818) );
  NAND2_X1 U909 ( .A1(n818), .A2(G868), .ZN(n822) );
  NAND2_X1 U910 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U911 ( .A1(n822), .A2(n821), .ZN(G295) );
  NAND2_X1 U912 ( .A1(G2078), .A2(G2084), .ZN(n823) );
  XNOR2_X1 U913 ( .A(n823), .B(KEYINPUT87), .ZN(n824) );
  XNOR2_X1 U914 ( .A(n824), .B(KEYINPUT20), .ZN(n825) );
  NAND2_X1 U915 ( .A1(n825), .A2(G2090), .ZN(n826) );
  XNOR2_X1 U916 ( .A(n826), .B(KEYINPUT21), .ZN(n827) );
  XNOR2_X1 U917 ( .A(n827), .B(KEYINPUT88), .ZN(n828) );
  NAND2_X1 U918 ( .A1(n828), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U919 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U920 ( .A1(G235), .A2(G236), .ZN(n829) );
  XNOR2_X1 U921 ( .A(n829), .B(KEYINPUT89), .ZN(n830) );
  NOR2_X1 U922 ( .A1(G237), .A2(n830), .ZN(n831) );
  XNOR2_X1 U923 ( .A(KEYINPUT90), .B(n831), .ZN(n832) );
  NAND2_X1 U924 ( .A1(n832), .A2(G108), .ZN(n844) );
  NAND2_X1 U925 ( .A1(n844), .A2(G567), .ZN(n837) );
  NOR2_X1 U926 ( .A1(G220), .A2(G219), .ZN(n833) );
  XOR2_X1 U927 ( .A(KEYINPUT22), .B(n833), .Z(n834) );
  NOR2_X1 U928 ( .A1(G218), .A2(n834), .ZN(n835) );
  NAND2_X1 U929 ( .A1(G96), .A2(n835), .ZN(n845) );
  NAND2_X1 U930 ( .A1(n845), .A2(G2106), .ZN(n836) );
  NAND2_X1 U931 ( .A1(n837), .A2(n836), .ZN(n846) );
  NAND2_X1 U932 ( .A1(G483), .A2(G661), .ZN(n838) );
  NOR2_X1 U933 ( .A1(n846), .A2(n838), .ZN(n843) );
  NAND2_X1 U934 ( .A1(n843), .A2(G36), .ZN(n839) );
  XOR2_X1 U935 ( .A(KEYINPUT91), .B(n839), .Z(G176) );
  NAND2_X1 U936 ( .A1(G2106), .A2(n840), .ZN(G217) );
  AND2_X1 U937 ( .A1(G15), .A2(G2), .ZN(n841) );
  NAND2_X1 U938 ( .A1(G661), .A2(n841), .ZN(G259) );
  NAND2_X1 U939 ( .A1(G3), .A2(G1), .ZN(n842) );
  NAND2_X1 U940 ( .A1(n843), .A2(n842), .ZN(G188) );
  INV_X1 U942 ( .A(G108), .ZN(G238) );
  INV_X1 U943 ( .A(G96), .ZN(G221) );
  NOR2_X1 U944 ( .A1(n845), .A2(n844), .ZN(G325) );
  INV_X1 U945 ( .A(G325), .ZN(G261) );
  INV_X1 U946 ( .A(n846), .ZN(G319) );
  XOR2_X1 U947 ( .A(G2096), .B(KEYINPUT43), .Z(n848) );
  XNOR2_X1 U948 ( .A(G2072), .B(KEYINPUT42), .ZN(n847) );
  XNOR2_X1 U949 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U950 ( .A(n849), .B(G2678), .Z(n851) );
  XNOR2_X1 U951 ( .A(G2067), .B(G2090), .ZN(n850) );
  XNOR2_X1 U952 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U953 ( .A(KEYINPUT112), .B(G2100), .Z(n853) );
  XNOR2_X1 U954 ( .A(G2078), .B(G2084), .ZN(n852) );
  XNOR2_X1 U955 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n855), .B(n854), .ZN(G227) );
  XOR2_X1 U957 ( .A(G1976), .B(G1981), .Z(n857) );
  XNOR2_X1 U958 ( .A(G1966), .B(G1956), .ZN(n856) );
  XNOR2_X1 U959 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U960 ( .A(n858), .B(G2474), .Z(n860) );
  XNOR2_X1 U961 ( .A(G1986), .B(G1971), .ZN(n859) );
  XNOR2_X1 U962 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U963 ( .A(KEYINPUT41), .B(G1961), .Z(n862) );
  XNOR2_X1 U964 ( .A(G1996), .B(G1991), .ZN(n861) );
  XNOR2_X1 U965 ( .A(n862), .B(n861), .ZN(n863) );
  XNOR2_X1 U966 ( .A(n864), .B(n863), .ZN(G229) );
  NAND2_X1 U967 ( .A1(G100), .A2(n889), .ZN(n866) );
  NAND2_X1 U968 ( .A1(G112), .A2(n883), .ZN(n865) );
  NAND2_X1 U969 ( .A1(n866), .A2(n865), .ZN(n867) );
  XNOR2_X1 U970 ( .A(n867), .B(KEYINPUT113), .ZN(n869) );
  NAND2_X1 U971 ( .A1(G136), .A2(n888), .ZN(n868) );
  NAND2_X1 U972 ( .A1(n869), .A2(n868), .ZN(n872) );
  NAND2_X1 U973 ( .A1(n884), .A2(G124), .ZN(n870) );
  XOR2_X1 U974 ( .A(KEYINPUT44), .B(n870), .Z(n871) );
  NOR2_X1 U975 ( .A1(n872), .A2(n871), .ZN(G162) );
  XOR2_X1 U976 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n882) );
  NAND2_X1 U977 ( .A1(G139), .A2(n888), .ZN(n874) );
  NAND2_X1 U978 ( .A1(G103), .A2(n889), .ZN(n873) );
  NAND2_X1 U979 ( .A1(n874), .A2(n873), .ZN(n880) );
  NAND2_X1 U980 ( .A1(n884), .A2(G127), .ZN(n875) );
  XNOR2_X1 U981 ( .A(n875), .B(KEYINPUT116), .ZN(n877) );
  NAND2_X1 U982 ( .A1(G115), .A2(n883), .ZN(n876) );
  NAND2_X1 U983 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U984 ( .A(KEYINPUT47), .B(n878), .Z(n879) );
  NOR2_X1 U985 ( .A1(n880), .A2(n879), .ZN(n956) );
  XNOR2_X1 U986 ( .A(n956), .B(G162), .ZN(n881) );
  XNOR2_X1 U987 ( .A(n882), .B(n881), .ZN(n899) );
  XNOR2_X1 U988 ( .A(G160), .B(n942), .ZN(n897) );
  NAND2_X1 U989 ( .A1(G118), .A2(n883), .ZN(n886) );
  NAND2_X1 U990 ( .A1(G130), .A2(n884), .ZN(n885) );
  NAND2_X1 U991 ( .A1(n886), .A2(n885), .ZN(n887) );
  XNOR2_X1 U992 ( .A(KEYINPUT114), .B(n887), .ZN(n895) );
  NAND2_X1 U993 ( .A1(G142), .A2(n888), .ZN(n891) );
  NAND2_X1 U994 ( .A1(G106), .A2(n889), .ZN(n890) );
  NAND2_X1 U995 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U996 ( .A(KEYINPUT45), .B(n892), .ZN(n893) );
  XNOR2_X1 U997 ( .A(KEYINPUT115), .B(n893), .ZN(n894) );
  NOR2_X1 U998 ( .A1(n895), .A2(n894), .ZN(n896) );
  XNOR2_X1 U999 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U1000 ( .A(n899), .B(n898), .Z(n903) );
  XNOR2_X1 U1001 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n903), .B(n902), .ZN(n906) );
  XOR2_X1 U1003 ( .A(n904), .B(G164), .Z(n905) );
  XNOR2_X1 U1004 ( .A(n906), .B(n905), .ZN(n907) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n907), .ZN(G395) );
  XNOR2_X1 U1006 ( .A(G286), .B(n908), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(G171), .B(n997), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(n910), .B(n909), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(n911), .B(n1017), .ZN(n912) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n912), .ZN(G397) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n913) );
  XOR2_X1 U1012 ( .A(KEYINPUT49), .B(n913), .Z(n914) );
  NAND2_X1 U1013 ( .A1(G319), .A2(n914), .ZN(n915) );
  NOR2_X1 U1014 ( .A1(G401), .A2(n915), .ZN(n918) );
  NOR2_X1 U1015 ( .A1(G395), .A2(G397), .ZN(n916) );
  XOR2_X1 U1016 ( .A(KEYINPUT117), .B(n916), .Z(n917) );
  NAND2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  XNOR2_X1 U1019 ( .A(G2090), .B(G35), .ZN(n932) );
  XOR2_X1 U1020 ( .A(G1996), .B(G32), .Z(n919) );
  NAND2_X1 U1021 ( .A1(n919), .A2(G28), .ZN(n929) );
  XNOR2_X1 U1022 ( .A(G2067), .B(G26), .ZN(n921) );
  XNOR2_X1 U1023 ( .A(G33), .B(G2072), .ZN(n920) );
  NOR2_X1 U1024 ( .A1(n921), .A2(n920), .ZN(n927) );
  XOR2_X1 U1025 ( .A(n922), .B(G25), .Z(n925) );
  XNOR2_X1 U1026 ( .A(G27), .B(n923), .ZN(n924) );
  NOR2_X1 U1027 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1028 ( .A1(n927), .A2(n926), .ZN(n928) );
  NOR2_X1 U1029 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1030 ( .A(KEYINPUT53), .B(n930), .ZN(n931) );
  NOR2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n935) );
  XOR2_X1 U1032 ( .A(G2084), .B(G34), .Z(n933) );
  XNOR2_X1 U1033 ( .A(KEYINPUT54), .B(n933), .ZN(n934) );
  NAND2_X1 U1034 ( .A1(n935), .A2(n934), .ZN(n938) );
  NOR2_X1 U1035 ( .A1(G29), .A2(KEYINPUT55), .ZN(n936) );
  NAND2_X1 U1036 ( .A1(n938), .A2(n936), .ZN(n937) );
  NAND2_X1 U1037 ( .A1(G11), .A2(n937), .ZN(n969) );
  INV_X1 U1038 ( .A(KEYINPUT55), .ZN(n963) );
  OR2_X1 U1039 ( .A1(n963), .A2(n938), .ZN(n967) );
  XOR2_X1 U1040 ( .A(G2090), .B(G162), .Z(n939) );
  NOR2_X1 U1041 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1042 ( .A(KEYINPUT51), .B(n941), .Z(n948) );
  NOR2_X1 U1043 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1044 ( .A(KEYINPUT118), .B(n944), .Z(n946) );
  XOR2_X1 U1045 ( .A(G2084), .B(G160), .Z(n945) );
  NOR2_X1 U1046 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1047 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1048 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1049 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1050 ( .A(n953), .B(KEYINPUT119), .ZN(n955) );
  NAND2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n961) );
  XOR2_X1 U1052 ( .A(G2072), .B(n956), .Z(n958) );
  XOR2_X1 U1053 ( .A(G164), .B(G2078), .Z(n957) );
  NOR2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1055 ( .A(KEYINPUT50), .B(n959), .Z(n960) );
  NOR2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(n962), .B(KEYINPUT52), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1059 ( .A1(G29), .A2(n965), .ZN(n966) );
  NAND2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1061 ( .A1(n969), .A2(n968), .ZN(n1027) );
  XNOR2_X1 U1062 ( .A(G20), .B(n970), .ZN(n974) );
  XNOR2_X1 U1063 ( .A(G1341), .B(G19), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(G1981), .B(G6), .ZN(n971) );
  NOR2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n977) );
  XOR2_X1 U1067 ( .A(KEYINPUT59), .B(G1348), .Z(n975) );
  XNOR2_X1 U1068 ( .A(G4), .B(n975), .ZN(n976) );
  NOR2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1070 ( .A(KEYINPUT60), .B(n978), .ZN(n979) );
  XNOR2_X1 U1071 ( .A(n979), .B(KEYINPUT124), .ZN(n982) );
  XNOR2_X1 U1072 ( .A(G1961), .B(G5), .ZN(n980) );
  XNOR2_X1 U1073 ( .A(n980), .B(KEYINPUT123), .ZN(n981) );
  NAND2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(G21), .B(G1966), .ZN(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1077 ( .A(KEYINPUT125), .B(n985), .Z(n992) );
  XOR2_X1 U1078 ( .A(G1976), .B(G23), .Z(n987) );
  XOR2_X1 U1079 ( .A(G1971), .B(G22), .Z(n986) );
  NAND2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n989) );
  XNOR2_X1 U1081 ( .A(G24), .B(G1986), .ZN(n988) );
  NOR2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1083 ( .A(KEYINPUT58), .B(n990), .ZN(n991) );
  NAND2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1085 ( .A(n993), .B(KEYINPUT126), .ZN(n994) );
  XNOR2_X1 U1086 ( .A(KEYINPUT61), .B(n994), .ZN(n995) );
  NOR2_X1 U1087 ( .A1(G16), .A2(n995), .ZN(n1024) );
  XOR2_X1 U1088 ( .A(G16), .B(KEYINPUT120), .Z(n996) );
  XNOR2_X1 U1089 ( .A(KEYINPUT56), .B(n996), .ZN(n1022) );
  XNOR2_X1 U1090 ( .A(n997), .B(G1341), .ZN(n999) );
  XNOR2_X1 U1091 ( .A(G171), .B(G1961), .ZN(n998) );
  NAND2_X1 U1092 ( .A1(n999), .A2(n998), .ZN(n1001) );
  XNOR2_X1 U1093 ( .A(G1971), .B(G303), .ZN(n1000) );
  NOR2_X1 U1094 ( .A1(n1001), .A2(n1000), .ZN(n1016) );
  XNOR2_X1 U1095 ( .A(n1002), .B(G1956), .ZN(n1004) );
  NAND2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1014) );
  XNOR2_X1 U1099 ( .A(G1966), .B(G168), .ZN(n1010) );
  NAND2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1101 ( .A(KEYINPUT121), .B(n1011), .ZN(n1012) );
  XNOR2_X1 U1102 ( .A(KEYINPUT57), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1019) );
  XNOR2_X1 U1105 ( .A(G1348), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(n1020), .B(KEYINPUT122), .ZN(n1021) );
  NOR2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1110 ( .A(KEYINPUT127), .B(n1025), .Z(n1026) );
  NAND2_X1 U1111 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1028), .Z(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

