//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 0 1 1 0 1 0 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 0 0 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n643, new_n644, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n841,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202));
  INV_X1    g001(.A(G169gat), .ZN(new_n203));
  INV_X1    g002(.A(G176gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT23), .ZN(new_n207));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n207), .A2(KEYINPUT25), .A3(new_n208), .ZN(new_n209));
  AND2_X1   g008(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n210));
  NOR2_X1   g009(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n205), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT67), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n212), .B(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G183gat), .ZN(new_n215));
  INV_X1    g014(.A(G190gat), .ZN(new_n216));
  OR3_X1    g015(.A1(new_n215), .A2(new_n216), .A3(KEYINPUT24), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT24), .B1(new_n215), .B2(new_n216), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT69), .B(G183gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(new_n216), .ZN(new_n221));
  AOI211_X1 g020(.A(new_n209), .B(new_n214), .C1(new_n219), .C2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT25), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n207), .B(KEYINPUT65), .ZN(new_n224));
  NOR2_X1   g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n225), .B(KEYINPUT64), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n219), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n224), .A2(new_n208), .A3(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n223), .B1(new_n228), .B2(new_n214), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n222), .B1(new_n229), .B2(KEYINPUT68), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n230), .B1(KEYINPUT68), .B2(new_n229), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n220), .A2(KEYINPUT27), .ZN(new_n232));
  NOR2_X1   g031(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n233));
  XOR2_X1   g032(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n234));
  OAI211_X1 g033(.A(new_n232), .B(new_n233), .C1(new_n215), .C2(new_n234), .ZN(new_n235));
  XOR2_X1   g034(.A(KEYINPUT27), .B(G183gat), .Z(new_n236));
  OAI21_X1  g035(.A(KEYINPUT28), .B1(new_n236), .B2(G190gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n238), .B(KEYINPUT71), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n206), .A2(KEYINPUT72), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n240), .A2(KEYINPUT26), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n208), .B1(new_n240), .B2(KEYINPUT26), .ZN(new_n242));
  OAI221_X1 g041(.A(new_n239), .B1(new_n215), .B2(new_n216), .C1(new_n241), .C2(new_n242), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n231), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(G226gat), .A2(G233gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n231), .A2(new_n243), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT29), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n247), .A2(new_n248), .B1(G226gat), .B2(G233gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G197gat), .B(G204gat), .ZN(new_n251));
  INV_X1    g050(.A(G211gat), .ZN(new_n252));
  INV_X1    g051(.A(G218gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n251), .B1(KEYINPUT22), .B2(new_n254), .ZN(new_n255));
  XOR2_X1   g054(.A(G211gat), .B(G218gat), .Z(new_n256));
  XOR2_X1   g055(.A(new_n255), .B(new_n256), .Z(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n250), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n249), .A2(KEYINPUT78), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n245), .B1(new_n244), .B2(KEYINPUT29), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n247), .A2(G226gat), .A3(G233gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n260), .B1(new_n263), .B2(KEYINPUT78), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n202), .B(new_n259), .C1(new_n264), .C2(new_n258), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT87), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G8gat), .B(G36gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(G64gat), .B(G92gat), .ZN(new_n269));
  XOR2_X1   g068(.A(new_n268), .B(new_n269), .Z(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(KEYINPUT78), .B1(new_n246), .B2(new_n249), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT78), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n261), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(new_n257), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n276), .A2(KEYINPUT87), .A3(new_n202), .A4(new_n259), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n258), .B1(new_n272), .B2(new_n274), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n263), .A2(new_n257), .ZN(new_n279));
  OAI21_X1  g078(.A(KEYINPUT37), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n267), .A2(new_n271), .A3(new_n277), .A4(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT38), .ZN(new_n282));
  XOR2_X1   g081(.A(G141gat), .B(G148gat), .Z(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT79), .ZN(new_n284));
  XNOR2_X1  g083(.A(G155gat), .B(G162gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(G155gat), .ZN(new_n287));
  INV_X1    g086(.A(G162gat), .ZN(new_n288));
  OAI21_X1  g087(.A(KEYINPUT2), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n286), .B(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G113gat), .B(G120gat), .ZN(new_n293));
  XOR2_X1   g092(.A(G127gat), .B(G134gat), .Z(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT74), .ZN(new_n295));
  AOI211_X1 g094(.A(KEYINPUT1), .B(new_n293), .C1(new_n295), .C2(KEYINPUT73), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n293), .A2(KEYINPUT73), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT74), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n298), .A2(KEYINPUT1), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n294), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  OR2_X1    g099(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n292), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n302), .B(KEYINPUT4), .ZN(new_n303));
  INV_X1    g102(.A(new_n301), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT80), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT80), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  OR2_X1    g106(.A1(new_n291), .A2(KEYINPUT3), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n291), .A2(KEYINPUT3), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n305), .A2(new_n307), .A3(new_n308), .A4(new_n309), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n303), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(G225gat), .A2(G233gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n311), .A2(KEYINPUT5), .A3(new_n312), .ZN(new_n313));
  XOR2_X1   g112(.A(G1gat), .B(G29gat), .Z(new_n314));
  XNOR2_X1  g113(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n314), .B(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G57gat), .B(G85gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n316), .B(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n303), .A2(new_n312), .A3(new_n310), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT5), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n305), .A2(new_n307), .A3(new_n291), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n312), .B1(new_n321), .B2(new_n302), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n319), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n313), .A2(new_n318), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n318), .B1(new_n313), .B2(new_n323), .ZN(new_n326));
  OR3_X1    g125(.A1(new_n325), .A2(KEYINPUT6), .A3(new_n326), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n313), .A2(new_n323), .A3(KEYINPUT6), .A4(new_n318), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(KEYINPUT82), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n276), .A2(new_n259), .A3(new_n270), .ZN(new_n331));
  AND2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n275), .A2(new_n257), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT85), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n334), .B1(new_n250), .B2(new_n258), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n263), .A2(KEYINPUT85), .A3(new_n257), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT37), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT86), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT38), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT86), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n341), .B(KEYINPUT37), .C1(new_n333), .C2(new_n337), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n339), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n267), .A2(new_n271), .A3(new_n277), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n282), .B(new_n332), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n271), .B1(new_n278), .B2(new_n279), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n331), .A2(KEYINPUT30), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT30), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n276), .A2(new_n348), .A3(new_n259), .A4(new_n270), .ZN(new_n349));
  AOI21_X1  g148(.A(KEYINPUT84), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n347), .A2(new_n349), .A3(KEYINPUT84), .ZN(new_n352));
  NOR3_X1   g151(.A1(new_n311), .A2(KEYINPUT39), .A3(new_n312), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n353), .A2(new_n318), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n321), .A2(new_n312), .A3(new_n302), .ZN(new_n355));
  OAI211_X1 g154(.A(KEYINPUT39), .B(new_n355), .C1(new_n311), .C2(new_n312), .ZN(new_n356));
  AND2_X1   g155(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n324), .B1(new_n357), .B2(KEYINPUT40), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n358), .B1(KEYINPUT40), .B2(new_n357), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n351), .A2(new_n352), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n258), .B1(new_n308), .B2(new_n248), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n361), .B1(G228gat), .B2(G233gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n255), .A2(new_n256), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n248), .B1(new_n363), .B2(KEYINPUT83), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n364), .B1(new_n257), .B2(KEYINPUT83), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n291), .B1(new_n365), .B2(KEYINPUT3), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT3), .B1(new_n258), .B2(new_n248), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n368), .A2(new_n292), .ZN(new_n369));
  OAI211_X1 g168(.A(G228gat), .B(G233gat), .C1(new_n361), .C2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  XOR2_X1   g170(.A(KEYINPUT31), .B(G50gat), .Z(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G78gat), .B(G106gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n374), .B(G22gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n373), .B(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n345), .A2(new_n360), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n247), .A2(new_n301), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n231), .A2(new_n243), .A3(new_n304), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT34), .ZN(new_n382));
  NAND2_X1  g181(.A1(G227gat), .A2(G233gat), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n382), .B1(new_n381), .B2(new_n383), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n379), .A2(G227gat), .A3(G233gat), .A4(new_n380), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT32), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT33), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  XOR2_X1   g191(.A(G15gat), .B(G43gat), .Z(new_n393));
  XNOR2_X1  g192(.A(G71gat), .B(G99gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n393), .B(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n390), .A2(new_n392), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n395), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n389), .B(KEYINPUT32), .C1(new_n391), .C2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(KEYINPUT77), .B1(new_n388), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n388), .A2(new_n399), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT77), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n387), .A2(new_n402), .A3(new_n396), .A4(new_n398), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n400), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  XOR2_X1   g203(.A(KEYINPUT76), .B(KEYINPUT36), .Z(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n399), .B1(KEYINPUT75), .B2(new_n387), .ZN(new_n407));
  INV_X1    g206(.A(new_n386), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT75), .B1(new_n408), .B2(new_n384), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n409), .A2(new_n396), .A3(new_n398), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT36), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n406), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n347), .A2(new_n349), .ZN(new_n414));
  INV_X1    g213(.A(new_n330), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n377), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n376), .B1(new_n407), .B2(new_n410), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n418), .A2(new_n414), .A3(new_n415), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT35), .ZN(new_n420));
  INV_X1    g219(.A(new_n404), .ZN(new_n421));
  NOR3_X1   g220(.A1(new_n330), .A2(KEYINPUT35), .A3(new_n376), .ZN(new_n422));
  AND3_X1   g221(.A1(new_n347), .A2(new_n349), .A3(KEYINPUT84), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n421), .B(new_n422), .C1(new_n423), .C2(new_n350), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n378), .A2(new_n417), .B1(new_n420), .B2(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT91), .B(G29gat), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT92), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(new_n428), .A3(G36gat), .ZN(new_n429));
  INV_X1    g228(.A(G36gat), .ZN(new_n430));
  OAI21_X1  g229(.A(KEYINPUT92), .B1(new_n426), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(G50gat), .ZN(new_n433));
  INV_X1    g232(.A(G43gat), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n434), .A2(KEYINPUT93), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n434), .A2(KEYINPUT93), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n433), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n434), .A2(G50gat), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT15), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n432), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(G29gat), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n441), .A2(new_n430), .A3(KEYINPUT14), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT14), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n443), .B1(G29gat), .B2(G36gat), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT15), .ZN(new_n446));
  XNOR2_X1  g245(.A(G43gat), .B(G50gat), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT89), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n438), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n434), .A2(G50gat), .ZN(new_n451));
  OAI21_X1  g250(.A(KEYINPUT89), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n445), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n449), .A2(new_n452), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n445), .A2(KEYINPUT90), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT90), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n442), .A2(new_n444), .A3(new_n456), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n429), .A2(new_n431), .A3(new_n455), .A4(new_n457), .ZN(new_n458));
  AOI22_X1  g257(.A1(new_n440), .A2(new_n453), .B1(new_n454), .B2(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(G15gat), .B(G22gat), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n460), .A2(G1gat), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(G8gat), .ZN(new_n463));
  INV_X1    g262(.A(G1gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT16), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  AND3_X1   g265(.A1(new_n462), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n463), .B1(new_n462), .B2(new_n466), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n459), .A2(new_n469), .ZN(new_n470));
  NOR3_X1   g269(.A1(new_n459), .A2(KEYINPUT94), .A3(new_n469), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT94), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n437), .A2(new_n438), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(new_n446), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n474), .A2(new_n453), .A3(new_n429), .A4(new_n431), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n458), .A2(new_n454), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OR2_X1    g276(.A1(new_n467), .A2(new_n468), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n472), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n470), .B1(new_n471), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(G229gat), .A2(G233gat), .ZN(new_n481));
  XOR2_X1   g280(.A(new_n481), .B(KEYINPUT13), .Z(new_n482));
  NAND2_X1  g281(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT94), .B1(new_n459), .B2(new_n469), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n477), .A2(new_n478), .A3(new_n472), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT17), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n475), .A2(new_n476), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n487), .B1(new_n475), .B2(new_n476), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n469), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n486), .A2(new_n490), .A3(KEYINPUT18), .A4(new_n481), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n483), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(G113gat), .B(G141gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n493), .B(new_n494), .ZN(new_n495));
  XOR2_X1   g294(.A(G169gat), .B(G197gat), .Z(new_n496));
  XNOR2_X1  g295(.A(new_n495), .B(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n497), .B(KEYINPUT12), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n486), .A2(new_n481), .A3(new_n490), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT18), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n492), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n498), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n483), .A2(new_n491), .A3(KEYINPUT95), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n501), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT95), .B1(new_n483), .B2(new_n491), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n503), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT96), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI211_X1 g308(.A(KEYINPUT96), .B(new_n503), .C1(new_n505), .C2(new_n506), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n502), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n425), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(G120gat), .B(G148gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(G176gat), .B(G204gat), .ZN(new_n514));
  XOR2_X1   g313(.A(new_n513), .B(new_n514), .Z(new_n515));
  NAND2_X1  g314(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n516), .A2(G85gat), .A3(G92gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(G85gat), .A2(G92gat), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n518), .A2(KEYINPUT100), .A3(KEYINPUT7), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(G99gat), .A2(G106gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT101), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT101), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n523), .A2(G99gat), .A3(G106gat), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n522), .A2(new_n524), .A3(KEYINPUT8), .ZN(new_n525));
  XNOR2_X1  g324(.A(G99gat), .B(G106gat), .ZN(new_n526));
  INV_X1    g325(.A(G85gat), .ZN(new_n527));
  INV_X1    g326(.A(G92gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n520), .A2(new_n525), .A3(new_n526), .A4(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT102), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AOI22_X1  g331(.A1(new_n517), .A2(new_n519), .B1(new_n527), .B2(new_n528), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n533), .A2(KEYINPUT102), .A3(new_n526), .A4(new_n525), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n520), .A2(new_n525), .A3(new_n529), .ZN(new_n536));
  INV_X1    g335(.A(new_n526), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT103), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT103), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n536), .A2(new_n540), .A3(new_n537), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n535), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(G71gat), .A2(G78gat), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT9), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(G64gat), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n546), .A2(G57gat), .ZN(new_n547));
  INV_X1    g346(.A(G57gat), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n548), .A2(G64gat), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n545), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(KEYINPUT97), .B1(new_n550), .B2(KEYINPUT98), .ZN(new_n551));
  XNOR2_X1  g350(.A(G71gat), .B(G78gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n548), .A2(G64gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n546), .A2(G57gat), .ZN(new_n554));
  AOI22_X1  g353(.A1(new_n553), .A2(new_n554), .B1(new_n544), .B2(new_n543), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT97), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n552), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n551), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g357(.A(KEYINPUT97), .B(new_n552), .C1(new_n550), .C2(KEYINPUT98), .ZN(new_n559));
  AND2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n542), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT10), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n558), .A2(new_n559), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n563), .A2(new_n530), .A3(new_n538), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n542), .A2(KEYINPUT104), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT104), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n535), .A2(new_n539), .A3(new_n567), .A4(new_n541), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n560), .A2(new_n562), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n565), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(G230gat), .A2(G233gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT105), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n571), .A2(KEYINPUT105), .A3(new_n572), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n564), .ZN(new_n578));
  INV_X1    g377(.A(new_n572), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n515), .B1(new_n577), .B2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT106), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n573), .A2(new_n515), .A3(new_n580), .ZN(new_n584));
  AOI21_X1  g383(.A(KEYINPUT107), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n577), .A2(new_n580), .ZN(new_n586));
  INV_X1    g385(.A(new_n515), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n582), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AOI211_X1 g387(.A(KEYINPUT106), .B(new_n515), .C1(new_n577), .C2(new_n580), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n584), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT107), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n585), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n563), .A2(KEYINPUT21), .ZN(new_n594));
  NAND2_X1  g393(.A1(G231gat), .A2(G233gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(G127gat), .ZN(new_n597));
  XOR2_X1   g396(.A(G183gat), .B(G211gat), .Z(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n478), .B1(KEYINPUT21), .B2(new_n563), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT99), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(G155gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n601), .B(new_n603), .ZN(new_n604));
  OR2_X1    g403(.A1(new_n599), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n599), .A2(new_n604), .ZN(new_n606));
  AND2_X1   g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G134gat), .B(G162gat), .ZN(new_n608));
  AOI21_X1  g407(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n566), .A2(new_n568), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n612), .B1(new_n489), .B2(new_n488), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n566), .A2(new_n477), .A3(new_n568), .ZN(new_n614));
  NAND3_X1  g413(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(G190gat), .B(G218gat), .Z(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n616), .A2(new_n617), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n611), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  OR2_X1    g420(.A1(new_n616), .A2(new_n617), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n622), .A2(new_n610), .A3(new_n618), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n607), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n593), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n512), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n629), .A2(new_n415), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(new_n464), .ZN(G1324gat));
  NOR2_X1   g430(.A1(new_n423), .A2(new_n350), .ZN(new_n632));
  XOR2_X1   g431(.A(KEYINPUT16), .B(G8gat), .Z(new_n633));
  NAND4_X1  g432(.A1(new_n512), .A2(new_n632), .A3(new_n628), .A4(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n632), .ZN(new_n635));
  OAI21_X1  g434(.A(G8gat), .B1(new_n629), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n634), .ZN(new_n637));
  MUX2_X1   g436(.A(new_n634), .B(new_n637), .S(KEYINPUT42), .Z(G1325gat));
  OR3_X1    g437(.A1(new_n629), .A2(G15gat), .A3(new_n404), .ZN(new_n639));
  INV_X1    g438(.A(new_n413), .ZN(new_n640));
  OAI21_X1  g439(.A(G15gat), .B1(new_n629), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(G1326gat));
  NOR2_X1   g441(.A1(new_n629), .A2(new_n377), .ZN(new_n643));
  XOR2_X1   g442(.A(KEYINPUT43), .B(G22gat), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(G1327gat));
  INV_X1    g444(.A(new_n607), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n646), .A2(new_n624), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n593), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT108), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n512), .A2(new_n330), .A3(new_n426), .A4(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT45), .ZN(new_n652));
  INV_X1    g451(.A(new_n511), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n593), .A2(new_n653), .A3(new_n607), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT110), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n624), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n621), .A2(KEYINPUT110), .A3(new_n623), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n658), .A2(KEYINPUT44), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n378), .A2(new_n417), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT109), .ZN(new_n662));
  AND3_X1   g461(.A1(new_n424), .A2(new_n420), .A3(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n662), .B1(new_n424), .B2(new_n420), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n659), .B1(new_n661), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(KEYINPUT44), .B1(new_n425), .B2(new_n624), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n654), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n668), .A2(new_n330), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n652), .B1(new_n426), .B2(new_n669), .ZN(G1328gat));
  NAND4_X1  g469(.A1(new_n512), .A2(new_n430), .A3(new_n632), .A4(new_n650), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT46), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n430), .B1(new_n668), .B2(new_n632), .ZN(new_n673));
  OR2_X1    g472(.A1(new_n672), .A2(new_n673), .ZN(G1329gat));
  XNOR2_X1  g473(.A(KEYINPUT93), .B(G43gat), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n413), .A2(new_n676), .ZN(new_n677));
  AOI211_X1 g476(.A(new_n654), .B(new_n677), .C1(new_n666), .C2(new_n667), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n512), .A2(new_n650), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n675), .B1(new_n680), .B2(new_n404), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n679), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n682), .ZN(new_n684));
  INV_X1    g483(.A(new_n681), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n684), .B1(new_n685), .B2(new_n678), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n683), .A2(new_n686), .ZN(G1330gat));
  INV_X1    g486(.A(KEYINPUT48), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n433), .B1(new_n668), .B2(new_n376), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n512), .A2(new_n433), .A3(new_n376), .A4(new_n650), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n688), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  AOI211_X1 g491(.A(new_n377), .B(new_n654), .C1(new_n666), .C2(new_n667), .ZN(new_n693));
  OAI211_X1 g492(.A(KEYINPUT48), .B(new_n690), .C1(new_n693), .C2(new_n433), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n694), .ZN(G1331gat));
  NAND2_X1  g494(.A1(new_n424), .A2(new_n420), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(KEYINPUT109), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n424), .A2(new_n420), .A3(new_n662), .ZN(new_n698));
  AOI22_X1  g497(.A1(new_n697), .A2(new_n698), .B1(new_n378), .B2(new_n417), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n593), .A2(new_n653), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n626), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(new_n330), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(G57gat), .ZN(G1332gat));
  INV_X1    g503(.A(KEYINPUT49), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n632), .B1(new_n705), .B2(new_n546), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n706), .B(KEYINPUT112), .Z(new_n707));
  NAND2_X1  g506(.A1(new_n702), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n705), .A2(new_n546), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1333gat));
  INV_X1    g509(.A(G71gat), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n702), .A2(new_n711), .A3(new_n421), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n699), .A2(new_n640), .A3(new_n701), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n712), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT50), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1334gat));
  NAND2_X1  g515(.A1(new_n702), .A2(new_n376), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g517(.A1(new_n700), .A2(new_n607), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n719), .B1(new_n666), .B2(new_n667), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n720), .A2(new_n330), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT51), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n647), .A2(new_n511), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(new_n699), .B2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n723), .ZN(new_n725));
  OAI211_X1 g524(.A(KEYINPUT51), .B(new_n725), .C1(new_n661), .C2(new_n665), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT113), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n724), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n593), .ZN(new_n729));
  OAI211_X1 g528(.A(KEYINPUT113), .B(new_n722), .C1(new_n699), .C2(new_n723), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n330), .A2(new_n527), .ZN(new_n732));
  OAI22_X1  g531(.A1(new_n721), .A2(new_n527), .B1(new_n731), .B2(new_n732), .ZN(G1336gat));
  AOI21_X1  g532(.A(new_n528), .B1(new_n720), .B2(new_n632), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n635), .A2(G92gat), .A3(new_n593), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n736), .B1(new_n724), .B2(new_n726), .ZN(new_n737));
  OAI21_X1  g536(.A(KEYINPUT52), .B1(new_n734), .B2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n719), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT44), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n660), .A2(new_n696), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n740), .B1(new_n741), .B2(new_n625), .ZN(new_n742));
  INV_X1    g541(.A(new_n659), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n699), .A2(new_n743), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n632), .B(new_n739), .C1(new_n742), .C2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G92gat), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n728), .A2(new_n730), .A3(new_n735), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT52), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n738), .A2(new_n749), .ZN(G1337gat));
  NAND2_X1  g549(.A1(new_n720), .A2(new_n413), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G99gat), .ZN(new_n752));
  OR2_X1    g551(.A1(new_n404), .A2(G99gat), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n731), .B2(new_n753), .ZN(G1338gat));
  INV_X1    g553(.A(G106gat), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n755), .B1(new_n720), .B2(new_n376), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n593), .A2(G106gat), .A3(new_n377), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n758), .B1(new_n724), .B2(new_n726), .ZN(new_n759));
  OAI21_X1  g558(.A(KEYINPUT53), .B1(new_n756), .B2(new_n759), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n376), .B(new_n739), .C1(new_n742), .C2(new_n744), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G106gat), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n728), .A2(new_n730), .A3(new_n757), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT53), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n760), .A2(new_n765), .ZN(G1339gat));
  AOI21_X1  g565(.A(KEYINPUT105), .B1(new_n571), .B2(new_n572), .ZN(new_n767));
  AOI211_X1 g566(.A(new_n574), .B(new_n579), .C1(new_n565), .C2(new_n570), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n767), .A2(new_n768), .A3(KEYINPUT54), .ZN(new_n769));
  OAI21_X1  g568(.A(KEYINPUT114), .B1(new_n769), .B2(new_n515), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT54), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n575), .A2(new_n771), .A3(new_n576), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT114), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n772), .A2(new_n773), .A3(new_n587), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n770), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n565), .A2(new_n570), .A3(new_n579), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n573), .A2(KEYINPUT54), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT55), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT116), .ZN(new_n780));
  OR3_X1    g579(.A1(new_n480), .A2(new_n780), .A3(new_n482), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n780), .B1(new_n480), .B2(new_n482), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n486), .A2(new_n490), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n781), .B(new_n782), .C1(new_n481), .C2(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n502), .B1(new_n784), .B2(new_n497), .ZN(new_n785));
  AND3_X1   g584(.A1(new_n656), .A2(new_n657), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n777), .A2(KEYINPUT55), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n787), .B1(new_n770), .B2(new_n774), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT115), .ZN(new_n789));
  INV_X1    g588(.A(new_n584), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n788), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n787), .ZN(new_n792));
  AND3_X1   g591(.A1(new_n772), .A2(new_n773), .A3(new_n587), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n773), .B1(new_n772), .B2(new_n587), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n792), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT115), .B1(new_n795), .B2(new_n584), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n779), .B(new_n786), .C1(new_n791), .C2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT117), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n789), .B1(new_n788), .B2(new_n790), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n795), .A2(KEYINPUT115), .A3(new_n584), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n778), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n802), .A2(KEYINPUT117), .A3(new_n786), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n799), .A2(new_n803), .ZN(new_n804));
  AOI211_X1 g603(.A(new_n511), .B(new_n778), .C1(new_n800), .C2(new_n801), .ZN(new_n805));
  INV_X1    g604(.A(new_n785), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n583), .A2(KEYINPUT107), .A3(new_n584), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n590), .A2(new_n591), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n658), .B1(new_n805), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n646), .B1(new_n804), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n627), .A2(new_n653), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n813), .A2(new_n415), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n418), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n815), .A2(new_n632), .ZN(new_n816));
  INV_X1    g615(.A(G113gat), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n816), .A2(new_n817), .A3(new_n653), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n330), .B(new_n421), .C1(new_n423), .C2(new_n350), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n377), .B(new_n820), .C1(new_n811), .C2(new_n812), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT118), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n812), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n653), .B(new_n779), .C1(new_n791), .C2(new_n796), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n785), .B1(new_n585), .B2(new_n592), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AOI22_X1  g626(.A1(new_n658), .A2(new_n827), .B1(new_n799), .B2(new_n803), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n824), .B1(new_n828), .B2(new_n646), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n829), .A2(KEYINPUT118), .A3(new_n377), .A4(new_n820), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n823), .A2(new_n653), .A3(new_n830), .ZN(new_n831));
  AND3_X1   g630(.A1(new_n831), .A2(KEYINPUT119), .A3(G113gat), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT119), .B1(new_n831), .B2(G113gat), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n818), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT120), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT120), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n818), .B(new_n836), .C1(new_n832), .C2(new_n833), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(G1340gat));
  AOI21_X1  g637(.A(G120gat), .B1(new_n816), .B2(new_n729), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n823), .A2(new_n830), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n729), .A2(G120gat), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n839), .B1(new_n840), .B2(new_n841), .ZN(G1341gat));
  NAND3_X1  g641(.A1(new_n840), .A2(G127gat), .A3(new_n646), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT121), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n843), .A2(new_n844), .ZN(new_n846));
  AOI21_X1  g645(.A(G127gat), .B1(new_n816), .B2(new_n646), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(G1342gat));
  NOR2_X1   g647(.A1(new_n632), .A2(new_n624), .ZN(new_n849));
  INV_X1    g648(.A(G134gat), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(KEYINPUT56), .B1(new_n815), .B2(new_n851), .ZN(new_n852));
  OR3_X1    g651(.A1(new_n815), .A2(KEYINPUT56), .A3(new_n851), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n840), .A2(new_n625), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n852), .B(new_n853), .C1(new_n854), .C2(new_n850), .ZN(G1343gat));
  NAND4_X1  g654(.A1(new_n779), .A2(new_n653), .A3(new_n584), .A4(new_n795), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n625), .B1(new_n826), .B2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n804), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n812), .B1(new_n859), .B2(new_n607), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT57), .B1(new_n860), .B2(new_n377), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n413), .A2(new_n632), .A3(new_n415), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n829), .A2(new_n376), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n861), .B(new_n862), .C1(KEYINPUT57), .C2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(G141gat), .B1(new_n864), .B2(new_n511), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n640), .A2(new_n376), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n866), .B1(new_n814), .B2(KEYINPUT122), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT122), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n868), .B1(new_n813), .B2(new_n415), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n511), .A2(G141gat), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n867), .A2(new_n635), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  XNOR2_X1  g670(.A(KEYINPUT123), .B(KEYINPUT58), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n865), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n872), .B1(new_n865), .B2(new_n871), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n873), .A2(new_n874), .ZN(G1344gat));
  NAND2_X1  g674(.A1(new_n863), .A2(KEYINPUT57), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n862), .A2(new_n729), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT125), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n802), .A2(new_n625), .A3(new_n785), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n607), .B1(new_n857), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n824), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n377), .A2(KEYINPUT57), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n876), .A2(new_n877), .A3(new_n878), .A4(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(G148gat), .ZN(new_n885));
  AOI22_X1  g684(.A1(new_n863), .A2(KEYINPUT57), .B1(new_n881), .B2(new_n882), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n878), .B1(new_n886), .B2(new_n877), .ZN(new_n887));
  OAI21_X1  g686(.A(KEYINPUT59), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT59), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n889), .B(G148gat), .C1(new_n864), .C2(new_n593), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n867), .A2(new_n869), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT124), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n593), .A2(G148gat), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n892), .A2(new_n893), .A3(new_n635), .A4(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n867), .A2(new_n635), .A3(new_n869), .ZN(new_n896));
  INV_X1    g695(.A(new_n894), .ZN(new_n897));
  OAI21_X1  g696(.A(KEYINPUT124), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n891), .A2(new_n899), .ZN(G1345gat));
  OAI21_X1  g699(.A(G155gat), .B1(new_n864), .B2(new_n607), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n646), .A2(new_n287), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n901), .B1(new_n896), .B2(new_n902), .ZN(G1346gat));
  NAND3_X1  g702(.A1(new_n892), .A2(new_n288), .A3(new_n849), .ZN(new_n904));
  OAI21_X1  g703(.A(G162gat), .B1(new_n864), .B2(new_n658), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(G1347gat));
  NAND4_X1  g705(.A1(new_n351), .A2(new_n415), .A3(new_n352), .A4(new_n421), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT126), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n907), .B(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(new_n377), .A3(new_n829), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n910), .A2(new_n203), .A3(new_n511), .ZN(new_n911));
  INV_X1    g710(.A(new_n418), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n632), .A2(new_n415), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n813), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(G169gat), .B1(new_n914), .B2(new_n653), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n911), .A2(new_n915), .ZN(G1348gat));
  OAI21_X1  g715(.A(G176gat), .B1(new_n910), .B2(new_n593), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n914), .A2(new_n204), .A3(new_n729), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(G1349gat));
  INV_X1    g718(.A(new_n236), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n914), .A2(new_n920), .A3(new_n646), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n910), .A2(new_n607), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n921), .B1(new_n922), .B2(new_n220), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT60), .ZN(G1350gat));
  NAND4_X1  g723(.A1(new_n914), .A2(new_n216), .A3(new_n657), .A4(new_n656), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n909), .A2(new_n377), .A3(new_n625), .A4(new_n829), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT61), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n926), .A2(new_n927), .A3(G190gat), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n927), .B1(new_n926), .B2(G190gat), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n925), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT127), .ZN(G1351gat));
  NOR2_X1   g731(.A1(new_n913), .A2(new_n413), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n886), .A2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(G197gat), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n934), .A2(new_n935), .A3(new_n511), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n829), .A2(new_n376), .A3(new_n933), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n937), .A2(new_n511), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n936), .B1(new_n935), .B2(new_n938), .ZN(G1352gat));
  NOR3_X1   g738(.A1(new_n937), .A2(G204gat), .A3(new_n593), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT62), .ZN(new_n941));
  OAI21_X1  g740(.A(G204gat), .B1(new_n934), .B2(new_n593), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(G1353gat));
  NAND3_X1  g742(.A1(new_n886), .A2(new_n646), .A3(new_n933), .ZN(new_n944));
  AND3_X1   g743(.A1(new_n944), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n945));
  AOI21_X1  g744(.A(KEYINPUT63), .B1(new_n944), .B2(G211gat), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n646), .A2(new_n252), .ZN(new_n947));
  OAI22_X1  g746(.A1(new_n945), .A2(new_n946), .B1(new_n937), .B2(new_n947), .ZN(G1354gat));
  OAI21_X1  g747(.A(G218gat), .B1(new_n934), .B2(new_n624), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n656), .A2(new_n253), .A3(new_n657), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n949), .B1(new_n937), .B2(new_n950), .ZN(G1355gat));
endmodule


