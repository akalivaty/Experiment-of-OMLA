

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592;

  XNOR2_X1 U325 ( .A(KEYINPUT91), .B(n402), .ZN(n552) );
  XNOR2_X1 U326 ( .A(n391), .B(n390), .ZN(n549) );
  NAND2_X1 U327 ( .A1(n520), .A2(n575), .ZN(n498) );
  NOR2_X1 U328 ( .A1(n399), .A2(n552), .ZN(n392) );
  INV_X1 U329 ( .A(n570), .ZN(n546) );
  NOR2_X1 U330 ( .A1(n560), .A2(n473), .ZN(n470) );
  AND2_X1 U331 ( .A1(n487), .A2(n463), .ZN(n465) );
  AND2_X1 U332 ( .A1(n293), .A2(n294), .ZN(n459) );
  OR2_X1 U333 ( .A1(n516), .A2(n393), .ZN(n293) );
  OR2_X1 U334 ( .A1(n403), .A2(n402), .ZN(n294) );
  XNOR2_X2 U335 ( .A(n465), .B(n464), .ZN(n473) );
  NOR2_X1 U336 ( .A1(n454), .A2(n531), .ZN(n517) );
  NOR2_X1 U337 ( .A1(n590), .A2(n461), .ZN(n462) );
  XOR2_X1 U338 ( .A(n363), .B(n362), .Z(n560) );
  XOR2_X1 U339 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n295) );
  XOR2_X1 U340 ( .A(n430), .B(n301), .Z(n296) );
  XNOR2_X1 U341 ( .A(n515), .B(n514), .ZN(n550) );
  INV_X1 U342 ( .A(KEYINPUT112), .ZN(n506) );
  XNOR2_X1 U343 ( .A(n506), .B(KEYINPUT47), .ZN(n507) );
  XNOR2_X1 U344 ( .A(n508), .B(n507), .ZN(n513) );
  XNOR2_X1 U345 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n514) );
  XNOR2_X1 U346 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U347 ( .A(n348), .B(n347), .ZN(n475) );
  NOR2_X1 U348 ( .A1(n560), .A2(n559), .ZN(n569) );
  XOR2_X1 U349 ( .A(KEYINPUT2), .B(G162GAT), .Z(n298) );
  XNOR2_X1 U350 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n297) );
  XNOR2_X1 U351 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U352 ( .A(G141GAT), .B(n299), .Z(n380) );
  XOR2_X1 U353 ( .A(G29GAT), .B(G134GAT), .Z(n430) );
  XNOR2_X1 U354 ( .A(G1GAT), .B(G85GAT), .ZN(n300) );
  XNOR2_X1 U355 ( .A(n295), .B(n300), .ZN(n301) );
  NAND2_X1 U356 ( .A1(G225GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U357 ( .A(n296), .B(n302), .ZN(n306) );
  XOR2_X1 U358 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n304) );
  XNOR2_X1 U359 ( .A(KEYINPUT90), .B(KEYINPUT89), .ZN(n303) );
  XNOR2_X1 U360 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U361 ( .A(n306), .B(n305), .Z(n311) );
  XOR2_X1 U362 ( .A(G127GAT), .B(KEYINPUT85), .Z(n308) );
  XNOR2_X1 U363 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n307) );
  XNOR2_X1 U364 ( .A(n308), .B(n307), .ZN(n359) );
  XNOR2_X1 U365 ( .A(G120GAT), .B(G148GAT), .ZN(n309) );
  XNOR2_X1 U366 ( .A(n309), .B(G57GAT), .ZN(n344) );
  XNOR2_X1 U367 ( .A(n359), .B(n344), .ZN(n310) );
  XNOR2_X1 U368 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U369 ( .A(n380), .B(n312), .ZN(n402) );
  XOR2_X1 U370 ( .A(G169GAT), .B(G8GAT), .Z(n381) );
  XOR2_X1 U371 ( .A(G1GAT), .B(KEYINPUT71), .Z(n314) );
  XNOR2_X1 U372 ( .A(G22GAT), .B(G15GAT), .ZN(n313) );
  XNOR2_X1 U373 ( .A(n314), .B(n313), .ZN(n420) );
  XOR2_X1 U374 ( .A(n381), .B(n420), .Z(n316) );
  XNOR2_X1 U375 ( .A(G29GAT), .B(G36GAT), .ZN(n315) );
  XNOR2_X1 U376 ( .A(n316), .B(n315), .ZN(n322) );
  XOR2_X1 U377 ( .A(G43GAT), .B(G50GAT), .Z(n318) );
  XNOR2_X1 U378 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n317) );
  XNOR2_X1 U379 ( .A(n318), .B(n317), .ZN(n429) );
  XOR2_X1 U380 ( .A(n429), .B(KEYINPUT67), .Z(n320) );
  NAND2_X1 U381 ( .A1(G229GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U382 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U383 ( .A(n322), .B(n321), .Z(n330) );
  XOR2_X1 U384 ( .A(KEYINPUT70), .B(G113GAT), .Z(n324) );
  XNOR2_X1 U385 ( .A(G141GAT), .B(G197GAT), .ZN(n323) );
  XNOR2_X1 U386 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U387 ( .A(KEYINPUT69), .B(KEYINPUT30), .Z(n326) );
  XNOR2_X1 U388 ( .A(KEYINPUT68), .B(KEYINPUT29), .ZN(n325) );
  XNOR2_X1 U389 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U390 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U391 ( .A(n330), .B(n329), .ZN(n575) );
  INV_X1 U392 ( .A(n575), .ZN(n534) );
  XNOR2_X1 U393 ( .A(G71GAT), .B(KEYINPUT72), .ZN(n331) );
  XNOR2_X1 U394 ( .A(n331), .B(KEYINPUT13), .ZN(n419) );
  INV_X1 U395 ( .A(n419), .ZN(n333) );
  INV_X1 U396 ( .A(KEYINPUT31), .ZN(n332) );
  NAND2_X1 U397 ( .A1(n333), .A2(n332), .ZN(n335) );
  NAND2_X1 U398 ( .A1(n419), .A2(KEYINPUT31), .ZN(n334) );
  NAND2_X1 U399 ( .A1(n335), .A2(n334), .ZN(n337) );
  AND2_X1 U400 ( .A1(G230GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U401 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U402 ( .A(KEYINPUT74), .B(KEYINPUT32), .Z(n339) );
  XNOR2_X1 U403 ( .A(KEYINPUT73), .B(KEYINPUT33), .ZN(n338) );
  XOR2_X1 U404 ( .A(n339), .B(n338), .Z(n340) );
  XNOR2_X1 U405 ( .A(n341), .B(n340), .ZN(n348) );
  XOR2_X1 U406 ( .A(G64GAT), .B(G92GAT), .Z(n343) );
  XNOR2_X1 U407 ( .A(G176GAT), .B(G204GAT), .ZN(n342) );
  XNOR2_X1 U408 ( .A(n343), .B(n342), .ZN(n386) );
  XNOR2_X1 U409 ( .A(n344), .B(n386), .ZN(n346) );
  XOR2_X1 U410 ( .A(G106GAT), .B(G78GAT), .Z(n369) );
  XOR2_X1 U411 ( .A(G99GAT), .B(G85GAT), .Z(n436) );
  XNOR2_X1 U412 ( .A(n369), .B(n436), .ZN(n345) );
  INV_X1 U413 ( .A(n475), .ZN(n580) );
  NOR2_X1 U414 ( .A1(n534), .A2(n580), .ZN(n463) );
  XOR2_X1 U415 ( .A(G99GAT), .B(G134GAT), .Z(n350) );
  NAND2_X1 U416 ( .A1(G227GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U417 ( .A(n350), .B(n349), .ZN(n363) );
  XOR2_X1 U418 ( .A(G71GAT), .B(G120GAT), .Z(n352) );
  XNOR2_X1 U419 ( .A(G169GAT), .B(G15GAT), .ZN(n351) );
  XNOR2_X1 U420 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U421 ( .A(G176GAT), .B(KEYINPUT20), .Z(n354) );
  XNOR2_X1 U422 ( .A(G43GAT), .B(G190GAT), .ZN(n353) );
  XNOR2_X1 U423 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U424 ( .A(n356), .B(n355), .Z(n361) );
  XOR2_X1 U425 ( .A(G183GAT), .B(KEYINPUT17), .Z(n358) );
  XNOR2_X1 U426 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n357) );
  XNOR2_X1 U427 ( .A(n358), .B(n357), .ZN(n391) );
  XNOR2_X1 U428 ( .A(n359), .B(n391), .ZN(n360) );
  XNOR2_X1 U429 ( .A(n361), .B(n360), .ZN(n362) );
  INV_X1 U430 ( .A(n560), .ZN(n516) );
  XOR2_X1 U431 ( .A(KEYINPUT87), .B(KEYINPUT88), .Z(n365) );
  XNOR2_X1 U432 ( .A(G22GAT), .B(G148GAT), .ZN(n364) );
  XNOR2_X1 U433 ( .A(n365), .B(n364), .ZN(n378) );
  XOR2_X1 U434 ( .A(G204GAT), .B(KEYINPUT24), .Z(n367) );
  XNOR2_X1 U435 ( .A(G50GAT), .B(KEYINPUT86), .ZN(n366) );
  XNOR2_X1 U436 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U437 ( .A(n369), .B(n368), .Z(n371) );
  NAND2_X1 U438 ( .A1(G228GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U439 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U440 ( .A(n372), .B(KEYINPUT22), .Z(n376) );
  XOR2_X1 U441 ( .A(G211GAT), .B(KEYINPUT21), .Z(n374) );
  XNOR2_X1 U442 ( .A(G197GAT), .B(G218GAT), .ZN(n373) );
  XNOR2_X1 U443 ( .A(n374), .B(n373), .ZN(n387) );
  XNOR2_X1 U444 ( .A(n387), .B(KEYINPUT23), .ZN(n375) );
  XNOR2_X1 U445 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U446 ( .A(n378), .B(n377), .Z(n379) );
  XNOR2_X1 U447 ( .A(n380), .B(n379), .ZN(n556) );
  XNOR2_X1 U448 ( .A(n556), .B(KEYINPUT28), .ZN(n454) );
  XOR2_X1 U449 ( .A(KEYINPUT92), .B(n381), .Z(n383) );
  NAND2_X1 U450 ( .A1(G226GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U451 ( .A(n383), .B(n382), .ZN(n385) );
  XNOR2_X1 U452 ( .A(G36GAT), .B(G190GAT), .ZN(n384) );
  XNOR2_X1 U453 ( .A(n384), .B(KEYINPUT79), .ZN(n423) );
  XOR2_X1 U454 ( .A(n385), .B(n423), .Z(n389) );
  XNOR2_X1 U455 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U456 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U457 ( .A(KEYINPUT27), .B(n549), .ZN(n399) );
  XNOR2_X1 U458 ( .A(n392), .B(KEYINPUT93), .ZN(n531) );
  XOR2_X1 U459 ( .A(n517), .B(KEYINPUT94), .Z(n393) );
  NOR2_X1 U460 ( .A1(n560), .A2(n549), .ZN(n394) );
  NOR2_X1 U461 ( .A1(n556), .A2(n394), .ZN(n396) );
  XOR2_X1 U462 ( .A(KEYINPUT25), .B(KEYINPUT96), .Z(n395) );
  XNOR2_X1 U463 ( .A(n396), .B(n395), .ZN(n401) );
  AND2_X1 U464 ( .A1(n556), .A2(n560), .ZN(n398) );
  XNOR2_X1 U465 ( .A(KEYINPUT95), .B(KEYINPUT26), .ZN(n397) );
  XNOR2_X1 U466 ( .A(n398), .B(n397), .ZN(n574) );
  NOR2_X1 U467 ( .A1(n399), .A2(n574), .ZN(n400) );
  NOR2_X1 U468 ( .A1(n401), .A2(n400), .ZN(n403) );
  XOR2_X1 U469 ( .A(G78GAT), .B(G211GAT), .Z(n405) );
  XNOR2_X1 U470 ( .A(G127GAT), .B(G155GAT), .ZN(n404) );
  XNOR2_X1 U471 ( .A(n405), .B(n404), .ZN(n409) );
  XOR2_X1 U472 ( .A(KEYINPUT12), .B(G64GAT), .Z(n407) );
  XNOR2_X1 U473 ( .A(G8GAT), .B(G183GAT), .ZN(n406) );
  XNOR2_X1 U474 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U475 ( .A(n409), .B(n408), .Z(n414) );
  XOR2_X1 U476 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n411) );
  NAND2_X1 U477 ( .A1(G231GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U478 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U479 ( .A(KEYINPUT82), .B(n412), .ZN(n413) );
  XNOR2_X1 U480 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U481 ( .A(KEYINPUT83), .B(KEYINPUT81), .Z(n416) );
  XNOR2_X1 U482 ( .A(G57GAT), .B(KEYINPUT80), .ZN(n415) );
  XNOR2_X1 U483 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U484 ( .A(n418), .B(n417), .Z(n422) );
  XNOR2_X1 U485 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U486 ( .A(n422), .B(n421), .ZN(n542) );
  INV_X1 U487 ( .A(n542), .ZN(n583) );
  XOR2_X1 U488 ( .A(n423), .B(KEYINPUT76), .Z(n428) );
  XOR2_X1 U489 ( .A(KEYINPUT78), .B(KEYINPUT75), .Z(n425) );
  XNOR2_X1 U490 ( .A(G162GAT), .B(KEYINPUT11), .ZN(n424) );
  XNOR2_X1 U491 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U492 ( .A(n426), .B(KEYINPUT66), .ZN(n427) );
  XNOR2_X1 U493 ( .A(n428), .B(n427), .ZN(n442) );
  XOR2_X1 U494 ( .A(n430), .B(n429), .Z(n432) );
  NAND2_X1 U495 ( .A1(G232GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U496 ( .A(n432), .B(n431), .ZN(n440) );
  XOR2_X1 U497 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n434) );
  XNOR2_X1 U498 ( .A(G106GAT), .B(G92GAT), .ZN(n433) );
  XNOR2_X1 U499 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U500 ( .A(n435), .B(KEYINPUT77), .Z(n438) );
  XNOR2_X1 U501 ( .A(G218GAT), .B(n436), .ZN(n437) );
  XNOR2_X1 U502 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U503 ( .A(n440), .B(n439), .Z(n441) );
  XNOR2_X1 U504 ( .A(n442), .B(n441), .ZN(n570) );
  NAND2_X1 U505 ( .A1(n583), .A2(n546), .ZN(n443) );
  XNOR2_X1 U506 ( .A(n443), .B(KEYINPUT84), .ZN(n444) );
  XNOR2_X1 U507 ( .A(n444), .B(KEYINPUT16), .ZN(n445) );
  NOR2_X1 U508 ( .A1(n459), .A2(n445), .ZN(n476) );
  NAND2_X1 U509 ( .A1(n463), .A2(n476), .ZN(n455) );
  NOR2_X1 U510 ( .A1(n552), .A2(n455), .ZN(n447) );
  XNOR2_X1 U511 ( .A(KEYINPUT34), .B(KEYINPUT97), .ZN(n446) );
  XNOR2_X1 U512 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U513 ( .A(G1GAT), .B(n448), .ZN(G1324GAT) );
  NOR2_X1 U514 ( .A1(n549), .A2(n455), .ZN(n449) );
  XOR2_X1 U515 ( .A(G8GAT), .B(n449), .Z(G1325GAT) );
  NOR2_X1 U516 ( .A1(n455), .A2(n560), .ZN(n453) );
  XOR2_X1 U517 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n451) );
  XNOR2_X1 U518 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n450) );
  XNOR2_X1 U519 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U520 ( .A(n453), .B(n452), .ZN(G1326GAT) );
  INV_X1 U521 ( .A(n454), .ZN(n495) );
  NOR2_X1 U522 ( .A1(n495), .A2(n455), .ZN(n457) );
  XNOR2_X1 U523 ( .A(KEYINPUT100), .B(KEYINPUT101), .ZN(n456) );
  XNOR2_X1 U524 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U525 ( .A(G22GAT), .B(n458), .ZN(G1327GAT) );
  XNOR2_X1 U526 ( .A(KEYINPUT36), .B(n546), .ZN(n590) );
  NOR2_X1 U527 ( .A1(n459), .A2(n583), .ZN(n460) );
  XOR2_X1 U528 ( .A(KEYINPUT102), .B(n460), .Z(n461) );
  XOR2_X1 U529 ( .A(KEYINPUT37), .B(n462), .Z(n487) );
  XNOR2_X1 U530 ( .A(KEYINPUT103), .B(KEYINPUT38), .ZN(n464) );
  NOR2_X1 U531 ( .A1(n552), .A2(n473), .ZN(n468) );
  XNOR2_X1 U532 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n466) );
  XNOR2_X1 U533 ( .A(n466), .B(KEYINPUT104), .ZN(n467) );
  XNOR2_X1 U534 ( .A(n468), .B(n467), .ZN(G1328GAT) );
  NOR2_X1 U535 ( .A1(n473), .A2(n549), .ZN(n469) );
  XOR2_X1 U536 ( .A(G36GAT), .B(n469), .Z(G1329GAT) );
  XNOR2_X1 U537 ( .A(KEYINPUT40), .B(KEYINPUT105), .ZN(n471) );
  XNOR2_X1 U538 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U539 ( .A(G43GAT), .B(n472), .ZN(G1330GAT) );
  NOR2_X1 U540 ( .A1(n473), .A2(n495), .ZN(n474) );
  XOR2_X1 U541 ( .A(G50GAT), .B(n474), .Z(G1331GAT) );
  XOR2_X1 U542 ( .A(n475), .B(KEYINPUT41), .Z(n536) );
  NOR2_X1 U543 ( .A1(n575), .A2(n536), .ZN(n486) );
  NAND2_X1 U544 ( .A1(n486), .A2(n476), .ZN(n482) );
  NOR2_X1 U545 ( .A1(n552), .A2(n482), .ZN(n477) );
  XOR2_X1 U546 ( .A(n477), .B(KEYINPUT42), .Z(n478) );
  XNOR2_X1 U547 ( .A(G57GAT), .B(n478), .ZN(G1332GAT) );
  NOR2_X1 U548 ( .A1(n549), .A2(n482), .ZN(n479) );
  XOR2_X1 U549 ( .A(KEYINPUT106), .B(n479), .Z(n480) );
  XNOR2_X1 U550 ( .A(G64GAT), .B(n480), .ZN(G1333GAT) );
  NOR2_X1 U551 ( .A1(n560), .A2(n482), .ZN(n481) );
  XOR2_X1 U552 ( .A(G71GAT), .B(n481), .Z(G1334GAT) );
  NOR2_X1 U553 ( .A1(n495), .A2(n482), .ZN(n484) );
  XNOR2_X1 U554 ( .A(KEYINPUT43), .B(KEYINPUT107), .ZN(n483) );
  XNOR2_X1 U555 ( .A(n484), .B(n483), .ZN(n485) );
  XOR2_X1 U556 ( .A(G78GAT), .B(n485), .Z(G1335GAT) );
  NAND2_X1 U557 ( .A1(n487), .A2(n486), .ZN(n494) );
  NOR2_X1 U558 ( .A1(n552), .A2(n494), .ZN(n488) );
  XOR2_X1 U559 ( .A(G85GAT), .B(n488), .Z(G1336GAT) );
  NOR2_X1 U560 ( .A1(n549), .A2(n494), .ZN(n489) );
  XOR2_X1 U561 ( .A(G92GAT), .B(n489), .Z(G1337GAT) );
  NOR2_X1 U562 ( .A1(n560), .A2(n494), .ZN(n490) );
  XOR2_X1 U563 ( .A(KEYINPUT108), .B(n490), .Z(n491) );
  XNOR2_X1 U564 ( .A(G99GAT), .B(n491), .ZN(G1338GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT109), .B(KEYINPUT44), .Z(n493) );
  XNOR2_X1 U566 ( .A(G106GAT), .B(KEYINPUT110), .ZN(n492) );
  XNOR2_X1 U567 ( .A(n493), .B(n492), .ZN(n497) );
  NOR2_X1 U568 ( .A1(n495), .A2(n494), .ZN(n496) );
  XOR2_X1 U569 ( .A(n497), .B(n496), .Z(G1339GAT) );
  INV_X1 U570 ( .A(n536), .ZN(n520) );
  XOR2_X1 U571 ( .A(KEYINPUT46), .B(KEYINPUT111), .Z(n499) );
  NAND2_X1 U572 ( .A1(n498), .A2(n499), .ZN(n503) );
  INV_X1 U573 ( .A(n498), .ZN(n501) );
  INV_X1 U574 ( .A(n499), .ZN(n500) );
  NAND2_X1 U575 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U576 ( .A1(n503), .A2(n502), .ZN(n505) );
  NAND2_X1 U577 ( .A1(n542), .A2(n546), .ZN(n504) );
  NOR2_X1 U578 ( .A1(n505), .A2(n504), .ZN(n508) );
  NOR2_X1 U579 ( .A1(n542), .A2(n590), .ZN(n509) );
  XNOR2_X1 U580 ( .A(KEYINPUT45), .B(n509), .ZN(n510) );
  NAND2_X1 U581 ( .A1(n510), .A2(n475), .ZN(n511) );
  NOR2_X1 U582 ( .A1(n511), .A2(n575), .ZN(n512) );
  NOR2_X1 U583 ( .A1(n513), .A2(n512), .ZN(n515) );
  NAND2_X1 U584 ( .A1(n517), .A2(n516), .ZN(n518) );
  NOR2_X1 U585 ( .A1(n550), .A2(n518), .ZN(n527) );
  NAND2_X1 U586 ( .A1(n527), .A2(n575), .ZN(n519) );
  XNOR2_X1 U587 ( .A(n519), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U588 ( .A(G120GAT), .B(KEYINPUT49), .Z(n522) );
  NAND2_X1 U589 ( .A1(n527), .A2(n520), .ZN(n521) );
  XNOR2_X1 U590 ( .A(n522), .B(n521), .ZN(G1341GAT) );
  XNOR2_X1 U591 ( .A(G127GAT), .B(KEYINPUT114), .ZN(n526) );
  XOR2_X1 U592 ( .A(KEYINPUT113), .B(KEYINPUT50), .Z(n524) );
  NAND2_X1 U593 ( .A1(n527), .A2(n583), .ZN(n523) );
  XNOR2_X1 U594 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U595 ( .A(n526), .B(n525), .ZN(G1342GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n529) );
  NAND2_X1 U597 ( .A1(n527), .A2(n570), .ZN(n528) );
  XNOR2_X1 U598 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U599 ( .A(G134GAT), .B(n530), .Z(G1343GAT) );
  NOR2_X1 U600 ( .A1(n574), .A2(n531), .ZN(n533) );
  INV_X1 U601 ( .A(n550), .ZN(n532) );
  NAND2_X1 U602 ( .A1(n533), .A2(n532), .ZN(n545) );
  NOR2_X1 U603 ( .A1(n534), .A2(n545), .ZN(n535) );
  XOR2_X1 U604 ( .A(G141GAT), .B(n535), .Z(G1344GAT) );
  NOR2_X1 U605 ( .A1(n536), .A2(n545), .ZN(n541) );
  XOR2_X1 U606 ( .A(KEYINPUT117), .B(KEYINPUT53), .Z(n538) );
  XNOR2_X1 U607 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n537) );
  XNOR2_X1 U608 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U609 ( .A(KEYINPUT116), .B(n539), .ZN(n540) );
  XNOR2_X1 U610 ( .A(n541), .B(n540), .ZN(G1345GAT) );
  NOR2_X1 U611 ( .A1(n542), .A2(n545), .ZN(n543) );
  XOR2_X1 U612 ( .A(KEYINPUT118), .B(n543), .Z(n544) );
  XNOR2_X1 U613 ( .A(G155GAT), .B(n544), .ZN(G1346GAT) );
  NOR2_X1 U614 ( .A1(n546), .A2(n545), .ZN(n548) );
  XNOR2_X1 U615 ( .A(G162GAT), .B(KEYINPUT119), .ZN(n547) );
  XNOR2_X1 U616 ( .A(n548), .B(n547), .ZN(G1347GAT) );
  XOR2_X1 U617 ( .A(G169GAT), .B(KEYINPUT121), .Z(n562) );
  NOR2_X1 U618 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n551), .B(KEYINPUT54), .ZN(n553) );
  NAND2_X1 U620 ( .A1(n553), .A2(n552), .ZN(n555) );
  INV_X1 U621 ( .A(KEYINPUT65), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n573) );
  OR2_X1 U623 ( .A1(n573), .A2(n556), .ZN(n558) );
  XOR2_X1 U624 ( .A(KEYINPUT120), .B(KEYINPUT55), .Z(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(n559) );
  NAND2_X1 U626 ( .A1(n569), .A2(n575), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(G1348GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n564) );
  XNOR2_X1 U629 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(n565) );
  XOR2_X1 U631 ( .A(KEYINPUT56), .B(n565), .Z(n567) );
  NAND2_X1 U632 ( .A1(n569), .A2(n520), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(G1349GAT) );
  NAND2_X1 U634 ( .A1(n583), .A2(n569), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n568), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(KEYINPUT58), .ZN(n572) );
  XNOR2_X1 U638 ( .A(G190GAT), .B(n572), .ZN(G1351GAT) );
  NOR2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n588) );
  NAND2_X1 U640 ( .A1(n588), .A2(n575), .ZN(n579) );
  XOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n577) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U645 ( .A(G204GAT), .B(KEYINPUT61), .Z(n582) );
  NAND2_X1 U646 ( .A1(n588), .A2(n580), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  XOR2_X1 U648 ( .A(G211GAT), .B(KEYINPUT125), .Z(n585) );
  NAND2_X1 U649 ( .A1(n588), .A2(n583), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1354GAT) );
  XOR2_X1 U651 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n587) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n586) );
  XNOR2_X1 U653 ( .A(n587), .B(n586), .ZN(n592) );
  INV_X1 U654 ( .A(n588), .ZN(n589) );
  NOR2_X1 U655 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U656 ( .A(n592), .B(n591), .Z(G1355GAT) );
endmodule

