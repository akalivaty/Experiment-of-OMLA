

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591;

  XNOR2_X2 U324 ( .A(n452), .B(KEYINPUT112), .ZN(n546) );
  NOR2_X2 U325 ( .A1(n451), .A2(n472), .ZN(n452) );
  NOR2_X1 U326 ( .A1(n483), .A2(n422), .ZN(n423) );
  XNOR2_X1 U327 ( .A(KEYINPUT109), .B(KEYINPUT47), .ZN(n389) );
  XNOR2_X1 U328 ( .A(n400), .B(n372), .ZN(n373) );
  XNOR2_X1 U329 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U330 ( .A(KEYINPUT48), .B(n399), .ZN(n457) );
  XOR2_X1 U331 ( .A(n387), .B(n386), .Z(n490) );
  XNOR2_X1 U332 ( .A(n314), .B(n313), .ZN(n393) );
  XNOR2_X1 U333 ( .A(n312), .B(n311), .ZN(n313) );
  NOR2_X1 U334 ( .A1(n465), .A2(n472), .ZN(n572) );
  XOR2_X1 U335 ( .A(n421), .B(n420), .Z(n531) );
  XOR2_X2 U336 ( .A(n393), .B(n315), .Z(n568) );
  XOR2_X1 U337 ( .A(G92GAT), .B(G106GAT), .Z(n292) );
  XNOR2_X1 U338 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U339 ( .A(n350), .B(n349), .ZN(n368) );
  XNOR2_X1 U340 ( .A(n390), .B(n389), .ZN(n398) );
  INV_X1 U341 ( .A(G162GAT), .ZN(n370) );
  XNOR2_X1 U342 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U343 ( .A(n459), .B(KEYINPUT119), .ZN(n460) );
  INV_X1 U344 ( .A(KEYINPUT36), .ZN(n391) );
  XNOR2_X1 U345 ( .A(n384), .B(n383), .ZN(n387) );
  XNOR2_X1 U346 ( .A(n560), .B(n391), .ZN(n588) );
  XNOR2_X1 U347 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U348 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U349 ( .A(n469), .B(n468), .ZN(G1351GAT) );
  XNOR2_X1 U350 ( .A(G57GAT), .B(KEYINPUT69), .ZN(n293) );
  XNOR2_X1 U351 ( .A(n293), .B(KEYINPUT13), .ZN(n354) );
  XNOR2_X1 U352 ( .A(n354), .B(G85GAT), .ZN(n295) );
  AND2_X1 U353 ( .A1(G230GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U354 ( .A(n295), .B(n294), .ZN(n297) );
  XNOR2_X1 U355 ( .A(G204GAT), .B(G92GAT), .ZN(n296) );
  XNOR2_X1 U356 ( .A(n296), .B(G64GAT), .ZN(n320) );
  NAND2_X1 U357 ( .A1(n297), .A2(n320), .ZN(n301) );
  INV_X1 U358 ( .A(n297), .ZN(n299) );
  INV_X1 U359 ( .A(n320), .ZN(n298) );
  NAND2_X1 U360 ( .A1(n299), .A2(n298), .ZN(n300) );
  NAND2_X1 U361 ( .A1(n301), .A2(n300), .ZN(n305) );
  XOR2_X1 U362 ( .A(G78GAT), .B(G148GAT), .Z(n303) );
  XNOR2_X1 U363 ( .A(G106GAT), .B(KEYINPUT70), .ZN(n302) );
  XNOR2_X1 U364 ( .A(n303), .B(n302), .ZN(n428) );
  XOR2_X1 U365 ( .A(G176GAT), .B(n428), .Z(n304) );
  XNOR2_X1 U366 ( .A(n305), .B(n304), .ZN(n307) );
  INV_X1 U367 ( .A(KEYINPUT32), .ZN(n306) );
  XNOR2_X1 U368 ( .A(n307), .B(n306), .ZN(n314) );
  XNOR2_X1 U369 ( .A(G99GAT), .B(G71GAT), .ZN(n308) );
  XNOR2_X1 U370 ( .A(n308), .B(G120GAT), .ZN(n441) );
  XNOR2_X1 U371 ( .A(n441), .B(KEYINPUT73), .ZN(n312) );
  XOR2_X1 U372 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n310) );
  XNOR2_X1 U373 ( .A(KEYINPUT72), .B(KEYINPUT71), .ZN(n309) );
  XOR2_X1 U374 ( .A(n310), .B(n309), .Z(n311) );
  XOR2_X1 U375 ( .A(KEYINPUT41), .B(KEYINPUT64), .Z(n315) );
  XOR2_X1 U376 ( .A(KEYINPUT89), .B(KEYINPUT88), .Z(n319) );
  XOR2_X1 U377 ( .A(G36GAT), .B(G8GAT), .Z(n342) );
  NAND2_X1 U378 ( .A1(G226GAT), .A2(G233GAT), .ZN(n316) );
  XOR2_X1 U379 ( .A(G183GAT), .B(G211GAT), .Z(n357) );
  XNOR2_X1 U380 ( .A(n316), .B(n357), .ZN(n317) );
  XNOR2_X1 U381 ( .A(n342), .B(n317), .ZN(n318) );
  XNOR2_X1 U382 ( .A(n319), .B(n318), .ZN(n321) );
  XOR2_X1 U383 ( .A(n321), .B(n320), .Z(n330) );
  XOR2_X1 U384 ( .A(KEYINPUT81), .B(KEYINPUT18), .Z(n323) );
  XNOR2_X1 U385 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n322) );
  XNOR2_X1 U386 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U387 ( .A(n324), .B(KEYINPUT19), .Z(n326) );
  XNOR2_X1 U388 ( .A(G169GAT), .B(G176GAT), .ZN(n325) );
  XNOR2_X1 U389 ( .A(n326), .B(n325), .ZN(n450) );
  XOR2_X1 U390 ( .A(KEYINPUT83), .B(KEYINPUT21), .Z(n328) );
  XNOR2_X1 U391 ( .A(G197GAT), .B(G218GAT), .ZN(n327) );
  XNOR2_X1 U392 ( .A(n328), .B(n327), .ZN(n424) );
  XNOR2_X1 U393 ( .A(n450), .B(n424), .ZN(n329) );
  XNOR2_X1 U394 ( .A(n330), .B(n329), .ZN(n533) );
  XOR2_X1 U395 ( .A(n533), .B(KEYINPUT90), .Z(n331) );
  XNOR2_X1 U396 ( .A(KEYINPUT27), .B(n331), .ZN(n483) );
  XNOR2_X1 U397 ( .A(G43GAT), .B(KEYINPUT7), .ZN(n332) );
  XNOR2_X1 U398 ( .A(n332), .B(G29GAT), .ZN(n333) );
  XOR2_X1 U399 ( .A(n333), .B(KEYINPUT67), .Z(n335) );
  XNOR2_X1 U400 ( .A(G50GAT), .B(KEYINPUT8), .ZN(n334) );
  XOR2_X1 U401 ( .A(n335), .B(n334), .Z(n385) );
  XOR2_X1 U402 ( .A(G197GAT), .B(G15GAT), .Z(n337) );
  XNOR2_X1 U403 ( .A(G169GAT), .B(G113GAT), .ZN(n336) );
  XNOR2_X1 U404 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U405 ( .A(n385), .B(n338), .Z(n346) );
  XOR2_X1 U406 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n340) );
  NAND2_X1 U407 ( .A1(G229GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U408 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U409 ( .A(n341), .B(G141GAT), .Z(n344) );
  XOR2_X1 U410 ( .A(G22GAT), .B(G1GAT), .Z(n365) );
  XNOR2_X1 U411 ( .A(n342), .B(n365), .ZN(n343) );
  XNOR2_X1 U412 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U413 ( .A(n346), .B(n345), .Z(n577) );
  INV_X1 U414 ( .A(n577), .ZN(n553) );
  AND2_X1 U415 ( .A1(n553), .A2(n568), .ZN(n350) );
  XNOR2_X1 U416 ( .A(KEYINPUT107), .B(KEYINPUT46), .ZN(n348) );
  INV_X1 U417 ( .A(KEYINPUT106), .ZN(n347) );
  XOR2_X1 U418 ( .A(KEYINPUT76), .B(KEYINPUT12), .Z(n356) );
  XOR2_X1 U419 ( .A(KEYINPUT14), .B(KEYINPUT77), .Z(n352) );
  XNOR2_X1 U420 ( .A(G8GAT), .B(KEYINPUT15), .ZN(n351) );
  XNOR2_X1 U421 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U422 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U423 ( .A(n356), .B(n355), .ZN(n361) );
  XOR2_X1 U424 ( .A(G15GAT), .B(G127GAT), .Z(n445) );
  XOR2_X1 U425 ( .A(n357), .B(n445), .Z(n359) );
  NAND2_X1 U426 ( .A1(G231GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U427 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U428 ( .A(n361), .B(n360), .Z(n367) );
  XOR2_X1 U429 ( .A(G64GAT), .B(G78GAT), .Z(n363) );
  XNOR2_X1 U430 ( .A(G71GAT), .B(G155GAT), .ZN(n362) );
  XNOR2_X1 U431 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U432 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U433 ( .A(n367), .B(n366), .Z(n558) );
  XOR2_X1 U434 ( .A(KEYINPUT105), .B(n558), .Z(n571) );
  NOR2_X1 U435 ( .A1(n368), .A2(n571), .ZN(n369) );
  XNOR2_X1 U436 ( .A(n369), .B(KEYINPUT108), .ZN(n388) );
  XOR2_X1 U437 ( .A(G134GAT), .B(G85GAT), .Z(n400) );
  NAND2_X1 U438 ( .A1(G232GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U439 ( .A(G190GAT), .B(n373), .ZN(n384) );
  XOR2_X1 U440 ( .A(KEYINPUT11), .B(KEYINPUT66), .Z(n375) );
  XNOR2_X1 U441 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n374) );
  XNOR2_X1 U442 ( .A(n375), .B(n374), .ZN(n378) );
  XNOR2_X1 U443 ( .A(G36GAT), .B(G99GAT), .ZN(n376) );
  XNOR2_X1 U444 ( .A(n292), .B(n376), .ZN(n377) );
  XOR2_X1 U445 ( .A(n378), .B(n377), .Z(n382) );
  XOR2_X1 U446 ( .A(KEYINPUT74), .B(KEYINPUT9), .Z(n380) );
  XNOR2_X1 U447 ( .A(KEYINPUT65), .B(KEYINPUT75), .ZN(n379) );
  XNOR2_X1 U448 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U449 ( .A(n382), .B(n381), .ZN(n383) );
  INV_X1 U450 ( .A(n385), .ZN(n386) );
  NAND2_X1 U451 ( .A1(n388), .A2(n490), .ZN(n390) );
  XOR2_X1 U452 ( .A(n577), .B(KEYINPUT68), .Z(n563) );
  INV_X1 U453 ( .A(n558), .ZN(n585) );
  INV_X1 U454 ( .A(n490), .ZN(n560) );
  NOR2_X1 U455 ( .A1(n585), .A2(n588), .ZN(n392) );
  XNOR2_X1 U456 ( .A(n392), .B(KEYINPUT45), .ZN(n394) );
  BUF_X1 U457 ( .A(n393), .Z(n582) );
  NAND2_X1 U458 ( .A1(n394), .A2(n582), .ZN(n395) );
  NOR2_X1 U459 ( .A1(n563), .A2(n395), .ZN(n396) );
  XOR2_X1 U460 ( .A(KEYINPUT110), .B(n396), .Z(n397) );
  NAND2_X1 U461 ( .A1(n398), .A2(n397), .ZN(n399) );
  XOR2_X1 U462 ( .A(n400), .B(G127GAT), .Z(n403) );
  XNOR2_X1 U463 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n401) );
  XNOR2_X1 U464 ( .A(n401), .B(KEYINPUT79), .ZN(n442) );
  XNOR2_X1 U465 ( .A(G29GAT), .B(n442), .ZN(n402) );
  XNOR2_X1 U466 ( .A(n403), .B(n402), .ZN(n416) );
  XOR2_X1 U467 ( .A(G57GAT), .B(G148GAT), .Z(n405) );
  XNOR2_X1 U468 ( .A(G1GAT), .B(G120GAT), .ZN(n404) );
  XNOR2_X1 U469 ( .A(n405), .B(n404), .ZN(n409) );
  XOR2_X1 U470 ( .A(KEYINPUT86), .B(KEYINPUT4), .Z(n407) );
  XNOR2_X1 U471 ( .A(KEYINPUT85), .B(KEYINPUT5), .ZN(n406) );
  XNOR2_X1 U472 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U473 ( .A(n409), .B(n408), .Z(n414) );
  XOR2_X1 U474 ( .A(KEYINPUT6), .B(KEYINPUT87), .Z(n411) );
  NAND2_X1 U475 ( .A1(G225GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U476 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U477 ( .A(KEYINPUT1), .B(n412), .ZN(n413) );
  XNOR2_X1 U478 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U479 ( .A(n416), .B(n415), .ZN(n421) );
  XOR2_X1 U480 ( .A(KEYINPUT2), .B(G162GAT), .Z(n418) );
  XNOR2_X1 U481 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n417) );
  XNOR2_X1 U482 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U483 ( .A(G141GAT), .B(n419), .ZN(n425) );
  INV_X1 U484 ( .A(n425), .ZN(n420) );
  NAND2_X1 U485 ( .A1(n457), .A2(n531), .ZN(n422) );
  XOR2_X1 U486 ( .A(KEYINPUT111), .B(n423), .Z(n551) );
  XOR2_X1 U487 ( .A(KEYINPUT24), .B(KEYINPUT84), .Z(n427) );
  XOR2_X1 U488 ( .A(n425), .B(n424), .Z(n426) );
  XNOR2_X1 U489 ( .A(n427), .B(n426), .ZN(n432) );
  XOR2_X1 U490 ( .A(G22GAT), .B(n428), .Z(n430) );
  NAND2_X1 U491 ( .A1(G228GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U492 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U493 ( .A(n432), .B(n431), .Z(n437) );
  XOR2_X1 U494 ( .A(G204GAT), .B(G211GAT), .Z(n434) );
  XNOR2_X1 U495 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n433) );
  XNOR2_X1 U496 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U497 ( .A(G50GAT), .B(n435), .ZN(n436) );
  XNOR2_X1 U498 ( .A(n437), .B(n436), .ZN(n479) );
  XOR2_X1 U499 ( .A(n479), .B(KEYINPUT28), .Z(n537) );
  INV_X1 U500 ( .A(n537), .ZN(n474) );
  NAND2_X1 U501 ( .A1(n551), .A2(n474), .ZN(n451) );
  XOR2_X1 U502 ( .A(KEYINPUT80), .B(G183GAT), .Z(n439) );
  NAND2_X1 U503 ( .A1(G227GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U504 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U505 ( .A(n440), .B(KEYINPUT20), .Z(n444) );
  XNOR2_X1 U506 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U507 ( .A(n444), .B(n443), .ZN(n446) );
  XOR2_X1 U508 ( .A(n446), .B(n445), .Z(n448) );
  XNOR2_X1 U509 ( .A(G43GAT), .B(G134GAT), .ZN(n447) );
  XNOR2_X1 U510 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X2 U511 ( .A(n450), .B(n449), .Z(n535) );
  INV_X1 U512 ( .A(n535), .ZN(n472) );
  NAND2_X1 U513 ( .A1(n568), .A2(n546), .ZN(n456) );
  XOR2_X1 U514 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n454) );
  XOR2_X1 U515 ( .A(G120GAT), .B(KEYINPUT114), .Z(n453) );
  XNOR2_X1 U516 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U517 ( .A(n456), .B(n455), .ZN(G1341GAT) );
  XNOR2_X1 U518 ( .A(KEYINPUT118), .B(n533), .ZN(n458) );
  NAND2_X1 U519 ( .A1(n458), .A2(n457), .ZN(n461) );
  INV_X1 U520 ( .A(KEYINPUT54), .ZN(n459) );
  NOR2_X1 U521 ( .A1(n531), .A2(n462), .ZN(n576) );
  NAND2_X1 U522 ( .A1(n576), .A2(n479), .ZN(n464) );
  XOR2_X1 U523 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n463) );
  XNOR2_X1 U524 ( .A(n464), .B(n463), .ZN(n465) );
  AND2_X1 U525 ( .A1(n572), .A2(n560), .ZN(n469) );
  XNOR2_X1 U526 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n467) );
  INV_X1 U527 ( .A(G190GAT), .ZN(n466) );
  XNOR2_X1 U528 ( .A(G1GAT), .B(KEYINPUT95), .ZN(n470) );
  XNOR2_X1 U529 ( .A(n470), .B(KEYINPUT34), .ZN(n471) );
  XOR2_X1 U530 ( .A(KEYINPUT94), .B(n471), .Z(n495) );
  NAND2_X1 U531 ( .A1(n582), .A2(n563), .ZN(n506) );
  XOR2_X1 U532 ( .A(KEYINPUT82), .B(n472), .Z(n473) );
  NOR2_X1 U533 ( .A1(n483), .A2(n473), .ZN(n475) );
  NAND2_X1 U534 ( .A1(n475), .A2(n474), .ZN(n476) );
  NAND2_X1 U535 ( .A1(n531), .A2(n476), .ZN(n488) );
  NAND2_X1 U536 ( .A1(n535), .A2(n533), .ZN(n477) );
  NAND2_X1 U537 ( .A1(n479), .A2(n477), .ZN(n478) );
  XOR2_X1 U538 ( .A(KEYINPUT25), .B(n478), .Z(n486) );
  NOR2_X1 U539 ( .A1(n479), .A2(n535), .ZN(n482) );
  XOR2_X1 U540 ( .A(KEYINPUT92), .B(KEYINPUT26), .Z(n480) );
  XNOR2_X1 U541 ( .A(KEYINPUT91), .B(n480), .ZN(n481) );
  XOR2_X1 U542 ( .A(n482), .B(n481), .Z(n550) );
  NOR2_X1 U543 ( .A1(n483), .A2(n550), .ZN(n484) );
  NOR2_X1 U544 ( .A1(n531), .A2(n484), .ZN(n485) );
  NAND2_X1 U545 ( .A1(n486), .A2(n485), .ZN(n487) );
  NAND2_X1 U546 ( .A1(n488), .A2(n487), .ZN(n489) );
  XNOR2_X1 U547 ( .A(KEYINPUT93), .B(n489), .ZN(n502) );
  XOR2_X1 U548 ( .A(KEYINPUT78), .B(KEYINPUT16), .Z(n492) );
  NAND2_X1 U549 ( .A1(n558), .A2(n490), .ZN(n491) );
  XNOR2_X1 U550 ( .A(n492), .B(n491), .ZN(n493) );
  NAND2_X1 U551 ( .A1(n502), .A2(n493), .ZN(n520) );
  NOR2_X1 U552 ( .A1(n506), .A2(n520), .ZN(n500) );
  NAND2_X1 U553 ( .A1(n500), .A2(n531), .ZN(n494) );
  XNOR2_X1 U554 ( .A(n495), .B(n494), .ZN(G1324GAT) );
  NAND2_X1 U555 ( .A1(n500), .A2(n533), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n496), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT96), .B(KEYINPUT35), .Z(n498) );
  NAND2_X1 U558 ( .A1(n500), .A2(n535), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U560 ( .A(G15GAT), .B(n499), .ZN(G1326GAT) );
  NAND2_X1 U561 ( .A1(n500), .A2(n537), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n501), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U563 ( .A(KEYINPUT97), .B(KEYINPUT39), .Z(n509) );
  AND2_X1 U564 ( .A1(n585), .A2(n502), .ZN(n503) );
  XOR2_X1 U565 ( .A(KEYINPUT98), .B(n503), .Z(n504) );
  NOR2_X1 U566 ( .A1(n588), .A2(n504), .ZN(n505) );
  XNOR2_X1 U567 ( .A(KEYINPUT37), .B(n505), .ZN(n530) );
  NOR2_X1 U568 ( .A1(n530), .A2(n506), .ZN(n507) );
  XNOR2_X1 U569 ( .A(KEYINPUT38), .B(n507), .ZN(n518) );
  NAND2_X1 U570 ( .A1(n518), .A2(n531), .ZN(n508) );
  XNOR2_X1 U571 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U572 ( .A(G29GAT), .B(n510), .Z(G1328GAT) );
  XOR2_X1 U573 ( .A(G36GAT), .B(KEYINPUT99), .Z(n512) );
  NAND2_X1 U574 ( .A1(n533), .A2(n518), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n512), .B(n511), .ZN(G1329GAT) );
  XOR2_X1 U576 ( .A(KEYINPUT40), .B(KEYINPUT102), .Z(n514) );
  XNOR2_X1 U577 ( .A(G43GAT), .B(KEYINPUT101), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n514), .B(n513), .ZN(n517) );
  NAND2_X1 U579 ( .A1(n518), .A2(n535), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n515), .B(KEYINPUT100), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n517), .B(n516), .ZN(G1330GAT) );
  NAND2_X1 U582 ( .A1(n537), .A2(n518), .ZN(n519) );
  XNOR2_X1 U583 ( .A(G50GAT), .B(n519), .ZN(G1331GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT103), .B(KEYINPUT42), .Z(n522) );
  NAND2_X1 U585 ( .A1(n568), .A2(n577), .ZN(n529) );
  NOR2_X1 U586 ( .A1(n529), .A2(n520), .ZN(n526) );
  NAND2_X1 U587 ( .A1(n526), .A2(n531), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U589 ( .A(G57GAT), .B(n523), .ZN(G1332GAT) );
  NAND2_X1 U590 ( .A1(n526), .A2(n533), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n524), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U592 ( .A1(n526), .A2(n535), .ZN(n525) );
  XNOR2_X1 U593 ( .A(n525), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U594 ( .A(G78GAT), .B(KEYINPUT43), .Z(n528) );
  NAND2_X1 U595 ( .A1(n526), .A2(n537), .ZN(n527) );
  XNOR2_X1 U596 ( .A(n528), .B(n527), .ZN(G1335GAT) );
  NOR2_X1 U597 ( .A1(n530), .A2(n529), .ZN(n538) );
  NAND2_X1 U598 ( .A1(n538), .A2(n531), .ZN(n532) );
  XNOR2_X1 U599 ( .A(G85GAT), .B(n532), .ZN(G1336GAT) );
  NAND2_X1 U600 ( .A1(n538), .A2(n533), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n534), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U602 ( .A1(n538), .A2(n535), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n536), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT44), .B(KEYINPUT104), .Z(n540) );
  NAND2_X1 U605 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U607 ( .A(G106GAT), .B(n541), .Z(G1339GAT) );
  XOR2_X1 U608 ( .A(G113GAT), .B(KEYINPUT113), .Z(n543) );
  NAND2_X1 U609 ( .A1(n546), .A2(n563), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(G1340GAT) );
  NAND2_X1 U611 ( .A1(n546), .A2(n571), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n544), .B(KEYINPUT50), .ZN(n545) );
  XNOR2_X1 U613 ( .A(G127GAT), .B(n545), .ZN(G1342GAT) );
  NAND2_X1 U614 ( .A1(n560), .A2(n546), .ZN(n548) );
  XOR2_X1 U615 ( .A(KEYINPUT51), .B(KEYINPUT116), .Z(n547) );
  XNOR2_X1 U616 ( .A(G134GAT), .B(n549), .ZN(G1343GAT) );
  INV_X1 U617 ( .A(n550), .ZN(n575) );
  NAND2_X1 U618 ( .A1(n575), .A2(n551), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n552), .B(KEYINPUT117), .ZN(n561) );
  NAND2_X1 U620 ( .A1(n561), .A2(n553), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n556) );
  NAND2_X1 U623 ( .A1(n561), .A2(n568), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U625 ( .A(G148GAT), .B(n557), .ZN(G1345GAT) );
  NAND2_X1 U626 ( .A1(n561), .A2(n558), .ZN(n559) );
  XNOR2_X1 U627 ( .A(G155GAT), .B(n559), .ZN(G1346GAT) );
  NAND2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U630 ( .A1(n572), .A2(n563), .ZN(n564) );
  XNOR2_X1 U631 ( .A(G169GAT), .B(n564), .ZN(G1348GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n566) );
  XNOR2_X1 U633 ( .A(G176GAT), .B(KEYINPUT121), .ZN(n565) );
  XNOR2_X1 U634 ( .A(n566), .B(n565), .ZN(n567) );
  XOR2_X1 U635 ( .A(KEYINPUT56), .B(n567), .Z(n570) );
  NAND2_X1 U636 ( .A1(n572), .A2(n568), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(G1349GAT) );
  XOR2_X1 U638 ( .A(G183GAT), .B(KEYINPUT123), .Z(n574) );
  NAND2_X1 U639 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1350GAT) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n587) );
  NOR2_X1 U642 ( .A1(n587), .A2(n577), .ZN(n581) );
  XOR2_X1 U643 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n579) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  NOR2_X1 U647 ( .A1(n582), .A2(n587), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  NOR2_X1 U650 ( .A1(n585), .A2(n587), .ZN(n586) );
  XOR2_X1 U651 ( .A(G211GAT), .B(n586), .Z(G1354GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n590) );
  XNOR2_X1 U653 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n590), .B(n589), .ZN(n591) );
  XOR2_X1 U655 ( .A(G218GAT), .B(n591), .Z(G1355GAT) );
endmodule

