//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 1 0 0 0 0 1 0 0 1 1 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0 0 0 1 0 0 0 0 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:55 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1290, new_n1291,
    new_n1292, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT0), .Z(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n202), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n211), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT64), .Z(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n208), .B1(new_n219), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  OR2_X1    g0025(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n217), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT65), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n231), .B(new_n232), .Z(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G87), .B(G97), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  AND2_X1   g0044(.A1(KEYINPUT8), .A2(G58), .ZN(new_n245));
  NOR2_X1   g0045(.A1(KEYINPUT8), .A2(G58), .ZN(new_n246));
  NOR2_X1   g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NOR2_X1   g0047(.A1(G20), .A2(G33), .ZN(new_n248));
  AOI22_X1  g0048(.A1(new_n247), .A2(new_n248), .B1(G20), .B2(G77), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n213), .A2(G33), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT15), .B(G87), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  AND3_X1   g0053(.A1(new_n253), .A2(KEYINPUT69), .A3(new_n212), .ZN(new_n254));
  AOI21_X1  g0054(.A(KEYINPUT69), .B1(new_n253), .B2(new_n212), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G77), .ZN(new_n257));
  INV_X1    g0057(.A(G13), .ZN(new_n258));
  NOR3_X1   g0058(.A1(new_n258), .A2(new_n213), .A3(G1), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n252), .A2(new_n256), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n253), .A2(new_n212), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT69), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n253), .A2(KEYINPUT69), .A3(new_n212), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n259), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(KEYINPUT72), .B1(new_n213), .B2(G1), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT72), .ZN(new_n267));
  INV_X1    g0067(.A(G1), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(new_n268), .A3(G20), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n265), .A2(G77), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n260), .A2(new_n271), .ZN(new_n272));
  AND2_X1   g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NOR2_X1   g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  OAI21_X1  g0074(.A(KEYINPUT66), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT3), .ZN(new_n276));
  INV_X1    g0076(.A(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT66), .ZN(new_n279));
  NAND2_X1  g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G238), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G1698), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n284), .B1(G232), .B2(G1698), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  AND2_X1   g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  NOR3_X1   g0087(.A1(new_n287), .A2(KEYINPUT67), .A3(new_n212), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT67), .ZN(new_n289));
  AND2_X1   g0089(.A1(G1), .A2(G13), .ZN(new_n290));
  NAND2_X1  g0090(.A1(G33), .A2(G41), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n286), .B(new_n293), .C1(G107), .C2(new_n282), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n290), .A2(new_n291), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n268), .B1(G41), .B2(G45), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G41), .ZN(new_n299));
  INV_X1    g0099(.A(G45), .ZN(new_n300));
  AOI21_X1  g0100(.A(G1), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G274), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n302), .B1(new_n290), .B2(new_n291), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n298), .A2(G244), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n294), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n272), .B1(G200), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G190), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n306), .B1(new_n307), .B2(new_n305), .ZN(new_n308));
  INV_X1    g0108(.A(G169), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n310), .B(new_n272), .C1(G179), .C2(new_n305), .ZN(new_n311));
  AND2_X1   g0111(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  XOR2_X1   g0112(.A(new_n312), .B(KEYINPUT73), .Z(new_n313));
  OAI21_X1  g0113(.A(KEYINPUT67), .B1(new_n287), .B2(new_n212), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n290), .A2(new_n289), .A3(new_n291), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(G33), .A2(G87), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n278), .A2(new_n280), .ZN(new_n318));
  OR2_X1    g0118(.A1(G223), .A2(G1698), .ZN(new_n319));
  INV_X1    g0119(.A(G226), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G1698), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n318), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n316), .B1(new_n317), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n303), .A2(new_n301), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n295), .A2(G232), .A3(new_n296), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(KEYINPUT79), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G200), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n319), .A2(new_n321), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n273), .A2(new_n274), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n317), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n293), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT79), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n332), .A2(new_n333), .A3(new_n324), .A4(new_n325), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n327), .A2(new_n328), .A3(new_n334), .ZN(new_n335));
  AND2_X1   g0135(.A1(KEYINPUT80), .A2(G190), .ZN(new_n336));
  NOR2_X1   g0136(.A1(KEYINPUT80), .A2(G190), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n339), .B1(new_n331), .B2(new_n293), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT78), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n326), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n324), .A2(new_n325), .A3(KEYINPUT78), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n340), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT81), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT81), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n340), .A2(new_n342), .A3(new_n346), .A4(new_n343), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n335), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n278), .A2(KEYINPUT7), .A3(new_n213), .A4(new_n280), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT76), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n330), .A2(KEYINPUT76), .A3(KEYINPUT7), .A4(new_n213), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n278), .A2(new_n213), .A3(new_n280), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT7), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n351), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(G68), .ZN(new_n357));
  INV_X1    g0157(.A(G58), .ZN(new_n358));
  INV_X1    g0158(.A(G68), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(G20), .B1(new_n360), .B2(new_n201), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n248), .A2(G159), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n357), .A2(KEYINPUT16), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(G20), .B1(new_n275), .B2(new_n281), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n349), .B1(new_n366), .B2(KEYINPUT7), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n363), .B1(new_n367), .B2(G68), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n365), .B(new_n256), .C1(new_n368), .C2(KEYINPUT16), .ZN(new_n369));
  OR2_X1    g0169(.A1(KEYINPUT8), .A2(G58), .ZN(new_n370));
  NAND2_X1  g0170(.A1(KEYINPUT8), .A2(G58), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(KEYINPUT70), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT70), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(new_n245), .B2(new_n246), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n259), .ZN(new_n376));
  INV_X1    g0176(.A(new_n259), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n254), .B2(new_n255), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n270), .A2(new_n372), .A3(new_n374), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n376), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT77), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT77), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n376), .B(new_n382), .C1(new_n378), .C2(new_n379), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n348), .A2(new_n369), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT17), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n349), .ZN(new_n389));
  NOR3_X1   g0189(.A1(new_n273), .A2(new_n274), .A3(KEYINPUT66), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n279), .B1(new_n278), .B2(new_n280), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n213), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n389), .B1(new_n392), .B2(new_n354), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n364), .B1(new_n393), .B2(new_n359), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT16), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n256), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n363), .B1(new_n356), .B2(G68), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n397), .B1(new_n398), .B2(KEYINPUT16), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n384), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n342), .A2(new_n343), .ZN(new_n401));
  INV_X1    g0201(.A(G179), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n332), .A2(new_n402), .ZN(new_n403));
  OR2_X1    g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n327), .A2(new_n309), .A3(new_n334), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(KEYINPUT18), .B1(new_n400), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n369), .A2(new_n385), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT18), .ZN(new_n409));
  AND2_X1   g0209(.A1(new_n404), .A2(new_n405), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n400), .A2(KEYINPUT17), .A3(new_n348), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n388), .A2(new_n407), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n313), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(G1698), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n282), .A2(G222), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n282), .A2(G223), .A3(G1698), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n416), .B(new_n417), .C1(new_n257), .C2(new_n282), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n293), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n324), .B1(new_n297), .B2(new_n320), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT68), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n419), .A2(KEYINPUT68), .A3(new_n421), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NOR3_X1   g0224(.A1(new_n422), .A2(new_n424), .A3(G169), .ZN(new_n425));
  INV_X1    g0225(.A(new_n422), .ZN(new_n426));
  AOI21_X1  g0226(.A(G179), .B1(new_n426), .B2(new_n423), .ZN(new_n427));
  INV_X1    g0227(.A(G150), .ZN(new_n428));
  INV_X1    g0228(.A(new_n248), .ZN(new_n429));
  OAI22_X1  g0229(.A1(new_n375), .A2(new_n250), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n430), .A2(KEYINPUT71), .ZN(new_n431));
  OAI21_X1  g0231(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(new_n430), .B2(KEYINPUT71), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n256), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(G50), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n435), .B1(new_n266), .B2(new_n269), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n265), .A2(new_n436), .B1(new_n435), .B2(new_n259), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NOR3_X1   g0239(.A1(new_n425), .A2(new_n427), .A3(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(G190), .B1(new_n424), .B2(new_n422), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n426), .A2(G200), .A3(new_n423), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT9), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n438), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n439), .A2(KEYINPUT9), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n441), .A2(new_n442), .A3(new_n444), .A4(new_n445), .ZN(new_n446));
  OR2_X1    g0246(.A1(new_n446), .A2(KEYINPUT10), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(KEYINPUT10), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n440), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n248), .A2(G50), .B1(G20), .B2(new_n359), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(new_n257), .B2(new_n250), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n256), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT11), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n259), .A2(new_n359), .ZN(new_n455));
  XNOR2_X1  g0255(.A(new_n455), .B(KEYINPUT12), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n265), .A2(G68), .A3(new_n270), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n256), .A2(new_n451), .A3(KEYINPUT11), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n454), .A2(new_n456), .A3(new_n457), .A4(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT14), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT13), .ZN(new_n462));
  NOR2_X1   g0262(.A1(G226), .A2(G1698), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n463), .B1(new_n230), .B2(G1698), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n275), .A2(new_n464), .A3(new_n281), .ZN(new_n465));
  NAND2_X1  g0265(.A1(G33), .A2(G97), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT74), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT74), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n468), .A2(G33), .A3(G97), .ZN(new_n469));
  AND2_X1   g0269(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n293), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n324), .B1(new_n297), .B2(new_n283), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n462), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n316), .B1(new_n465), .B2(new_n470), .ZN(new_n476));
  NOR3_X1   g0276(.A1(new_n476), .A2(KEYINPUT13), .A3(new_n473), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n461), .B(G169), .C1(new_n475), .C2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n472), .A2(new_n462), .A3(new_n474), .ZN(new_n479));
  OAI21_X1  g0279(.A(KEYINPUT13), .B1(new_n476), .B2(new_n473), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n479), .A2(G179), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n479), .A2(new_n480), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n461), .B1(new_n483), .B2(G169), .ZN(new_n484));
  OAI21_X1  g0284(.A(KEYINPUT75), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(G169), .B1(new_n475), .B2(new_n477), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT14), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT75), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n487), .A2(new_n488), .A3(new_n481), .A4(new_n478), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n460), .B1(new_n485), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n483), .A2(G200), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n479), .A2(G190), .A3(new_n480), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n491), .A2(new_n460), .A3(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n414), .A2(new_n449), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n268), .A2(G33), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n265), .A2(KEYINPUT82), .A3(new_n498), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n377), .B(new_n498), .C1(new_n254), .C2(new_n255), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT82), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n499), .A2(new_n502), .A3(G97), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n259), .A2(new_n204), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n248), .A2(G77), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT6), .ZN(new_n506));
  NOR3_X1   g0306(.A1(new_n506), .A2(new_n204), .A3(G107), .ZN(new_n507));
  XNOR2_X1  g0307(.A(G97), .B(G107), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n507), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n505), .B1(new_n509), .B2(new_n213), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n510), .B1(new_n367), .B2(G107), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n503), .B(new_n504), .C1(new_n511), .C2(new_n397), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n300), .A2(G1), .ZN(new_n514));
  AND2_X1   g0314(.A1(KEYINPUT5), .A2(G41), .ZN(new_n515));
  NOR2_X1   g0315(.A1(KEYINPUT5), .A2(G41), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n517), .A2(G257), .A3(new_n295), .ZN(new_n518));
  XNOR2_X1  g0318(.A(KEYINPUT5), .B(G41), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n303), .A2(new_n514), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(G244), .B(new_n415), .C1(new_n273), .C2(new_n274), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT4), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n522), .A2(new_n523), .B1(G33), .B2(G283), .ZN(new_n524));
  INV_X1    g0324(.A(G244), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n275), .A2(new_n281), .A3(new_n415), .A4(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n275), .A2(new_n281), .A3(G250), .A4(G1698), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n524), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n521), .B1(new_n529), .B2(new_n293), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n307), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n531), .B1(G200), .B2(new_n530), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n513), .A2(new_n532), .ZN(new_n533));
  AOI211_X1 g0333(.A(G179), .B(new_n521), .C1(new_n529), .C2(new_n293), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n529), .A2(new_n293), .ZN(new_n536));
  INV_X1    g0336(.A(new_n521), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n309), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n512), .A2(new_n535), .A3(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(G87), .ZN(new_n541));
  NOR3_X1   g0341(.A1(new_n541), .A2(KEYINPUT22), .A3(G20), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n275), .A2(new_n281), .A3(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n213), .B(G87), .C1(new_n273), .C2(new_n274), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(KEYINPUT22), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NOR3_X1   g0346(.A1(new_n213), .A2(KEYINPUT23), .A3(G107), .ZN(new_n547));
  AOI21_X1  g0347(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n548));
  OAI22_X1  g0348(.A1(new_n547), .A2(KEYINPUT86), .B1(G20), .B2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT23), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n550), .A2(new_n205), .A3(G20), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT86), .ZN(new_n552));
  OAI22_X1  g0352(.A1(new_n551), .A2(new_n552), .B1(new_n550), .B2(new_n205), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  XOR2_X1   g0354(.A(KEYINPUT87), .B(KEYINPUT24), .Z(new_n555));
  AND3_X1   g0355(.A1(new_n546), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  OR2_X1    g0356(.A1(KEYINPUT87), .A2(KEYINPUT24), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n557), .B1(new_n546), .B2(new_n554), .ZN(new_n558));
  OR3_X1    g0358(.A1(new_n556), .A2(new_n558), .A3(new_n397), .ZN(new_n559));
  INV_X1    g0359(.A(G257), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(G1698), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n561), .B1(G250), .B2(G1698), .ZN(new_n562));
  INV_X1    g0362(.A(G294), .ZN(new_n563));
  OAI22_X1  g0363(.A1(new_n562), .A2(new_n330), .B1(new_n277), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n287), .A2(new_n212), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n514), .B2(new_n519), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n293), .A2(new_n564), .B1(new_n566), .B2(G264), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n567), .A2(KEYINPUT88), .A3(new_n307), .A4(new_n520), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT88), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n517), .A2(G264), .A3(new_n295), .ZN(new_n570));
  NOR2_X1   g0370(.A1(G250), .A2(G1698), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n571), .B1(new_n560), .B2(G1698), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n572), .A2(new_n318), .B1(G33), .B2(G294), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n520), .B(new_n570), .C1(new_n573), .C2(new_n316), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n569), .B1(new_n574), .B2(new_n328), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n574), .A2(G190), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n568), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n499), .A2(new_n502), .A3(G107), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n259), .A2(new_n205), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT25), .ZN(new_n580));
  XNOR2_X1  g0380(.A(new_n579), .B(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n559), .A2(new_n577), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n574), .A2(new_n309), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n564), .A2(new_n293), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n586), .A2(new_n402), .A3(new_n520), .A4(new_n570), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NOR3_X1   g0388(.A1(new_n556), .A2(new_n558), .A3(new_n397), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n588), .B1(new_n589), .B2(new_n582), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n533), .A2(new_n540), .A3(new_n584), .A4(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(G33), .A2(G283), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n592), .B(new_n213), .C1(G33), .C2(new_n204), .ZN(new_n593));
  INV_X1    g0393(.A(G116), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G20), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n593), .A2(new_n261), .A3(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT20), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n593), .A2(new_n261), .A3(KEYINPUT20), .A4(new_n595), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n258), .A2(G1), .ZN(new_n600));
  INV_X1    g0400(.A(new_n595), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n598), .A2(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n265), .A2(G116), .A3(new_n498), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT85), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n560), .A2(new_n415), .ZN(new_n606));
  INV_X1    g0406(.A(G264), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(G1698), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n606), .B(new_n608), .C1(new_n273), .C2(new_n274), .ZN(new_n609));
  INV_X1    g0409(.A(G303), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n605), .B(new_n609), .C1(new_n282), .C2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n610), .B1(new_n275), .B2(new_n281), .ZN(new_n612));
  INV_X1    g0412(.A(new_n609), .ZN(new_n613));
  OAI21_X1  g0413(.A(KEYINPUT85), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n611), .A2(new_n293), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n520), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(G270), .B2(new_n566), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n615), .A2(new_n339), .A3(new_n617), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n615), .A2(new_n617), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n604), .B(new_n618), .C1(new_n619), .C2(new_n328), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n604), .A2(new_n402), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n619), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT21), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n615), .A2(new_n617), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n309), .B1(new_n602), .B2(new_n603), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n624), .A2(new_n623), .A3(new_n625), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n620), .B(new_n622), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n251), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n629), .A2(new_n377), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT19), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n467), .B2(new_n469), .ZN(new_n632));
  OAI22_X1  g0432(.A1(new_n632), .A2(G20), .B1(G87), .B2(new_n206), .ZN(new_n633));
  AOI21_X1  g0433(.A(G20), .B1(new_n278), .B2(new_n280), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n213), .A2(G33), .A3(G97), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n634), .A2(G68), .B1(new_n635), .B2(new_n631), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n630), .B1(new_n637), .B2(new_n256), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n499), .A2(new_n502), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n638), .B1(new_n639), .B2(new_n251), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT84), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n638), .B(KEYINPUT84), .C1(new_n639), .C2(new_n251), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n303), .A2(new_n514), .ZN(new_n644));
  NOR2_X1   g0444(.A1(G238), .A2(G1698), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n645), .B1(new_n525), .B2(G1698), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n646), .A2(new_n318), .B1(G33), .B2(G116), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n644), .B1(new_n647), .B2(new_n316), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT83), .ZN(new_n649));
  OAI21_X1  g0449(.A(G250), .B1(new_n300), .B2(G1), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n649), .B1(new_n565), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n268), .A2(G45), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n295), .A2(KEYINPUT83), .A3(G250), .A4(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(G169), .B1(new_n648), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n525), .A2(G1698), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(G238), .B2(G1698), .ZN(new_n658));
  OAI22_X1  g0458(.A1(new_n658), .A2(new_n330), .B1(new_n277), .B2(new_n594), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(new_n293), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n660), .A2(G179), .A3(new_n654), .A4(new_n644), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n642), .A2(new_n643), .A3(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n499), .A2(new_n502), .A3(G87), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n638), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n648), .A2(new_n655), .A3(new_n307), .ZN(new_n667));
  AOI22_X1  g0467(.A1(new_n659), .A2(new_n293), .B1(new_n303), .B2(new_n514), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n328), .B1(new_n668), .B2(new_n654), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n663), .A2(new_n671), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n591), .A2(new_n628), .A3(new_n672), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n497), .A2(new_n673), .ZN(G372));
  NAND2_X1  g0474(.A1(new_n447), .A2(new_n448), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n388), .A2(new_n412), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n494), .A2(new_n311), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n676), .B1(new_n490), .B2(new_n677), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n407), .A2(new_n411), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n440), .B1(new_n675), .B2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT91), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n540), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n640), .A2(new_n662), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT89), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n638), .A2(new_n664), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n685), .B1(new_n638), .B2(new_n664), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n670), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n512), .A2(new_n539), .A3(KEYINPUT91), .A4(new_n535), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n683), .A2(new_n684), .A3(new_n688), .A4(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT26), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT92), .ZN(new_n693));
  AOI22_X1  g0493(.A1(new_n640), .A2(new_n641), .B1(new_n656), .B2(new_n661), .ZN(new_n694));
  AOI22_X1  g0494(.A1(new_n694), .A2(new_n643), .B1(new_n666), .B2(new_n670), .ZN(new_n695));
  INV_X1    g0495(.A(new_n540), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(KEYINPUT26), .A3(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n692), .A2(new_n693), .A3(new_n697), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n695), .A2(KEYINPUT92), .A3(KEYINPUT26), .A4(new_n696), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n699), .A2(new_n684), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n533), .A2(new_n540), .A3(new_n584), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n688), .A2(new_n684), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n622), .B(new_n590), .C1(new_n627), .C2(new_n626), .ZN(new_n704));
  AOI21_X1  g0504(.A(KEYINPUT90), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n704), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT90), .ZN(new_n707));
  NOR4_X1   g0507(.A1(new_n706), .A2(new_n701), .A3(new_n707), .A4(new_n702), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n698), .B(new_n700), .C1(new_n705), .C2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n681), .B1(new_n496), .B2(new_n710), .ZN(G369));
  OAI21_X1  g0511(.A(new_n622), .B1(new_n627), .B2(new_n626), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n600), .A2(new_n213), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n713), .A2(KEYINPUT27), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(KEYINPUT27), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n714), .A2(G213), .A3(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(G343), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n604), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n712), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(new_n628), .B2(new_n720), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n722), .A2(G330), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n718), .B1(new_n589), .B2(new_n582), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n584), .A2(new_n590), .A3(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n725), .B1(new_n590), .B2(new_n719), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n712), .A2(new_n719), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(new_n725), .ZN(new_n729));
  INV_X1    g0529(.A(new_n590), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n729), .B1(new_n730), .B2(new_n719), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n727), .A2(new_n731), .ZN(G399));
  INV_X1    g0532(.A(new_n209), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(G41), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n735), .A2(G1), .A3(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(new_n215), .B2(new_n735), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n738), .B(KEYINPUT28), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n709), .A2(new_n719), .ZN(new_n740));
  XNOR2_X1  g0540(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n665), .A2(KEYINPUT89), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n638), .A2(new_n664), .A3(new_n685), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AOI22_X1  g0545(.A1(new_n745), .A2(new_n670), .B1(new_n640), .B2(new_n662), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n746), .A2(new_n540), .A3(new_n533), .A4(new_n584), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n684), .B1(new_n747), .B2(new_n706), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n690), .A2(KEYINPUT26), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n695), .A2(new_n691), .A3(new_n696), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OAI211_X1 g0551(.A(KEYINPUT29), .B(new_n719), .C1(new_n748), .C2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n742), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n591), .ZN(new_n754));
  INV_X1    g0554(.A(new_n620), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n712), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n754), .A2(new_n756), .A3(new_n695), .A4(new_n719), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n586), .A2(new_n570), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n661), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n759), .A2(new_n615), .A3(new_n617), .A4(new_n530), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT30), .ZN(new_n761));
  OAI211_X1 g0561(.A(new_n574), .B(new_n402), .C1(new_n648), .C2(new_n655), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n530), .ZN(new_n763));
  AOI22_X1  g0563(.A1(new_n760), .A2(new_n761), .B1(new_n763), .B2(new_n624), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT93), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n765), .B1(new_n760), .B2(new_n761), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n567), .A2(G179), .A3(new_n668), .A4(new_n654), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n538), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n768), .A2(new_n619), .A3(KEYINPUT93), .A4(KEYINPUT30), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n764), .A2(new_n766), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(new_n718), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT31), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n770), .A2(KEYINPUT31), .A3(new_n718), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n757), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G330), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n753), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n739), .B1(new_n778), .B2(G1), .ZN(G364));
  NOR2_X1   g0579(.A1(new_n722), .A2(G330), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n258), .A2(G20), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n268), .B1(new_n781), .B2(G45), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n734), .A2(new_n783), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n723), .A2(new_n780), .A3(new_n784), .ZN(new_n785));
  XOR2_X1   g0585(.A(new_n785), .B(KEYINPUT95), .Z(new_n786));
  XNOR2_X1  g0586(.A(new_n784), .B(KEYINPUT96), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n733), .A2(new_n318), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n788), .B1(G45), .B2(new_n215), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n789), .B1(new_n243), .B2(G45), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n282), .A2(new_n209), .ZN(new_n791));
  INV_X1    g0591(.A(G355), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n791), .A2(new_n792), .B1(G116), .B2(new_n209), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(G13), .A2(G33), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(G20), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n212), .B1(G20), .B2(new_n309), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n799), .B(KEYINPUT97), .Z(new_n800));
  OAI21_X1  g0600(.A(new_n787), .B1(new_n794), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n797), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n722), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n338), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT98), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n805), .A2(new_n806), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G326), .ZN(new_n812));
  INV_X1    g0612(.A(new_n282), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n213), .A2(G179), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n814), .A2(G190), .A3(G200), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n813), .B1(new_n610), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n814), .A2(new_n307), .A3(new_n328), .ZN(new_n817));
  OR2_X1    g0617(.A1(new_n817), .A2(KEYINPUT101), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(KEYINPUT101), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n816), .B1(G329), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n804), .A2(G190), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  XNOR2_X1  g0624(.A(KEYINPUT33), .B(G317), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n824), .B1(KEYINPUT102), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(KEYINPUT102), .B2(new_n826), .ZN(new_n828));
  NOR3_X1   g0628(.A1(new_n213), .A2(new_n402), .A3(G200), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n339), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(G322), .ZN(new_n831));
  NOR3_X1   g0631(.A1(new_n307), .A2(G179), .A3(G200), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n832), .A2(new_n213), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n830), .A2(new_n831), .B1(new_n563), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n829), .A2(new_n307), .ZN(new_n835));
  INV_X1    g0635(.A(G311), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n814), .A2(new_n307), .A3(G200), .ZN(new_n837));
  INV_X1    g0637(.A(G283), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n835), .A2(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n834), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n812), .A2(new_n822), .A3(new_n828), .A4(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n815), .A2(new_n541), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n282), .B1(new_n205), .B2(new_n837), .ZN(new_n843));
  INV_X1    g0643(.A(new_n830), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n842), .B(new_n843), .C1(G58), .C2(new_n844), .ZN(new_n845));
  XOR2_X1   g0645(.A(KEYINPUT99), .B(G159), .Z(new_n846));
  NOR2_X1   g0646(.A1(new_n846), .A2(new_n817), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT32), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n847), .A2(new_n848), .B1(new_n257), .B2(new_n835), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(new_n848), .B2(new_n847), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n845), .B(new_n850), .C1(new_n435), .C2(new_n810), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n833), .A2(new_n204), .B1(new_n824), .B2(new_n359), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT100), .Z(new_n853));
  OAI21_X1  g0653(.A(new_n841), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n801), .B(new_n803), .C1(new_n798), .C2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n786), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(G396));
  OR3_X1    g0657(.A1(new_n311), .A2(KEYINPUT104), .A3(new_n719), .ZN(new_n858));
  OAI21_X1  g0658(.A(KEYINPUT104), .B1(new_n311), .B2(new_n719), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n272), .A2(new_n718), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n312), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n740), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n709), .A2(new_n719), .A3(new_n863), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n784), .B1(new_n867), .B2(new_n776), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n776), .B2(new_n867), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n835), .A2(new_n594), .B1(new_n824), .B2(new_n838), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n811), .B2(G303), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n871), .B(KEYINPUT103), .ZN(new_n872));
  INV_X1    g0672(.A(new_n837), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n844), .A2(G294), .B1(G87), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n205), .B2(new_n815), .ZN(new_n875));
  OAI221_X1 g0675(.A(new_n813), .B1(new_n204), .B2(new_n833), .C1(new_n820), .C2(new_n836), .ZN(new_n876));
  NOR3_X1   g0676(.A1(new_n872), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n835), .ZN(new_n878));
  INV_X1    g0678(.A(new_n846), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n878), .A2(new_n879), .B1(new_n823), .B2(G150), .ZN(new_n880));
  INV_X1    g0680(.A(G143), .ZN(new_n881));
  INV_X1    g0681(.A(G137), .ZN(new_n882));
  OAI221_X1 g0682(.A(new_n880), .B1(new_n881), .B2(new_n830), .C1(new_n810), .C2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n884), .A2(KEYINPUT34), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n884), .A2(KEYINPUT34), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n837), .A2(new_n359), .ZN(new_n887));
  INV_X1    g0687(.A(new_n815), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n887), .B1(G50), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n833), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n330), .B1(new_n890), .B2(G58), .ZN(new_n891));
  INV_X1    g0691(.A(G132), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n889), .B(new_n891), .C1(new_n820), .C2(new_n892), .ZN(new_n893));
  NOR3_X1   g0693(.A1(new_n885), .A2(new_n886), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n798), .B1(new_n877), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n787), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n798), .A2(new_n795), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n896), .B1(new_n257), .B2(new_n897), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n895), .B(new_n898), .C1(new_n863), .C2(new_n796), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n869), .A2(new_n899), .ZN(G384));
  INV_X1    g0700(.A(G330), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT106), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n460), .A2(new_n719), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n903), .B(KEYINPUT105), .ZN(new_n904));
  NOR3_X1   g0704(.A1(new_n490), .A2(new_n494), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n485), .A2(new_n489), .A3(new_n493), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n906), .A2(new_n903), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n902), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n485), .A2(new_n489), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n459), .ZN(new_n910));
  INV_X1    g0710(.A(new_n904), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n910), .A2(new_n493), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n906), .A2(new_n903), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n912), .A2(KEYINPUT106), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n908), .A2(new_n914), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n335), .A2(new_n345), .A3(new_n347), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n357), .A2(new_n364), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n395), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n384), .B1(new_n918), .B2(new_n399), .ZN(new_n919));
  OAI22_X1  g0719(.A1(new_n408), .A2(new_n916), .B1(new_n919), .B2(new_n406), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n919), .A2(new_n716), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT37), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n408), .A2(new_n410), .ZN(new_n923));
  INV_X1    g0723(.A(new_n716), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n408), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT37), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n923), .A2(new_n925), .A3(new_n926), .A4(new_n386), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n922), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n413), .A2(new_n921), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT38), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n928), .A2(new_n929), .A3(KEYINPUT38), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT31), .B1(new_n770), .B2(new_n718), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(new_n673), .B2(new_n719), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n864), .B1(new_n936), .B2(new_n774), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n915), .A2(new_n934), .A3(new_n937), .ZN(new_n938));
  XOR2_X1   g0738(.A(KEYINPUT108), .B(KEYINPUT40), .Z(new_n939));
  NAND2_X1  g0739(.A1(new_n775), .A2(new_n863), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(new_n908), .B2(new_n914), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT40), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n923), .A2(new_n925), .A3(new_n386), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(new_n926), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n925), .B1(new_n676), .B2(new_n679), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n931), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n942), .B1(new_n946), .B2(new_n933), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n938), .A2(new_n939), .B1(new_n941), .B2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n497), .A2(new_n775), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n901), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT109), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n952), .A2(new_n953), .B1(new_n949), .B2(new_n950), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n953), .B2(new_n952), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n490), .A2(new_n719), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT107), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT39), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n946), .A2(new_n958), .A3(new_n959), .A4(new_n933), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n946), .A2(new_n959), .A3(new_n933), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(KEYINPUT107), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n959), .B1(new_n932), .B2(new_n933), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n957), .B(new_n960), .C1(new_n962), .C2(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n311), .A2(new_n718), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n866), .A2(new_n966), .B1(new_n908), .B2(new_n914), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n934), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n679), .A2(new_n924), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n964), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n497), .A2(new_n742), .A3(new_n752), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n971), .A2(new_n681), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n970), .B(new_n972), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n955), .A2(new_n973), .B1(new_n268), .B2(new_n781), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(new_n973), .B2(new_n955), .ZN(new_n975));
  INV_X1    g0775(.A(new_n509), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n976), .A2(KEYINPUT35), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(KEYINPUT35), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n977), .A2(G116), .A3(new_n214), .A4(new_n978), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT36), .Z(new_n980));
  OR3_X1    g0780(.A1(new_n215), .A2(new_n257), .A3(new_n360), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n435), .A2(G68), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n268), .B(G13), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  OR3_X1    g0783(.A1(new_n975), .A2(new_n980), .A3(new_n983), .ZN(G367));
  INV_X1    g0784(.A(new_n788), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n799), .B1(new_n209), .B2(new_n251), .C1(new_n236), .C2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n787), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n873), .A2(G77), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n358), .B2(new_n815), .ZN(new_n989));
  INV_X1    g0789(.A(new_n817), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n813), .B(new_n989), .C1(G137), .C2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n811), .A2(G143), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n878), .A2(G50), .B1(new_n879), .B2(new_n823), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n844), .A2(G150), .B1(G68), .B2(new_n890), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n991), .A2(new_n992), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n810), .A2(new_n836), .ZN(new_n996));
  XNOR2_X1  g0796(.A(KEYINPUT113), .B(G317), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n330), .B1(new_n817), .B2(new_n997), .C1(new_n830), .C2(new_n610), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n833), .A2(new_n205), .B1(new_n837), .B2(new_n204), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n835), .A2(new_n838), .B1(new_n824), .B2(new_n563), .ZN(new_n1000));
  OR4_X1    g0800(.A1(new_n996), .A2(new_n998), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(KEYINPUT112), .B1(new_n888), .B2(G116), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT46), .Z(new_n1003));
  OAI21_X1  g0803(.A(new_n995), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT47), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n987), .B1(new_n1005), .B2(new_n798), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n743), .A2(new_n744), .A3(new_n718), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n746), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n684), .B2(new_n1007), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1006), .B1(new_n1009), .B2(new_n802), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n727), .A2(KEYINPUT111), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n533), .B(new_n540), .C1(new_n513), .C2(new_n719), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n696), .A2(new_n718), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n731), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT45), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n731), .A2(KEYINPUT45), .A3(new_n1014), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1011), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n727), .A2(KEYINPUT111), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT44), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n1021), .A2(KEYINPUT110), .ZN(new_n1022));
  OR3_X1    g0822(.A1(new_n731), .A2(new_n1014), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1021), .A2(KEYINPUT110), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1022), .B1(new_n731), .B2(new_n1014), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1019), .A2(new_n1020), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1020), .B1(new_n1019), .B2(new_n1026), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n729), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n728), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1031), .B1(new_n726), .B2(new_n1032), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(new_n723), .Z(new_n1034));
  OAI21_X1  g0834(.A(new_n778), .B1(new_n1030), .B2(new_n1034), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n734), .B(KEYINPUT41), .Z(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n783), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n1012), .A2(new_n590), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n718), .B1(new_n1039), .B2(new_n540), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n729), .A2(new_n1014), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1040), .B1(new_n1041), .B2(KEYINPUT42), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1041), .A2(KEYINPUT42), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n1042), .A2(new_n1043), .B1(KEYINPUT43), .B2(new_n1009), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1009), .A2(KEYINPUT43), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1044), .B(new_n1045), .Z(new_n1046));
  INV_X1    g0846(.A(new_n1014), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n727), .A2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1046), .B(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1010), .B1(new_n1038), .B2(new_n1050), .ZN(G387));
  INV_X1    g0851(.A(new_n1034), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n783), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n791), .A2(new_n736), .B1(G107), .B2(new_n209), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n233), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT114), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n247), .A2(new_n435), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT50), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n736), .B(new_n300), .C1(new_n359), .C2(new_n257), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n788), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n1055), .A2(G45), .B1(new_n1056), .B2(new_n1060), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1060), .A2(new_n1056), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1054), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n787), .B1(new_n1063), .B2(new_n800), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n833), .A2(new_n251), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n835), .A2(new_n359), .B1(new_n815), .B2(new_n257), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1065), .B(new_n1066), .C1(G50), .C2(new_n844), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n318), .B1(new_n817), .B2(new_n428), .C1(new_n204), .C2(new_n837), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n375), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1068), .B1(new_n1069), .B2(new_n823), .ZN(new_n1070));
  INV_X1    g0870(.A(G159), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1067), .B(new_n1070), .C1(new_n1071), .C2(new_n810), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n830), .A2(new_n997), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(G311), .B2(new_n823), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1074), .B1(new_n610), .B2(new_n835), .C1(new_n810), .C2(new_n831), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT115), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT48), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n833), .A2(new_n838), .B1(new_n815), .B2(new_n563), .ZN(new_n1080));
  NOR3_X1   g0880(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(KEYINPUT49), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n318), .B1(new_n990), .B2(G326), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1082), .B(new_n1083), .C1(new_n594), .C2(new_n837), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1081), .A2(KEYINPUT49), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1072), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1064), .B1(new_n1086), .B2(new_n798), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(KEYINPUT116), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n726), .B2(new_n802), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1087), .A2(KEYINPUT116), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n777), .A2(new_n1034), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n734), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n778), .A2(new_n1052), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n1053), .B1(new_n1089), .B2(new_n1090), .C1(new_n1093), .C2(new_n1094), .ZN(G393));
  INV_X1    g0895(.A(new_n1030), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n1091), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1030), .A2(new_n1092), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1097), .A2(new_n1098), .A3(new_n734), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1096), .A2(new_n783), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n240), .A2(new_n788), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1101), .B(new_n799), .C1(new_n204), .C2(new_n209), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n896), .B1(new_n1102), .B2(KEYINPUT117), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(KEYINPUT117), .B2(new_n1102), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n811), .A2(G317), .B1(G311), .B2(new_n844), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT52), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n282), .B1(G322), .B2(new_n990), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n890), .A2(G116), .B1(G303), .B2(new_n823), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n888), .A2(G283), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n878), .A2(G294), .B1(new_n873), .B2(G107), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n810), .A2(new_n428), .B1(new_n1071), .B2(new_n830), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1112), .B(KEYINPUT51), .Z(new_n1113));
  NOR2_X1   g0913(.A1(new_n833), .A2(new_n257), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(G50), .B2(new_n823), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n318), .B1(new_n817), .B2(new_n881), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(G87), .B2(new_n873), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n878), .A2(new_n247), .B1(new_n888), .B2(G68), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1115), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n1106), .A2(new_n1111), .B1(new_n1113), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1104), .B1(new_n1120), .B2(new_n798), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n802), .B2(new_n1014), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1099), .A2(new_n1100), .A3(new_n1122), .ZN(G390));
  OR2_X1    g0923(.A1(new_n496), .A2(new_n776), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n971), .A2(new_n1124), .A3(new_n681), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n915), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n901), .B2(new_n940), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n915), .A2(new_n937), .A3(G330), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n699), .A2(new_n684), .ZN(new_n1130));
  AOI21_X1  g0930(.A(KEYINPUT92), .B1(new_n690), .B2(new_n691), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1130), .B1(new_n697), .B2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n707), .B1(new_n747), .B2(new_n706), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n703), .A2(KEYINPUT90), .A3(new_n704), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n718), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n965), .B1(new_n1136), .B2(new_n863), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1129), .A2(new_n1138), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n719), .B(new_n863), .C1(new_n748), .C2(new_n751), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n1140), .A2(new_n966), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1127), .A2(new_n1128), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1125), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(KEYINPUT119), .B1(new_n967), .B2(new_n957), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n960), .B1(new_n962), .B2(new_n963), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT119), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1147), .B(new_n956), .C1(new_n1137), .C2(new_n1126), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1145), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n957), .B1(new_n946), .B2(new_n933), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n1141), .B2(new_n1126), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT118), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1150), .B(KEYINPUT118), .C1(new_n1141), .C2(new_n1126), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n1149), .A2(new_n1128), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1128), .B1(new_n1149), .B2(new_n1155), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1144), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1149), .A2(new_n1155), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1128), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1149), .A2(new_n1128), .A3(new_n1155), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1161), .A2(new_n1162), .A3(new_n1143), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1158), .A2(new_n1163), .A3(new_n734), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n783), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1146), .A2(new_n795), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n897), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n787), .B1(new_n1069), .B2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n282), .B1(new_n824), .B2(new_n882), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(KEYINPUT54), .B(G143), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n878), .A2(new_n1172), .B1(new_n873), .B2(G50), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1173), .B1(new_n892), .B2(new_n830), .C1(new_n1071), .C2(new_n833), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1170), .B(new_n1174), .C1(G125), .C2(new_n821), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n815), .A2(new_n428), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT53), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n811), .A2(G128), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1175), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n830), .A2(new_n594), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n835), .A2(new_n204), .B1(new_n824), .B2(new_n205), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1180), .B(new_n1181), .C1(new_n811), .C2(G283), .ZN(new_n1182));
  NOR4_X1   g0982(.A1(new_n282), .A2(new_n1114), .A3(new_n842), .A4(new_n887), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1182), .B(new_n1183), .C1(new_n563), .C2(new_n820), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1179), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1169), .B1(new_n1185), .B2(new_n798), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1167), .A2(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1187), .B(KEYINPUT120), .ZN(new_n1188));
  AND3_X1   g0988(.A1(new_n1166), .A2(KEYINPUT121), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(KEYINPUT121), .B1(new_n1166), .B2(new_n1188), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1164), .B1(new_n1189), .B2(new_n1190), .ZN(G378));
  NAND2_X1  g0991(.A1(new_n938), .A2(new_n939), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n947), .A2(new_n915), .A3(new_n937), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1192), .A2(KEYINPUT124), .A3(G330), .A4(new_n1193), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n439), .A2(new_n716), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  OR2_X1    g0997(.A1(new_n449), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n449), .A2(new_n1197), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1195), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n449), .A2(new_n1197), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n440), .B(new_n1196), .C1(new_n447), .C2(new_n448), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1195), .ZN(new_n1203));
  NOR3_X1   g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1200), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1194), .A2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(KEYINPUT124), .B1(new_n948), .B2(G330), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1192), .A2(G330), .A3(new_n1193), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT124), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1198), .A2(new_n1199), .A3(new_n1195), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1203), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  AND3_X1   g1013(.A1(new_n1209), .A2(new_n1210), .A3(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n970), .B1(new_n1208), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1216), .A2(new_n1194), .A3(new_n1205), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n970), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1215), .A2(new_n783), .A3(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n784), .B1(G50), .B2(new_n1168), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT123), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n318), .A2(G41), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1224), .B1(new_n358), .B2(new_n837), .C1(new_n257), .C2(new_n815), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n821), .B2(G283), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1226), .B(KEYINPUT122), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n835), .A2(new_n251), .B1(new_n833), .B2(new_n359), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n830), .A2(new_n205), .B1(new_n204), .B2(new_n824), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n1228), .B(new_n1229), .C1(new_n811), .C2(G116), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1227), .A2(new_n1230), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1231), .B(KEYINPUT58), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n435), .B1(G33), .B2(G41), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n824), .A2(new_n892), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n833), .A2(new_n428), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n1234), .B(new_n1235), .C1(new_n844), .C2(G128), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1236), .B1(new_n882), .B2(new_n835), .C1(new_n815), .C2(new_n1171), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(G125), .B2(new_n811), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(KEYINPUT59), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n879), .A2(new_n873), .ZN(new_n1241));
  AOI211_X1 g1041(.A(G33), .B(G41), .C1(new_n990), .C2(G124), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1240), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1239), .A2(KEYINPUT59), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n1232), .B1(new_n1224), .B2(new_n1233), .C1(new_n1243), .C2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1223), .B1(new_n1245), .B2(new_n798), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n1213), .B2(new_n796), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1221), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT57), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1125), .B1(new_n1165), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1215), .A2(new_n1220), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1250), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  AND3_X1   g1054(.A1(new_n1215), .A2(KEYINPUT57), .A3(new_n1220), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1125), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1163), .A2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n735), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT125), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1254), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  AOI211_X1 g1060(.A(KEYINPUT125), .B(new_n735), .C1(new_n1255), .C2(new_n1257), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1249), .B1(new_n1260), .B2(new_n1261), .ZN(G375));
  NAND3_X1  g1062(.A1(new_n1139), .A2(new_n1125), .A3(new_n1142), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1144), .A2(new_n1037), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1126), .A2(new_n795), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n787), .B1(G68), .B2(new_n1168), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n813), .A2(new_n988), .ZN(new_n1267));
  AOI211_X1 g1067(.A(new_n1065), .B(new_n1267), .C1(G97), .C2(new_n888), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n821), .A2(G303), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n811), .A2(G294), .ZN(new_n1270));
  OAI22_X1  g1070(.A1(new_n830), .A2(new_n838), .B1(new_n205), .B2(new_n835), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1271), .B1(G116), .B2(new_n823), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1268), .A2(new_n1269), .A3(new_n1270), .A4(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n811), .A2(G132), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n821), .A2(G128), .ZN(new_n1275));
  OAI22_X1  g1075(.A1(new_n835), .A2(new_n428), .B1(new_n815), .B2(new_n1071), .ZN(new_n1276));
  AOI211_X1 g1076(.A(new_n330), .B(new_n1276), .C1(G58), .C2(new_n873), .ZN(new_n1277));
  OAI22_X1  g1077(.A1(new_n833), .A2(new_n435), .B1(new_n824), .B2(new_n1171), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1278), .B1(G137), .B2(new_n844), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1274), .A2(new_n1275), .A3(new_n1277), .A4(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1273), .A2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1266), .B1(new_n1281), .B2(new_n798), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n1251), .A2(new_n783), .B1(new_n1265), .B2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1264), .A2(new_n1283), .ZN(G381));
  INV_X1    g1084(.A(G375), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1164), .A2(new_n1188), .A3(new_n1166), .ZN(new_n1286));
  OR4_X1    g1086(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1287));
  NOR3_X1   g1087(.A1(new_n1287), .A2(G387), .A3(G381), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1285), .A2(new_n1286), .A3(new_n1288), .ZN(G407));
  NAND2_X1  g1089(.A1(new_n717), .A2(G213), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1285), .A2(new_n1286), .A3(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(G407), .A2(new_n1292), .A3(G213), .ZN(G409));
  INV_X1    g1093(.A(KEYINPUT63), .ZN(new_n1294));
  OAI211_X1 g1094(.A(G378), .B(new_n1249), .C1(new_n1260), .C2(new_n1261), .ZN(new_n1295));
  NOR3_X1   g1095(.A1(new_n1252), .A2(new_n1036), .A3(new_n1253), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1286), .B1(new_n1296), .B2(new_n1248), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1290), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1144), .A2(KEYINPUT60), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1300), .A2(new_n1263), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n734), .B1(new_n1300), .B2(new_n1263), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n869), .A2(KEYINPUT126), .A3(new_n899), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1283), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT126), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(G384), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  NOR3_X1   g1108(.A1(new_n1303), .A2(new_n1305), .A3(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1308), .B1(new_n1303), .B2(new_n1305), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1294), .B1(new_n1299), .B2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1291), .A2(G2897), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1311), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1315), .B1(new_n1316), .B2(new_n1309), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1315), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1310), .A2(new_n1311), .A3(new_n1318), .ZN(new_n1319));
  AND2_X1   g1119(.A1(new_n1317), .A2(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(KEYINPUT61), .B1(new_n1299), .B2(new_n1320), .ZN(new_n1321));
  OR2_X1    g1121(.A1(new_n1038), .A2(new_n1050), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1322), .A2(new_n1010), .A3(G390), .ZN(new_n1323));
  INV_X1    g1123(.A(G390), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(G387), .ZN(new_n1325));
  XNOR2_X1  g1125(.A(G393), .B(new_n856), .ZN(new_n1326));
  AND3_X1   g1126(.A1(new_n1323), .A2(new_n1325), .A3(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1326), .B1(new_n1323), .B2(new_n1325), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1291), .B1(new_n1295), .B2(new_n1297), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1330), .A2(KEYINPUT63), .A3(new_n1312), .ZN(new_n1331));
  NAND4_X1  g1131(.A1(new_n1314), .A2(new_n1321), .A3(new_n1329), .A4(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT62), .ZN(new_n1333));
  AND3_X1   g1133(.A1(new_n1330), .A2(new_n1333), .A3(new_n1312), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT61), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1317), .A2(new_n1319), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1335), .B1(new_n1330), .B2(new_n1336), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1333), .B1(new_n1330), .B2(new_n1312), .ZN(new_n1338));
  NOR3_X1   g1138(.A1(new_n1334), .A2(new_n1337), .A3(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT127), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1340), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1326), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1324), .A2(G387), .ZN(new_n1343));
  AOI21_X1  g1143(.A(G390), .B1(new_n1322), .B2(new_n1010), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1342), .B1(new_n1343), .B2(new_n1344), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1323), .A2(new_n1325), .A3(new_n1326), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1345), .A2(KEYINPUT127), .A3(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1341), .A2(new_n1347), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1332), .B1(new_n1339), .B2(new_n1348), .ZN(G405));
  NAND2_X1  g1149(.A1(G375), .A2(new_n1286), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1350), .A2(new_n1295), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1351), .A2(new_n1347), .A3(new_n1341), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1348), .A2(new_n1295), .A3(new_n1350), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1352), .A2(new_n1353), .ZN(new_n1354));
  XNOR2_X1  g1154(.A(new_n1354), .B(new_n1312), .ZN(G402));
endmodule


