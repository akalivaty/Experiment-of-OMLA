//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 1 1 1 1 1 1 0 0 1 0 0 0 1 1 1 0 1 0 0 1 1 0 0 1 1 1 0 0 1 0 0 1 1 1 1 0 1 1 0 0 1 0 0 0 0 1 0 0 0 1 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1184, new_n1185, new_n1186, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n207));
  INV_X1    g0007(.A(G77), .ZN(new_n208));
  INV_X1    g0008(.A(G244), .ZN(new_n209));
  INV_X1    g0009(.A(G107), .ZN(new_n210));
  INV_X1    g0010(.A(G264), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G58), .ZN(new_n214));
  INV_X1    g0014(.A(G232), .ZN(new_n215));
  INV_X1    g0015(.A(G97), .ZN(new_n216));
  INV_X1    g0016(.A(G257), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n206), .B1(new_n212), .B2(new_n218), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT64), .Z(new_n220));
  INV_X1    g0020(.A(KEYINPUT1), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n220), .A2(new_n221), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n206), .A2(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT0), .Z(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n227), .A2(new_n204), .ZN(new_n228));
  OAI21_X1  g0028(.A(G50), .B1(G58), .B2(G68), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n226), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  AND3_X1   g0031(.A1(new_n222), .A2(new_n223), .A3(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(new_n215), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  AOI21_X1  g0047(.A(new_n227), .B1(G33), .B2(G41), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT3), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G33), .ZN(new_n252));
  AND2_X1   g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G1698), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n254), .B(KEYINPUT66), .ZN(new_n255));
  INV_X1    g0055(.A(G223), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n253), .A2(G222), .A3(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n259), .B1(new_n208), .B2(new_n253), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n248), .B1(new_n257), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G41), .ZN(new_n262));
  OAI21_X1  g0062(.A(KEYINPUT65), .B1(new_n249), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n227), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT65), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(G33), .A3(G41), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n263), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G45), .ZN(new_n268));
  AOI21_X1  g0068(.A(G1), .B1(new_n262), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n267), .A2(G274), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n269), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n267), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n271), .B1(G226), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n261), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT67), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT67), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n261), .A2(new_n278), .A3(new_n275), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G190), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n277), .A2(new_n279), .A3(G200), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G50), .A2(G58), .ZN(new_n283));
  INV_X1    g0083(.A(G68), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n204), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n204), .A2(G33), .ZN(new_n287));
  INV_X1    g0087(.A(G150), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G20), .A2(G33), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  OAI22_X1  g0090(.A1(new_n286), .A2(new_n287), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n285), .B1(new_n291), .B2(KEYINPUT68), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n292), .B1(KEYINPUT68), .B2(new_n291), .ZN(new_n293));
  NAND3_X1  g0093(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n227), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G13), .ZN(new_n297));
  NOR3_X1   g0097(.A1(new_n297), .A2(new_n204), .A3(G1), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n298), .A2(new_n295), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n203), .A2(G20), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n299), .A2(G50), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n298), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n296), .B(new_n301), .C1(G50), .C2(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT9), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n281), .A2(new_n282), .A3(new_n304), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n305), .B(KEYINPUT10), .ZN(new_n306));
  INV_X1    g0106(.A(G179), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n280), .A2(new_n307), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n308), .B(new_n303), .C1(G169), .C2(new_n280), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT74), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(new_n251), .B2(G33), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n249), .A2(KEYINPUT74), .A3(KEYINPUT3), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n313), .A2(new_n252), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n204), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n284), .B1(new_n316), .B2(KEYINPUT7), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT75), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n313), .A2(new_n314), .A3(KEYINPUT75), .A4(new_n252), .ZN(new_n320));
  NOR2_X1   g0120(.A1(KEYINPUT7), .A2(G20), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n317), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT76), .ZN(new_n324));
  XNOR2_X1  g0124(.A(G58), .B(G68), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n325), .A2(G20), .B1(G159), .B2(new_n289), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT76), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n317), .A2(new_n327), .A3(new_n322), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n324), .A2(KEYINPUT16), .A3(new_n326), .A4(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n250), .A2(new_n252), .ZN(new_n330));
  AND3_X1   g0130(.A1(new_n330), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n331));
  AOI21_X1  g0131(.A(KEYINPUT7), .B1(new_n330), .B2(new_n204), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n326), .B1(new_n333), .B2(new_n284), .ZN(new_n334));
  XNOR2_X1  g0134(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n329), .A2(new_n336), .A3(new_n295), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n286), .B1(new_n203), .B2(G20), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n338), .A2(new_n299), .B1(new_n298), .B2(new_n286), .ZN(new_n339));
  INV_X1    g0139(.A(new_n248), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n256), .A2(new_n258), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(G226), .B2(new_n258), .ZN(new_n342));
  INV_X1    g0142(.A(G87), .ZN(new_n343));
  OAI22_X1  g0143(.A1(new_n315), .A2(new_n342), .B1(new_n249), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT78), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n340), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(new_n345), .B2(new_n344), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n271), .B1(G232), .B2(new_n274), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n347), .A2(G190), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n347), .A2(new_n348), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(G200), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n337), .A2(new_n339), .A3(new_n349), .A4(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(KEYINPUT79), .A2(KEYINPUT17), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT79), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT17), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OR3_X1    g0156(.A1(new_n352), .A2(new_n353), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n337), .A2(new_n339), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n350), .A2(G169), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n307), .B2(new_n350), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT18), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT18), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n358), .A2(new_n360), .A3(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n352), .A2(new_n354), .A3(new_n355), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n357), .A2(new_n362), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n215), .A2(G1698), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(G226), .B2(G1698), .ZN(new_n369));
  OAI22_X1  g0169(.A1(new_n369), .A2(new_n330), .B1(new_n249), .B2(new_n216), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n248), .ZN(new_n371));
  INV_X1    g0171(.A(G238), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n371), .B(new_n270), .C1(new_n372), .C2(new_n273), .ZN(new_n373));
  OR2_X1    g0173(.A1(new_n373), .A2(KEYINPUT13), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(KEYINPUT13), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT14), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n376), .A2(new_n377), .A3(G169), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(new_n307), .B2(new_n376), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n377), .B1(new_n376), .B2(G169), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n298), .A2(new_n284), .ZN(new_n383));
  XNOR2_X1  g0183(.A(new_n383), .B(KEYINPUT12), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n284), .A2(G20), .ZN(new_n385));
  INV_X1    g0185(.A(G50), .ZN(new_n386));
  OAI221_X1 g0186(.A(new_n385), .B1(new_n287), .B2(new_n208), .C1(new_n290), .C2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n387), .A2(KEYINPUT11), .A3(new_n295), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n299), .A2(G68), .A3(new_n300), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n384), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT11), .B1(new_n387), .B2(new_n295), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n382), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n376), .A2(G200), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n374), .A2(G190), .A3(new_n375), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n395), .A2(new_n392), .A3(new_n396), .ZN(new_n397));
  XNOR2_X1  g0197(.A(new_n397), .B(KEYINPUT73), .ZN(new_n398));
  NOR3_X1   g0198(.A1(new_n330), .A2(new_n215), .A3(G1698), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT70), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT70), .ZN(new_n401));
  XOR2_X1   g0201(.A(KEYINPUT71), .B(G107), .Z(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n401), .B1(new_n403), .B2(new_n330), .ZN(new_n404));
  OAI221_X1 g0204(.A(new_n400), .B1(new_n404), .B2(new_n399), .C1(new_n255), .C2(new_n372), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n248), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n270), .B1(new_n273), .B2(new_n209), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT69), .ZN(new_n408));
  OR2_X1    g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n407), .A2(new_n408), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n406), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT72), .ZN(new_n412));
  OR3_X1    g0212(.A1(new_n411), .A2(new_n412), .A3(G179), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n412), .B1(new_n411), .B2(G179), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n299), .A2(G77), .A3(new_n300), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(G77), .B2(new_n302), .ZN(new_n416));
  NAND2_X1  g0216(.A1(G20), .A2(G77), .ZN(new_n417));
  XNOR2_X1  g0217(.A(KEYINPUT15), .B(G87), .ZN(new_n418));
  OAI221_X1 g0218(.A(new_n417), .B1(new_n286), .B2(new_n290), .C1(new_n287), .C2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n416), .B1(new_n419), .B2(new_n295), .ZN(new_n420));
  INV_X1    g0220(.A(G169), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n420), .B1(new_n411), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n413), .A2(new_n414), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n411), .A2(G200), .ZN(new_n424));
  INV_X1    g0224(.A(G190), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n424), .B(new_n420), .C1(new_n425), .C2(new_n411), .ZN(new_n426));
  AND4_X1   g0226(.A1(new_n394), .A2(new_n398), .A3(new_n423), .A4(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n311), .A2(new_n367), .A3(new_n427), .ZN(new_n428));
  XNOR2_X1  g0228(.A(KEYINPUT5), .B(G41), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n203), .A2(G45), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  AND2_X1   g0232(.A1(new_n432), .A2(new_n267), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(G270), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n267), .A2(G274), .A3(new_n431), .A4(new_n429), .ZN(new_n435));
  AND3_X1   g0235(.A1(new_n313), .A2(new_n252), .A3(new_n314), .ZN(new_n436));
  NOR2_X1   g0236(.A1(G257), .A2(G1698), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n437), .B1(new_n211), .B2(G1698), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n436), .A2(new_n438), .B1(G303), .B2(new_n330), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n434), .B(new_n435), .C1(new_n340), .C2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n441), .A2(new_n421), .ZN(new_n442));
  NAND2_X1  g0242(.A1(G33), .A2(G283), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n443), .B(new_n204), .C1(G33), .C2(new_n216), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n444), .B(new_n295), .C1(new_n204), .C2(G116), .ZN(new_n445));
  XOR2_X1   g0245(.A(new_n445), .B(KEYINPUT20), .Z(new_n446));
  NOR2_X1   g0246(.A1(new_n302), .A2(G116), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n299), .B1(G1), .B2(new_n249), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n447), .B1(new_n449), .B2(G116), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(KEYINPUT21), .B1(new_n442), .B2(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n451), .A2(KEYINPUT21), .A3(G169), .A4(new_n440), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n441), .A2(new_n451), .A3(G179), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n451), .B1(G200), .B2(new_n440), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n457), .B1(new_n425), .B2(new_n440), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n436), .A2(new_n204), .A3(G68), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT19), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n402), .A2(new_n343), .A3(new_n216), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n204), .B1(new_n249), .B2(new_n216), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n287), .A2(KEYINPUT19), .A3(new_n216), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n460), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n466), .A2(new_n295), .B1(new_n298), .B2(new_n418), .ZN(new_n467));
  INV_X1    g0267(.A(new_n418), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n449), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  OR2_X1    g0270(.A1(new_n430), .A2(G274), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n267), .B(new_n471), .C1(G250), .C2(new_n431), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT82), .ZN(new_n473));
  OR2_X1    g0273(.A1(new_n431), .A2(G250), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT82), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n267), .A2(new_n474), .A3(new_n475), .A4(new_n471), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G116), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n209), .A2(G1698), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n479), .B1(G238), .B2(G1698), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n478), .B1(new_n315), .B2(new_n480), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n481), .A2(new_n248), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n421), .B1(new_n477), .B2(new_n483), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n477), .A2(new_n483), .A3(G179), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n470), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n482), .B1(new_n473), .B2(new_n476), .ZN(new_n487));
  INV_X1    g0287(.A(G200), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n449), .A2(G87), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n477), .A2(new_n483), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n467), .B(new_n490), .C1(new_n425), .C2(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n486), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n459), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n433), .A2(G264), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n217), .A2(G1698), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(G250), .B2(G1698), .ZN(new_n497));
  INV_X1    g0297(.A(G294), .ZN(new_n498));
  OAI22_X1  g0298(.A1(new_n315), .A2(new_n497), .B1(new_n249), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n248), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n495), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT84), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT84), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n495), .A2(new_n503), .A3(new_n500), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n502), .A2(new_n435), .A3(new_n504), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n495), .A2(new_n435), .A3(new_n500), .ZN(new_n506));
  OAI22_X1  g0306(.A1(new_n505), .A2(new_n307), .B1(new_n421), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT25), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(new_n302), .B2(G107), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n298), .A2(KEYINPUT25), .A3(new_n210), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n449), .A2(G107), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT24), .ZN(new_n512));
  AND2_X1   g0312(.A1(new_n512), .A2(KEYINPUT83), .ZN(new_n513));
  OR2_X1    g0313(.A1(new_n204), .A2(KEYINPUT23), .ZN(new_n514));
  OAI22_X1  g0314(.A1(new_n514), .A2(G107), .B1(KEYINPUT83), .B2(new_n512), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n402), .A2(G20), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n515), .B1(new_n516), .B2(KEYINPUT23), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n204), .A2(G87), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n330), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n517), .B1(KEYINPUT22), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n436), .A2(KEYINPUT22), .A3(G87), .ZN(new_n521));
  AOI21_X1  g0321(.A(G20), .B1(new_n521), .B2(new_n478), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n513), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n295), .ZN(new_n524));
  NOR3_X1   g0324(.A1(new_n520), .A2(new_n522), .A3(new_n513), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n511), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n507), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n505), .A2(new_n488), .B1(new_n425), .B2(new_n506), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n529), .A2(new_n526), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT4), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n258), .A2(G244), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n532), .B1(new_n315), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n533), .A2(new_n532), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n535), .B1(G250), .B2(G1698), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n534), .B(new_n443), .C1(new_n536), .C2(new_n330), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n248), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n432), .A2(new_n267), .A3(G257), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n435), .A2(new_n539), .A3(KEYINPUT81), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n435), .A2(new_n539), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT81), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n538), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  OR2_X1    g0344(.A1(new_n544), .A2(G179), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT6), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n216), .A2(new_n210), .ZN(new_n547));
  NOR2_X1   g0347(.A1(G97), .A2(G107), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n210), .A2(KEYINPUT6), .A3(G97), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n204), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT80), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n290), .A2(new_n208), .ZN(new_n553));
  OR3_X1    g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n552), .B1(new_n551), .B2(new_n553), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n403), .B1(new_n331), .B2(new_n332), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n295), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n302), .A2(G97), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n559), .B1(new_n449), .B2(G97), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n544), .A2(new_n421), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n545), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n560), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n564), .B1(new_n557), .B2(new_n295), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n544), .A2(G200), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n565), .B(new_n566), .C1(new_n425), .C2(new_n544), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n494), .A2(new_n531), .A3(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n428), .A2(new_n569), .ZN(G372));
  INV_X1    g0370(.A(new_n397), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n394), .B1(new_n571), .B2(new_n423), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n572), .A2(new_n365), .A3(new_n357), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n362), .A2(new_n364), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n306), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n575), .A2(new_n309), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n487), .A2(G179), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n577), .B(KEYINPUT85), .C1(new_n421), .C2(new_n487), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT85), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(new_n485), .B2(new_n484), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n578), .A2(new_n580), .B1(new_n467), .B2(new_n469), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT86), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n487), .B2(new_n488), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n491), .A2(KEYINPUT86), .A3(G200), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n585), .A2(new_n492), .ZN(new_n586));
  NOR3_X1   g0386(.A1(new_n581), .A2(new_n586), .A3(new_n563), .ZN(new_n587));
  OAI21_X1  g0387(.A(KEYINPUT88), .B1(new_n587), .B2(KEYINPUT26), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n578), .A2(new_n580), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n470), .ZN(new_n590));
  INV_X1    g0390(.A(new_n563), .ZN(new_n591));
  OR2_X1    g0391(.A1(new_n585), .A2(new_n492), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT88), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT26), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n493), .A2(new_n563), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(KEYINPUT26), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n588), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n442), .A2(new_n451), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT21), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n455), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT87), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(KEYINPUT87), .B1(new_n452), .B2(new_n455), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n527), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n590), .A2(new_n592), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n563), .B(new_n567), .C1(new_n529), .C2(new_n526), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n581), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n599), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n576), .B1(new_n428), .B2(new_n613), .ZN(G369));
  NAND3_X1  g0414(.A1(new_n203), .A2(new_n204), .A3(G13), .ZN(new_n615));
  OR2_X1    g0415(.A1(new_n615), .A2(KEYINPUT27), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(KEYINPUT27), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n616), .A2(G213), .A3(new_n617), .ZN(new_n618));
  XOR2_X1   g0418(.A(KEYINPUT89), .B(G343), .Z(new_n619));
  NOR2_X1   g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n451), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n456), .A2(new_n458), .A3(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n622), .B1(new_n607), .B2(new_n621), .ZN(new_n623));
  XNOR2_X1  g0423(.A(new_n623), .B(KEYINPUT90), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n526), .A2(new_n620), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n531), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n620), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n626), .B1(new_n527), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n624), .A2(G330), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n528), .A2(new_n627), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n456), .A2(new_n620), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n531), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n629), .A2(new_n630), .A3(new_n632), .ZN(G399));
  INV_X1    g0433(.A(new_n224), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n634), .A2(G41), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n462), .A2(G116), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n636), .A2(G1), .A3(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n638), .B1(new_n229), .B2(new_n636), .ZN(new_n639));
  XNOR2_X1  g0439(.A(new_n639), .B(KEYINPUT28), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n456), .A2(new_n527), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n611), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n593), .A2(KEYINPUT26), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n597), .A2(new_n595), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(new_n644), .A3(new_n590), .ZN(new_n645));
  OAI211_X1 g0445(.A(KEYINPUT29), .B(new_n627), .C1(new_n642), .C2(new_n645), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n646), .A2(KEYINPUT91), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(KEYINPUT91), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n613), .A2(new_n620), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n647), .B(new_n648), .C1(KEYINPUT29), .C2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n441), .A2(G179), .A3(new_n487), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n502), .A2(new_n504), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n651), .A2(new_n652), .A3(new_n544), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n653), .A2(KEYINPUT30), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(KEYINPUT30), .ZN(new_n655));
  NOR3_X1   g0455(.A1(new_n441), .A2(new_n487), .A3(G179), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n656), .A2(new_n505), .A3(new_n544), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n654), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n620), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT31), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n494), .A2(new_n531), .A3(new_n568), .A4(new_n627), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n658), .A2(KEYINPUT31), .A3(new_n620), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(G330), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n650), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n640), .B1(new_n666), .B2(G1), .ZN(G364));
  NOR2_X1   g0467(.A1(new_n297), .A2(G20), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n203), .B1(new_n668), .B2(G45), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n636), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n671), .B1(new_n624), .B2(G330), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(G330), .B2(new_n624), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n227), .B1(G20), .B2(new_n421), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NOR4_X1   g0475(.A1(new_n204), .A2(new_n488), .A3(G179), .A4(G190), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(new_n210), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n204), .A2(new_n307), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(G200), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(new_n425), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(G179), .A2(G200), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n204), .B1(new_n683), .B2(G190), .ZN(new_n684));
  OAI22_X1  g0484(.A1(new_n682), .A2(new_n386), .B1(new_n684), .B2(new_n216), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n680), .A2(G190), .ZN(new_n686));
  AOI211_X1 g0486(.A(new_n678), .B(new_n685), .C1(G68), .C2(new_n686), .ZN(new_n687));
  NOR4_X1   g0487(.A1(new_n204), .A2(new_n425), .A3(new_n488), .A4(G179), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n688), .A2(KEYINPUT96), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(KEYINPUT96), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G87), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n683), .A2(G20), .A3(new_n425), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  XNOR2_X1  g0495(.A(KEYINPUT94), .B(G159), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g0497(.A(KEYINPUT95), .B(KEYINPUT32), .Z(new_n698));
  XNOR2_X1  g0498(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n679), .A2(G190), .A3(new_n488), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n253), .B1(new_n700), .B2(new_n214), .ZN(new_n701));
  NOR2_X1   g0501(.A1(G190), .A2(G200), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n679), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n701), .B1(G77), .B2(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n687), .A2(new_n693), .A3(new_n699), .A4(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n692), .A2(G303), .ZN(new_n707));
  INV_X1    g0507(.A(G311), .ZN(new_n708));
  INV_X1    g0508(.A(G329), .ZN(new_n709));
  OAI22_X1  g0509(.A1(new_n703), .A2(new_n708), .B1(new_n694), .B2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n700), .ZN(new_n711));
  AOI211_X1 g0511(.A(new_n253), .B(new_n710), .C1(G322), .C2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n684), .ZN(new_n713));
  AOI22_X1  g0513(.A1(new_n713), .A2(G294), .B1(new_n676), .B2(G283), .ZN(new_n714));
  XNOR2_X1  g0514(.A(KEYINPUT33), .B(G317), .ZN(new_n715));
  AOI22_X1  g0515(.A1(new_n715), .A2(new_n686), .B1(new_n681), .B2(G326), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n707), .A2(new_n712), .A3(new_n714), .A4(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n675), .B1(new_n706), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(G13), .A2(G33), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n204), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT93), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n721), .A2(new_n675), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n224), .A2(new_n253), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n723), .B1(KEYINPUT92), .B2(G355), .ZN(new_n724));
  OR2_X1    g0524(.A1(G355), .A2(KEYINPUT92), .ZN(new_n725));
  INV_X1    g0525(.A(G116), .ZN(new_n726));
  AOI22_X1  g0526(.A1(new_n724), .A2(new_n725), .B1(new_n726), .B2(new_n634), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n319), .A2(new_n320), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(new_n634), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n230), .A2(new_n268), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n731), .B1(new_n243), .B2(new_n268), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n727), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  AOI211_X1 g0533(.A(new_n670), .B(new_n718), .C1(new_n722), .C2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(new_n623), .B2(new_n721), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n673), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(G396));
  NOR2_X1   g0537(.A1(new_n420), .A2(new_n627), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n413), .A2(new_n414), .A3(new_n422), .A4(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n423), .A2(new_n426), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n739), .B1(new_n740), .B2(new_n738), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n649), .B(new_n741), .ZN(new_n742));
  OR2_X1    g0542(.A1(new_n742), .A2(new_n665), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n671), .B1(new_n742), .B2(new_n665), .ZN(new_n744));
  INV_X1    g0544(.A(new_n741), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(new_n719), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n692), .A2(G107), .ZN(new_n747));
  OAI22_X1  g0547(.A1(new_n703), .A2(new_n726), .B1(new_n694), .B2(new_n708), .ZN(new_n748));
  AOI211_X1 g0548(.A(new_n253), .B(new_n748), .C1(G294), .C2(new_n711), .ZN(new_n749));
  AOI22_X1  g0549(.A1(new_n713), .A2(G97), .B1(new_n676), .B2(G87), .ZN(new_n750));
  AOI22_X1  g0550(.A1(new_n686), .A2(G283), .B1(new_n681), .B2(G303), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n747), .A2(new_n749), .A3(new_n750), .A4(new_n751), .ZN(new_n752));
  AOI22_X1  g0552(.A1(new_n711), .A2(G143), .B1(new_n704), .B2(new_n696), .ZN(new_n753));
  INV_X1    g0553(.A(G137), .ZN(new_n754));
  INV_X1    g0554(.A(new_n686), .ZN(new_n755));
  OAI221_X1 g0555(.A(new_n753), .B1(new_n682), .B2(new_n754), .C1(new_n288), .C2(new_n755), .ZN(new_n756));
  XOR2_X1   g0556(.A(new_n756), .B(KEYINPUT34), .Z(new_n757));
  INV_X1    g0557(.A(G132), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n677), .A2(new_n284), .B1(new_n758), .B2(new_n694), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n759), .B1(G58), .B2(new_n713), .ZN(new_n760));
  OAI211_X1 g0560(.A(new_n760), .B(new_n728), .C1(new_n386), .C2(new_n691), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n752), .B1(new_n757), .B2(new_n761), .ZN(new_n762));
  AND2_X1   g0562(.A1(new_n762), .A2(new_n674), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n674), .A2(new_n719), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n670), .B(new_n763), .C1(new_n208), .C2(new_n764), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n743), .A2(new_n744), .B1(new_n746), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(G384));
  NOR2_X1   g0567(.A1(new_n668), .A2(new_n203), .ZN(new_n768));
  INV_X1    g0568(.A(G330), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n392), .A2(new_n627), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(new_n398), .B2(new_n381), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n394), .A2(new_n397), .A3(new_n771), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n775), .A2(new_n664), .A3(new_n741), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(KEYINPUT40), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n329), .A2(new_n295), .ZN(new_n778));
  INV_X1    g0578(.A(new_n335), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n327), .B1(new_n317), .B2(new_n322), .ZN(new_n780));
  INV_X1    g0580(.A(new_n326), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n779), .B1(new_n782), .B2(new_n328), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n339), .B1(new_n778), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n360), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(new_n352), .ZN(new_n786));
  INV_X1    g0586(.A(KEYINPUT98), .ZN(new_n787));
  AND3_X1   g0587(.A1(new_n317), .A2(new_n327), .A3(new_n322), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n788), .A2(new_n780), .A3(new_n781), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n295), .B(new_n329), .C1(new_n789), .C2(new_n779), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n787), .B(new_n618), .C1(new_n790), .C2(new_n339), .ZN(new_n791));
  INV_X1    g0591(.A(new_n618), .ZN(new_n792));
  AOI21_X1  g0592(.A(KEYINPUT98), .B1(new_n784), .B2(new_n792), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n786), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(KEYINPUT37), .ZN(new_n795));
  OAI21_X1  g0595(.A(KEYINPUT99), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n358), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n351), .A2(new_n349), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n797), .A2(new_n798), .B1(new_n784), .B2(new_n360), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n784), .A2(new_n792), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n787), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n784), .A2(KEYINPUT98), .A3(new_n792), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n799), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT99), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n803), .A2(new_n804), .A3(KEYINPUT37), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n358), .A2(new_n792), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n361), .A2(new_n806), .A3(new_n795), .A4(new_n352), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n796), .A2(new_n805), .A3(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n791), .A2(new_n793), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n366), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n808), .A2(KEYINPUT38), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(KEYINPUT38), .B1(new_n808), .B2(new_n811), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT100), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AND2_X1   g0615(.A1(new_n366), .A2(new_n810), .ZN(new_n816));
  INV_X1    g0616(.A(new_n807), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n803), .A2(KEYINPUT37), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n817), .B1(new_n818), .B2(KEYINPUT99), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n816), .B1(new_n819), .B2(new_n805), .ZN(new_n820));
  NOR3_X1   g0620(.A1(new_n820), .A2(KEYINPUT100), .A3(KEYINPUT38), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n777), .B1(new_n815), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT38), .ZN(new_n823));
  INV_X1    g0623(.A(new_n806), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n366), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n361), .A2(new_n806), .A3(new_n352), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(KEYINPUT37), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n827), .A2(KEYINPUT101), .A3(new_n807), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(KEYINPUT101), .B1(new_n827), .B2(new_n807), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n823), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n812), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n776), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(KEYINPUT40), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n822), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n428), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n837), .A2(new_n664), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n769), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n838), .B2(new_n836), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT102), .ZN(new_n841));
  OAI21_X1  g0641(.A(KEYINPUT100), .B1(new_n820), .B2(KEYINPUT38), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n808), .A2(new_n811), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n843), .A2(new_n814), .A3(new_n823), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n842), .A2(new_n844), .A3(new_n812), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n599), .A2(new_n612), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n846), .A2(new_n627), .A3(new_n741), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n423), .A2(new_n620), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n775), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n845), .A2(new_n852), .B1(new_n574), .B2(new_n618), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT39), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n812), .A2(new_n854), .A3(new_n831), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(new_n845), .B2(KEYINPUT39), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n382), .A2(new_n393), .A3(new_n627), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n853), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n576), .B1(new_n650), .B2(new_n428), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n858), .B(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n768), .B1(new_n841), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(new_n841), .B2(new_n860), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n228), .A2(G116), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n549), .A2(new_n550), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n863), .B1(new_n864), .B2(KEYINPUT35), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(KEYINPUT35), .B2(new_n864), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT36), .ZN(new_n867));
  OAI21_X1  g0667(.A(G77), .B1(new_n214), .B2(new_n284), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n868), .A2(new_n229), .B1(G50), .B2(new_n284), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n869), .A2(G1), .A3(new_n297), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n871), .B(KEYINPUT97), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n862), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n873), .B(KEYINPUT103), .ZN(G367));
  OAI221_X1 g0674(.A(new_n722), .B1(new_n224), .B2(new_n418), .C1(new_n730), .C2(new_n239), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n875), .A2(new_n671), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n627), .B1(new_n467), .B2(new_n490), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n581), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(new_n609), .B2(new_n877), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n711), .A2(G303), .B1(new_n704), .B2(G283), .ZN(new_n880));
  INV_X1    g0680(.A(G317), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n880), .B1(new_n881), .B2(new_n694), .ZN(new_n882));
  OAI22_X1  g0682(.A1(new_n755), .A2(new_n498), .B1(new_n682), .B2(new_n708), .ZN(new_n883));
  OAI22_X1  g0683(.A1(new_n677), .A2(new_n216), .B1(new_n402), .B2(new_n684), .ZN(new_n884));
  OR4_X1    g0684(.A1(new_n728), .A2(new_n882), .A3(new_n883), .A4(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n691), .A2(new_n726), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n886), .B(KEYINPUT46), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n691), .A2(new_n214), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n696), .A2(new_n686), .B1(new_n681), .B2(G143), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n330), .B1(new_n704), .B2(G50), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n711), .A2(G150), .B1(G137), .B2(new_n695), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n713), .A2(G68), .B1(new_n676), .B2(G77), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n889), .A2(new_n890), .A3(new_n891), .A4(new_n892), .ZN(new_n893));
  OAI22_X1  g0693(.A1(new_n885), .A2(new_n887), .B1(new_n888), .B2(new_n893), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(KEYINPUT107), .ZN(new_n895));
  XOR2_X1   g0695(.A(new_n895), .B(KEYINPUT47), .Z(new_n896));
  OAI221_X1 g0696(.A(new_n876), .B1(new_n721), .B2(new_n879), .C1(new_n896), .C2(new_n675), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n568), .B1(new_n565), .B2(new_n627), .ZN(new_n898));
  OR2_X1    g0698(.A1(new_n898), .A2(new_n527), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n620), .B1(new_n899), .B2(new_n563), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n591), .A2(new_n620), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n898), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(new_n531), .A3(new_n631), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n904), .B(KEYINPUT105), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT42), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n905), .A2(KEYINPUT42), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n901), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n879), .A2(KEYINPUT104), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT43), .B1(new_n879), .B2(KEYINPUT104), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n905), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT42), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n900), .B1(new_n916), .B2(new_n906), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n879), .A2(KEYINPUT43), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n912), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n903), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n913), .A2(new_n921), .B1(new_n629), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n909), .A2(new_n919), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n629), .A2(new_n922), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n924), .B(new_n925), .C1(new_n909), .C2(new_n912), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n669), .B(KEYINPUT106), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n632), .A2(new_n630), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n922), .A2(new_n930), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n931), .B(KEYINPUT44), .Z(new_n932));
  NOR2_X1   g0732(.A1(new_n922), .A2(new_n930), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT45), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n629), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n932), .A2(new_n629), .A3(new_n934), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n624), .A2(G330), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n632), .B1(new_n628), .B2(new_n631), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n940), .B(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n666), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n635), .B(KEYINPUT41), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n929), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n897), .B1(new_n927), .B2(new_n945), .ZN(G387));
  NOR2_X1   g0746(.A1(new_n628), .A2(new_n721), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n236), .A2(new_n268), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT109), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n637), .B(new_n268), .C1(new_n284), .C2(new_n208), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n950), .A2(KEYINPUT110), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(KEYINPUT110), .ZN(new_n952));
  OR3_X1    g0752(.A1(new_n286), .A2(KEYINPUT50), .A3(G50), .ZN(new_n953));
  OAI21_X1  g0753(.A(KEYINPUT50), .B1(new_n286), .B2(G50), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n951), .A2(new_n952), .A3(new_n953), .A4(new_n954), .ZN(new_n955));
  AND3_X1   g0755(.A1(new_n949), .A2(new_n729), .A3(new_n955), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n637), .A2(new_n723), .B1(G107), .B2(new_n224), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n722), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n728), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n700), .A2(new_n386), .B1(new_n288), .B2(new_n694), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(G68), .B2(new_n704), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n681), .A2(G159), .B1(G97), .B2(new_n676), .ZN(new_n962));
  INV_X1    g0762(.A(new_n286), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n686), .A2(new_n963), .B1(new_n468), .B2(new_n713), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n961), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n959), .B(new_n965), .C1(G77), .C2(new_n692), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n711), .A2(G317), .B1(new_n704), .B2(G303), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n681), .A2(G322), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n967), .B(new_n968), .C1(new_n708), .C2(new_n755), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT48), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n969), .A2(new_n970), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n692), .A2(G294), .B1(G283), .B2(new_n713), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT49), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n677), .A2(new_n726), .ZN(new_n976));
  AOI211_X1 g0776(.A(new_n976), .B(new_n728), .C1(G326), .C2(new_n695), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n966), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n958), .B(new_n671), .C1(new_n978), .C2(new_n675), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n947), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n942), .A2(new_n928), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n981), .A2(KEYINPUT108), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(KEYINPUT108), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n942), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n636), .B1(new_n666), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n666), .B2(new_n985), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n984), .A2(new_n987), .ZN(G393));
  NAND2_X1  g0788(.A1(new_n666), .A2(new_n985), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n989), .A2(new_n939), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n990), .A2(new_n636), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n939), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n937), .A2(new_n938), .A3(new_n929), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n722), .B1(new_n216), .B2(new_n224), .C1(new_n730), .C2(new_n246), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n670), .B1(new_n995), .B2(KEYINPUT111), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(KEYINPUT111), .B2(new_n995), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n682), .A2(new_n881), .B1(new_n708), .B2(new_n700), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT52), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n692), .A2(G283), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n684), .A2(new_n726), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n1001), .B(new_n678), .C1(G303), .C2(new_n686), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n330), .B1(new_n703), .B2(new_n498), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(G322), .B2(new_n695), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n999), .A2(new_n1000), .A3(new_n1002), .A4(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(G143), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n677), .A2(new_n343), .B1(new_n1006), .B2(new_n694), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n959), .B(new_n1007), .C1(new_n692), .C2(G68), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT113), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(G150), .A2(new_n681), .B1(new_n711), .B2(G159), .ZN(new_n1010));
  XOR2_X1   g0810(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n1011));
  XOR2_X1   g0811(.A(new_n1010), .B(new_n1011), .Z(new_n1012));
  AOI22_X1  g0812(.A1(new_n686), .A2(G50), .B1(new_n704), .B2(new_n963), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1012), .B(new_n1013), .C1(new_n208), .C2(new_n684), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1005), .B1(new_n1009), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n997), .B1(new_n1015), .B2(new_n674), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n903), .B2(new_n721), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n994), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n993), .A2(new_n1019), .ZN(G390));
  OR2_X1    g0820(.A1(new_n428), .A2(new_n665), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1021), .B(new_n576), .C1(new_n650), .C2(new_n428), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n773), .B(new_n774), .C1(new_n665), .C2(new_n745), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n775), .A2(new_n664), .A3(G330), .A4(new_n741), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n850), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n627), .B1(new_n642), .B2(new_n645), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n849), .B1(new_n1028), .B2(new_n745), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1024), .A2(new_n1030), .A3(new_n1025), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1027), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1023), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  AOI221_X4 g0834(.A(new_n855), .B1(new_n851), .B2(new_n857), .C1(new_n845), .C2(KEYINPUT39), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT114), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1025), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n857), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(new_n1029), .B2(new_n775), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1037), .B1(new_n1039), .B2(new_n832), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1025), .A2(new_n1036), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  NOR3_X1   g0843(.A1(new_n1035), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n845), .A2(KEYINPUT39), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n855), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1045), .B(new_n1046), .C1(new_n1038), .C2(new_n852), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1042), .B1(new_n1047), .B2(new_n1040), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1034), .B1(new_n1044), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1043), .B1(new_n1035), .B2(new_n1041), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1047), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1050), .A2(new_n1051), .A3(new_n1033), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1049), .A2(new_n635), .A3(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n929), .B1(new_n1044), .B2(new_n1048), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n670), .B1(new_n286), .B2(new_n764), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n691), .A2(new_n288), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT53), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n711), .A2(G132), .B1(G125), .B2(new_n695), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(KEYINPUT54), .B(G143), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1058), .B(new_n253), .C1(new_n703), .C2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n713), .A2(G159), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n755), .B2(new_n754), .ZN(new_n1062));
  INV_X1    g0862(.A(G128), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n682), .A2(new_n1063), .B1(new_n386), .B2(new_n677), .ZN(new_n1064));
  NOR3_X1   g0864(.A1(new_n1060), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1057), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT115), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1057), .A2(KEYINPUT115), .A3(new_n1065), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n686), .A2(new_n403), .B1(new_n704), .B2(G97), .ZN(new_n1070));
  INV_X1    g0870(.A(G283), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1070), .B1(new_n1071), .B2(new_n682), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT116), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n330), .B1(new_n694), .B2(new_n498), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(G116), .B2(new_n711), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n713), .A2(G77), .B1(new_n676), .B2(G68), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1073), .A2(new_n693), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  AND3_X1   g0877(.A1(new_n1068), .A2(new_n1069), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n719), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1055), .B1(new_n675), .B2(new_n1078), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1053), .A2(new_n1054), .A3(new_n1081), .ZN(G378));
  XOR2_X1   g0882(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n303), .A2(new_n792), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT55), .Z(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n306), .A2(new_n309), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1087), .B1(new_n306), .B2(new_n309), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1084), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1090), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1092), .A2(new_n1083), .A3(new_n1088), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n836), .B2(G330), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n769), .B(new_n1094), .C1(new_n822), .C2(new_n835), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n858), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n845), .A2(new_n777), .B1(new_n834), .B2(KEYINPUT40), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1094), .B1(new_n1099), .B2(new_n769), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n836), .A2(G330), .A3(new_n1095), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1079), .A2(new_n1038), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .A4(new_n853), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1098), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n929), .ZN(new_n1105));
  OR2_X1    g0905(.A1(new_n691), .A2(new_n1059), .ZN(new_n1106));
  OR2_X1    g0906(.A1(new_n1106), .A2(KEYINPUT117), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(KEYINPUT117), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n700), .A2(new_n1063), .B1(new_n703), .B2(new_n754), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(G132), .B2(new_n686), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n681), .A2(G125), .B1(G150), .B2(new_n713), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1107), .A2(new_n1108), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(KEYINPUT59), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n676), .A2(new_n696), .ZN(new_n1114));
  AOI211_X1 g0914(.A(G33), .B(G41), .C1(new_n695), .C2(G124), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1112), .A2(KEYINPUT59), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n711), .A2(G107), .B1(G283), .B2(new_n695), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n418), .B2(new_n703), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n755), .A2(new_n216), .B1(new_n684), .B2(new_n284), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n682), .A2(new_n726), .B1(new_n214), .B2(new_n677), .ZN(new_n1122));
  NOR3_X1   g0922(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n728), .A2(G41), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1123), .B(new_n1124), .C1(new_n208), .C2(new_n691), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT58), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1124), .ZN(new_n1127));
  AOI21_X1  g0927(.A(G50), .B1(new_n249), .B2(new_n262), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n1125), .A2(new_n1126), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n1126), .B2(new_n1125), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n674), .B1(new_n1118), .B2(new_n1130), .ZN(new_n1131));
  XOR2_X1   g0931(.A(new_n1131), .B(KEYINPUT118), .Z(new_n1132));
  AOI21_X1  g0932(.A(new_n670), .B1(new_n386), .B2(new_n764), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT119), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1132), .B(new_n1134), .C1(new_n1095), .C2(new_n1080), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1105), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT121), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1138), .B1(new_n1139), .B2(new_n858), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n1104), .B2(new_n1138), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1033), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1142));
  OAI21_X1  g0942(.A(KEYINPUT57), .B1(new_n1142), .B2(new_n1022), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n635), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1049), .A2(new_n1023), .ZN(new_n1145));
  AOI21_X1  g0945(.A(KEYINPUT57), .B1(new_n1145), .B2(new_n1104), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1137), .B1(new_n1144), .B2(new_n1146), .ZN(G375));
  AND2_X1   g0947(.A1(new_n1027), .A2(new_n1031), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n1022), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1033), .A2(new_n1149), .A3(new_n944), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n670), .B1(new_n284), .B2(new_n764), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n253), .B1(G303), .B2(new_n695), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1152), .B1(new_n1071), .B2(new_n700), .C1(new_n402), .C2(new_n703), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n755), .A2(new_n726), .B1(new_n682), .B2(new_n498), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n677), .A2(new_n208), .B1(new_n418), .B2(new_n684), .ZN(new_n1155));
  NOR3_X1   g0955(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n692), .A2(G97), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n704), .A2(G150), .B1(new_n695), .B2(G128), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n754), .B2(new_n700), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n755), .A2(new_n1059), .B1(new_n214), .B2(new_n677), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n682), .A2(new_n758), .B1(new_n684), .B2(new_n386), .ZN(new_n1161));
  NOR3_X1   g0961(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n959), .B1(new_n692), .B2(G159), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1156), .A2(new_n1157), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1151), .B1(new_n675), .B2(new_n1164), .C1(new_n775), .C2(new_n1080), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n1148), .B2(new_n928), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1150), .A2(new_n1167), .ZN(G381));
  AOI21_X1  g0968(.A(new_n1018), .B1(new_n991), .B2(new_n992), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1169), .B(new_n897), .C1(new_n945), .C2(new_n927), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n984), .A2(new_n987), .A3(new_n736), .A4(new_n766), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n1170), .A2(G381), .A3(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT122), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n1053), .A2(new_n1054), .A3(new_n1081), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1104), .A2(new_n1138), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1140), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT57), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n1049), .B2(new_n1023), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n636), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1146), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1136), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1173), .A2(new_n1174), .A3(new_n1182), .ZN(G407));
  NAND2_X1  g0983(.A1(new_n619), .A2(G213), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT123), .Z(new_n1185));
  NAND3_X1  g0985(.A1(new_n1182), .A2(new_n1174), .A3(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(G407), .A2(G213), .A3(new_n1186), .ZN(G409));
  OAI211_X1 g0987(.A(G378), .B(new_n1137), .C1(new_n1144), .C2(new_n1146), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1141), .A2(new_n928), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1104), .B(new_n944), .C1(new_n1142), .C2(new_n1022), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n1135), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1174), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1188), .A2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1148), .A2(KEYINPUT60), .A3(new_n1022), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n1194), .A2(new_n635), .ZN(new_n1195));
  OAI21_X1  g0995(.A(KEYINPUT60), .B1(new_n1148), .B2(new_n1022), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(new_n1149), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1195), .A2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(G384), .B1(new_n1198), .B2(new_n1167), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n766), .B(new_n1166), .C1(new_n1195), .C2(new_n1197), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1193), .A2(new_n1184), .A3(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT63), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1201), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n1185), .A2(G2897), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT125), .ZN(new_n1208));
  XOR2_X1   g1008(.A(KEYINPUT124), .B(G2897), .Z(new_n1209));
  NAND3_X1  g1009(.A1(new_n619), .A2(new_n1209), .A3(G213), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1208), .B1(new_n1201), .B2(new_n1210), .ZN(new_n1211));
  AND3_X1   g1011(.A1(new_n619), .A2(new_n1209), .A3(G213), .ZN(new_n1212));
  NOR4_X1   g1012(.A1(new_n1199), .A2(new_n1200), .A3(KEYINPUT125), .A4(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1207), .B1(new_n1211), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1193), .A2(new_n1184), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(G390), .A2(G387), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT126), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1170), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(G393), .B(new_n736), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT127), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1220), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1170), .A2(new_n1218), .A3(KEYINPUT127), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1220), .A2(new_n1223), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n1221), .ZN(new_n1228));
  AOI21_X1  g1028(.A(KEYINPUT61), .B1(new_n1226), .B2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1185), .B1(new_n1188), .B2(new_n1192), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1230), .A2(KEYINPUT63), .A3(new_n1201), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1204), .A2(new_n1217), .A3(new_n1229), .A4(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT61), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(new_n1230), .B2(new_n1214), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT62), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1202), .A2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1230), .A2(KEYINPUT62), .A3(new_n1201), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1234), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1226), .A2(new_n1228), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1232), .B1(new_n1238), .B2(new_n1240), .ZN(G405));
  NAND2_X1  g1041(.A1(G375), .A2(new_n1174), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1242), .A2(new_n1205), .A3(new_n1188), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1188), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1201), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1239), .A2(new_n1243), .A3(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1239), .B1(new_n1245), .B2(new_n1243), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1246), .A2(new_n1247), .ZN(G402));
endmodule


