//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 1 0 1 0 0 1 0 0 0 1 1 0 0 0 1 1 0 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n456, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n562, new_n564, new_n565, new_n566,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n579, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n616, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1211, new_n1212, new_n1213;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  XOR2_X1   g028(.A(G325), .B(KEYINPUT66), .Z(G261));
  AOI22_X1  g029(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n452), .ZN(G319));
  NAND2_X1  g030(.A1(G113), .A2(G2104), .ZN(new_n456));
  INV_X1    g031(.A(G2104), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(KEYINPUT3), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G125), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n456), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n465), .A2(G101), .A3(G2104), .ZN(new_n466));
  XNOR2_X1  g041(.A(new_n466), .B(KEYINPUT68), .ZN(new_n467));
  INV_X1    g042(.A(G137), .ZN(new_n468));
  OAI21_X1  g043(.A(KEYINPUT67), .B1(new_n457), .B2(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(new_n458), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n457), .A2(KEYINPUT67), .A3(KEYINPUT3), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n470), .A2(new_n465), .A3(new_n471), .ZN(new_n472));
  OAI211_X1 g047(.A(new_n464), .B(new_n467), .C1(new_n468), .C2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  NAND3_X1  g049(.A1(new_n470), .A2(G2105), .A3(new_n471), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  INV_X1    g052(.A(new_n472), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  OAI21_X1  g058(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  OAI21_X1  g060(.A(KEYINPUT69), .B1(new_n465), .B2(G114), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n487), .A2(new_n488), .A3(G2105), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n485), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT70), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n485), .A2(new_n486), .A3(new_n489), .A4(new_n492), .ZN(new_n493));
  AOI22_X1  g068(.A1(new_n476), .A2(G126), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n470), .A2(G138), .A3(new_n465), .A4(new_n471), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n461), .A2(KEYINPUT4), .ZN(new_n497));
  AND2_X1   g072(.A1(new_n465), .A2(G138), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT6), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(KEYINPUT71), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT6), .A3(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT5), .B(G543), .ZN(new_n510));
  AND3_X1   g085(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n509), .B1(new_n508), .B2(new_n510), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G88), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n515), .B1(new_n505), .B2(new_n507), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G50), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(KEYINPUT5), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT5), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G62), .ZN(new_n522));
  OAI21_X1  g097(.A(KEYINPUT73), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(G75), .A2(G543), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT73), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n510), .A2(new_n525), .A3(G62), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n523), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n514), .A2(new_n517), .A3(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  INV_X1    g105(.A(KEYINPUT74), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n508), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n505), .A2(KEYINPUT74), .A3(new_n507), .ZN(new_n533));
  AND3_X1   g108(.A1(new_n532), .A2(G543), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G51), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n508), .A2(new_n510), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(KEYINPUT72), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n537), .A2(G89), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n510), .A2(G63), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n541));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n541), .B(new_n542), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n535), .A2(new_n539), .A3(new_n540), .A4(new_n543), .ZN(G286));
  INV_X1    g119(.A(G286), .ZN(G168));
  NAND2_X1  g120(.A1(G77), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G64), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n521), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G651), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n532), .A2(G543), .A3(new_n533), .ZN(new_n550));
  INV_X1    g125(.A(G52), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n552), .B1(G90), .B2(new_n513), .ZN(G171));
  AOI22_X1  g128(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n554));
  OR2_X1    g129(.A1(new_n554), .A2(new_n504), .ZN(new_n555));
  INV_X1    g130(.A(G43), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n537), .A2(new_n538), .ZN(new_n557));
  INV_X1    g132(.A(G81), .ZN(new_n558));
  OAI221_X1 g133(.A(new_n555), .B1(new_n550), .B2(new_n556), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  AND3_X1   g136(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G36), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  XOR2_X1   g141(.A(new_n566), .B(KEYINPUT76), .Z(G188));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n534), .A2(KEYINPUT77), .A3(new_n568), .A4(G53), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n532), .A2(KEYINPUT77), .A3(G543), .A4(new_n533), .ZN(new_n570));
  INV_X1    g145(.A(G53), .ZN(new_n571));
  OAI21_X1  g146(.A(KEYINPUT9), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G65), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n521), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n513), .A2(G91), .B1(G651), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n573), .A2(new_n577), .ZN(G299));
  INV_X1    g153(.A(G90), .ZN(new_n579));
  OAI221_X1 g154(.A(new_n549), .B1(new_n550), .B2(new_n551), .C1(new_n557), .C2(new_n579), .ZN(G301));
  NAND2_X1  g155(.A1(new_n513), .A2(G87), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n534), .A2(G49), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(G288));
  INV_X1    g159(.A(G86), .ZN(new_n585));
  NOR3_X1   g160(.A1(new_n511), .A2(new_n512), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G61), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n521), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(G651), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n516), .A2(G48), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n586), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G305));
  INV_X1    g169(.A(G47), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  OAI22_X1  g171(.A1(new_n550), .A2(new_n595), .B1(new_n504), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n597), .B1(G85), .B2(new_n513), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  INV_X1    g175(.A(G92), .ZN(new_n601));
  OAI21_X1  g176(.A(KEYINPUT10), .B1(new_n557), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(G79), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G66), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n521), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n534), .A2(G54), .B1(G651), .B2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n513), .A2(new_n607), .A3(G92), .ZN(new_n608));
  AND3_X1   g183(.A1(new_n602), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n600), .B1(new_n609), .B2(G868), .ZN(G284));
  OAI21_X1  g185(.A(new_n600), .B1(new_n609), .B2(G868), .ZN(G321));
  NAND2_X1  g186(.A1(G286), .A2(G868), .ZN(new_n612));
  AND2_X1   g187(.A1(new_n573), .A2(new_n577), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(G868), .ZN(G297));
  OAI21_X1  g189(.A(new_n612), .B1(new_n613), .B2(G868), .ZN(G280));
  XNOR2_X1  g190(.A(KEYINPUT78), .B(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n609), .B1(G860), .B2(new_n616), .ZN(G148));
  NAND2_X1  g192(.A1(new_n609), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G868), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(G868), .B2(new_n560), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT80), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n624), .B(new_n625), .C1(G111), .C2(new_n465), .ZN(new_n626));
  INV_X1    g201(.A(G135), .ZN(new_n627));
  INV_X1    g202(.A(G123), .ZN(new_n628));
  OAI221_X1 g203(.A(new_n626), .B1(new_n472), .B2(new_n627), .C1(new_n628), .C2(new_n475), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(G2096), .Z(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n465), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT13), .B(G2100), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n630), .A2(new_n635), .ZN(G156));
  XOR2_X1   g211(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n637));
  XNOR2_X1  g212(.A(G2451), .B(G2454), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n637), .B(new_n638), .Z(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2427), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT83), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n642), .B(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT14), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT82), .B(KEYINPUT84), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  OR3_X1    g223(.A1(new_n645), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n648), .B1(new_n645), .B2(new_n646), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n649), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n652), .B1(new_n649), .B2(new_n650), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n640), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n655), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n657), .A2(new_n639), .A3(new_n653), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1341), .B(G1348), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT85), .Z(new_n661));
  AND3_X1   g236(.A1(new_n659), .A2(KEYINPUT86), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(G14), .B1(new_n659), .B2(new_n661), .ZN(new_n663));
  AOI21_X1  g238(.A(KEYINPUT86), .B1(new_n659), .B2(new_n661), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(G401));
  XOR2_X1   g240(.A(G2072), .B(G2078), .Z(new_n666));
  XOR2_X1   g241(.A(G2067), .B(G2678), .Z(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n666), .B1(new_n670), .B2(KEYINPUT18), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2096), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G2100), .ZN(new_n673));
  AND2_X1   g248(.A1(new_n670), .A2(KEYINPUT17), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n668), .A2(new_n669), .ZN(new_n675));
  AOI21_X1  g250(.A(KEYINPUT18), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n673), .B(new_n676), .Z(G227));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1971), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n678), .A2(new_n679), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT20), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n684), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n681), .A2(new_n683), .A3(new_n685), .ZN(new_n689));
  OAI211_X1 g264(.A(new_n688), .B(new_n689), .C1(new_n687), .C2(new_n686), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G1981), .ZN(new_n691));
  XOR2_X1   g266(.A(G1991), .B(G1996), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT87), .B(KEYINPUT88), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n693), .B(new_n697), .Z(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(G229));
  NOR2_X1   g274(.A1(G29), .A2(G35), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(G162), .B2(G29), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT29), .B(G2090), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G26), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT96), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT28), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n476), .A2(G128), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n478), .A2(G140), .ZN(new_n709));
  OR2_X1    g284(.A1(G104), .A2(G2105), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n710), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT94), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n708), .A2(new_n709), .A3(new_n713), .ZN(new_n714));
  AND3_X1   g289(.A1(new_n714), .A2(KEYINPUT95), .A3(G29), .ZN(new_n715));
  AOI21_X1  g290(.A(KEYINPUT95), .B1(new_n714), .B2(G29), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n707), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G2067), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n717), .A2(new_n718), .ZN(new_n720));
  INV_X1    g295(.A(G1966), .ZN(new_n721));
  NAND2_X1  g296(.A1(G168), .A2(G16), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G16), .B2(G21), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n719), .A2(new_n720), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT97), .B(KEYINPUT23), .Z(new_n725));
  INV_X1    g300(.A(G16), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G20), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n725), .B(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(new_n613), .B2(new_n726), .ZN(new_n729));
  INV_X1    g304(.A(G1956), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n723), .A2(new_n721), .ZN(new_n732));
  AND3_X1   g307(.A1(new_n724), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n726), .A2(G19), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n560), .B2(new_n726), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G1341), .ZN(new_n736));
  OR2_X1    g311(.A1(KEYINPUT24), .A2(G34), .ZN(new_n737));
  NAND2_X1  g312(.A1(KEYINPUT24), .A2(G34), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n737), .A2(new_n704), .A3(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G160), .B2(new_n704), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n740), .A2(G2084), .ZN(new_n741));
  OR2_X1    g316(.A1(G29), .A2(G32), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n476), .A2(G129), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n478), .A2(G141), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n465), .A2(G105), .A3(G2104), .ZN(new_n745));
  NAND3_X1  g320(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT26), .Z(new_n747));
  NAND4_X1  g322(.A1(new_n743), .A2(new_n744), .A3(new_n745), .A4(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n742), .B1(new_n748), .B2(new_n704), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT27), .B(G1996), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT30), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n753), .A2(G28), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(G28), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n754), .A2(new_n755), .A3(new_n704), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n751), .A2(new_n752), .A3(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT31), .B(G11), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  NOR4_X1   g334(.A1(new_n736), .A2(new_n741), .A3(new_n757), .A4(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n704), .A2(G27), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G164), .B2(new_n704), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n762), .A2(G2078), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n762), .A2(G2078), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n733), .A2(new_n760), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n740), .A2(G2084), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT25), .Z(new_n770));
  INV_X1    g345(.A(G139), .ZN(new_n771));
  INV_X1    g346(.A(new_n461), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n772), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n773));
  OAI221_X1 g348(.A(new_n770), .B1(new_n472), .B2(new_n771), .C1(new_n773), .C2(new_n465), .ZN(new_n774));
  MUX2_X1   g349(.A(G33), .B(new_n774), .S(G29), .Z(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(G2072), .Z(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n726), .A2(G5), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G171), .B2(new_n726), .ZN(new_n779));
  INV_X1    g354(.A(G1961), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  NOR4_X1   g357(.A1(new_n766), .A2(new_n768), .A3(new_n777), .A4(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT36), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n726), .A2(G23), .ZN(new_n785));
  INV_X1    g360(.A(G288), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n785), .B1(new_n786), .B2(new_n726), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT33), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(G1976), .ZN(new_n790));
  INV_X1    g365(.A(G1976), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n787), .A2(KEYINPUT33), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n787), .A2(KEYINPUT33), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n790), .A2(new_n794), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT91), .B(KEYINPUT34), .Z(new_n796));
  NAND2_X1  g371(.A1(new_n593), .A2(G16), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G6), .B2(G16), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n798), .A2(KEYINPUT32), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(KEYINPUT32), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(G1981), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n799), .A2(G1981), .A3(new_n800), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(G16), .A2(G22), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G166), .B2(G16), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT92), .B(G1971), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n795), .A2(new_n796), .A3(new_n805), .A4(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n796), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n790), .A2(new_n809), .A3(new_n794), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n803), .A2(new_n804), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n811), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(G25), .ZN(new_n816));
  OAI21_X1  g391(.A(KEYINPUT89), .B1(new_n816), .B2(G29), .ZN(new_n817));
  OR3_X1    g392(.A1(new_n816), .A2(KEYINPUT89), .A3(G29), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n476), .A2(G119), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n478), .A2(G131), .ZN(new_n820));
  OAI21_X1  g395(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n465), .A2(G107), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n819), .B(new_n820), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT90), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n817), .B(new_n818), .C1(new_n825), .C2(new_n704), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT35), .B(G1991), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n826), .B(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(G16), .A2(G24), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(new_n598), .B2(G16), .ZN(new_n831));
  INV_X1    g406(.A(G1986), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n784), .B1(new_n815), .B2(new_n835), .ZN(new_n836));
  AOI211_X1 g411(.A(KEYINPUT36), .B(new_n834), .C1(new_n810), .C2(new_n814), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n703), .B(new_n783), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT93), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(G4), .B2(G16), .ZN(new_n840));
  OR3_X1    g415(.A1(new_n839), .A2(G4), .A3(G16), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n602), .A2(new_n606), .A3(new_n608), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n840), .B(new_n841), .C1(new_n842), .C2(new_n726), .ZN(new_n843));
  INV_X1    g418(.A(G1348), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n629), .A2(new_n704), .ZN(new_n846));
  NOR3_X1   g421(.A1(new_n838), .A2(new_n845), .A3(new_n846), .ZN(G311));
  NOR2_X1   g422(.A1(new_n766), .A2(new_n782), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n848), .A2(new_n767), .A3(new_n776), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n815), .A2(new_n835), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(KEYINPUT36), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n815), .A2(new_n784), .A3(new_n835), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n849), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n845), .ZN(new_n854));
  INV_X1    g429(.A(new_n846), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n853), .A2(new_n854), .A3(new_n855), .A4(new_n703), .ZN(G150));
  XOR2_X1   g431(.A(KEYINPUT98), .B(G93), .Z(new_n857));
  AND3_X1   g432(.A1(new_n537), .A2(new_n538), .A3(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n534), .A2(G55), .ZN(new_n860));
  AOI22_X1  g435(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n861), .A2(new_n504), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n859), .A2(new_n860), .A3(KEYINPUT99), .A4(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT99), .ZN(new_n864));
  INV_X1    g439(.A(G55), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n862), .B1(new_n550), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n864), .B1(new_n866), .B2(new_n858), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(G860), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT37), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n609), .A2(G559), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT38), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n868), .A2(new_n559), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n866), .A2(new_n858), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n875), .A2(new_n559), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n873), .B(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n879), .A2(KEYINPUT39), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT100), .ZN(new_n881));
  INV_X1    g456(.A(new_n879), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT39), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n869), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n871), .B1(new_n881), .B2(new_n884), .ZN(G145));
  XNOR2_X1  g460(.A(new_n482), .B(new_n629), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n473), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n774), .A2(KEYINPUT101), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n774), .A2(KEYINPUT101), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n748), .B(new_n501), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(new_n714), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n892), .A2(new_n714), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n891), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n823), .B(KEYINPUT103), .ZN(new_n897));
  OAI21_X1  g472(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n898));
  OR2_X1    g473(.A1(new_n898), .A2(KEYINPUT102), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(KEYINPUT102), .ZN(new_n900));
  OAI211_X1 g475(.A(new_n899), .B(new_n900), .C1(G118), .C2(new_n465), .ZN(new_n901));
  INV_X1    g476(.A(G142), .ZN(new_n902));
  INV_X1    g477(.A(G130), .ZN(new_n903));
  OAI221_X1 g478(.A(new_n901), .B1(new_n472), .B2(new_n902), .C1(new_n903), .C2(new_n475), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(new_n633), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n897), .B(new_n905), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n892), .A2(new_n714), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n907), .A2(new_n890), .A3(new_n893), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n896), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n906), .B1(new_n896), .B2(new_n908), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n888), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n896), .A2(new_n908), .ZN(new_n912));
  INV_X1    g487(.A(new_n906), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n896), .A2(new_n906), .A3(new_n908), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(new_n915), .A3(new_n887), .ZN(new_n916));
  INV_X1    g491(.A(G37), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n911), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT104), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n911), .A2(new_n916), .A3(KEYINPUT104), .A4(new_n917), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g498(.A(KEYINPUT107), .ZN(new_n924));
  AND2_X1   g499(.A1(G303), .A2(G288), .ZN(new_n925));
  NOR2_X1   g500(.A1(G303), .A2(G288), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n593), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(G166), .A2(new_n786), .ZN(new_n928));
  NAND2_X1  g503(.A1(G303), .A2(G288), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n928), .A2(G305), .A3(new_n929), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n927), .A2(new_n930), .A3(new_n598), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n598), .B1(new_n927), .B2(new_n930), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT106), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(KEYINPUT42), .ZN(new_n935));
  OR2_X1    g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n934), .A2(KEYINPUT42), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n933), .A2(new_n937), .A3(new_n935), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  OR2_X1    g514(.A1(new_n618), .A2(KEYINPUT105), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n618), .A2(KEYINPUT105), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n878), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n940), .A2(new_n874), .A3(new_n877), .A4(new_n941), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n613), .A2(new_n609), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT41), .ZN(new_n947));
  NAND2_X1  g522(.A1(G299), .A2(new_n842), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n946), .A2(new_n948), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT41), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n945), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n943), .A2(new_n944), .A3(new_n950), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n939), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n943), .A2(new_n944), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n951), .A2(new_n949), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n953), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n957), .A2(new_n938), .A3(new_n936), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(G868), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n868), .A2(G868), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n924), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G868), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n964), .B1(new_n954), .B2(new_n958), .ZN(new_n965));
  NOR3_X1   g540(.A1(new_n965), .A2(KEYINPUT107), .A3(new_n961), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n963), .A2(new_n966), .ZN(G295));
  NAND2_X1  g542(.A1(new_n960), .A2(new_n962), .ZN(G331));
  XNOR2_X1  g543(.A(G301), .B(G286), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n969), .A2(new_n874), .A3(new_n877), .ZN(new_n970));
  XNOR2_X1  g545(.A(G171), .B(G286), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n560), .B1(new_n863), .B2(new_n867), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n971), .B1(new_n972), .B2(new_n876), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n956), .A2(new_n974), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n946), .A2(new_n948), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n970), .A2(new_n973), .A3(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n975), .A2(new_n933), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT108), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n975), .A2(new_n977), .ZN(new_n981));
  INV_X1    g556(.A(new_n933), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n975), .A2(new_n933), .A3(KEYINPUT108), .A4(new_n977), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n980), .A2(new_n983), .A3(new_n917), .A4(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT43), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n980), .A2(new_n917), .A3(new_n984), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n951), .A2(KEYINPUT110), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n976), .A2(new_n990), .A3(new_n947), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT110), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n950), .A2(new_n992), .A3(KEYINPUT41), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n949), .A2(KEYINPUT109), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n989), .A2(new_n991), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n974), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n933), .B1(new_n996), .B2(new_n977), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n988), .A2(new_n986), .A3(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(KEYINPUT44), .B1(new_n987), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n985), .A2(KEYINPUT43), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n988), .A2(KEYINPUT43), .A3(new_n997), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n999), .B1(new_n1003), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g579(.A(G1384), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n491), .A2(new_n493), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n470), .A2(G126), .A3(G2105), .A4(new_n471), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  AOI22_X1  g583(.A1(new_n495), .A2(KEYINPUT4), .B1(new_n498), .B2(new_n497), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1005), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT45), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n1013));
  OR2_X1    g588(.A1(new_n1013), .A2(G40), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(G40), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(G160), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1012), .A2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n714), .B(new_n718), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n748), .B(G1996), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1018), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  XOR2_X1   g597(.A(new_n827), .B(KEYINPUT112), .Z(new_n1023));
  NAND2_X1  g598(.A1(new_n823), .A2(new_n1023), .ZN(new_n1024));
  OR2_X1    g599(.A1(new_n823), .A2(new_n1023), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1018), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1022), .A2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n598), .B(new_n832), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1027), .B1(new_n1018), .B2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n1029), .B(KEYINPUT113), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT45), .B1(new_n501), .B2(new_n1005), .ZN(new_n1032));
  OAI211_X1 g607(.A(KEYINPUT45), .B(new_n1005), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1031), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G2078), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1017), .B1(new_n1012), .B2(KEYINPUT114), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(G1384), .B1(new_n494), .B2(new_n500), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT50), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1010), .A2(KEYINPUT50), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n473), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n780), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1039), .A2(G2078), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1048), .A2(G40), .A3(G160), .A4(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1040), .A2(new_n1047), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT125), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT125), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1040), .A2(new_n1053), .A3(new_n1047), .A4(new_n1050), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1052), .A2(G171), .A3(new_n1054), .ZN(new_n1055));
  AND4_X1   g630(.A1(new_n1012), .A2(new_n1045), .A3(new_n1033), .A4(new_n1049), .ZN(new_n1056));
  AOI221_X4 g631(.A(new_n1056), .B1(new_n780), .B2(new_n1046), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(G301), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1055), .A2(KEYINPUT54), .A3(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1040), .A2(G301), .A3(new_n1047), .A4(new_n1050), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1060), .B1(new_n1057), .B2(G301), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1012), .A2(new_n1045), .A3(new_n1033), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n721), .ZN(new_n1064));
  INV_X1    g639(.A(G2084), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1043), .A2(new_n1044), .A3(new_n1065), .A4(new_n1045), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1064), .A2(G168), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT51), .ZN(new_n1068));
  INV_X1    g643(.A(G8), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1069), .A2(KEYINPUT124), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1067), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1068), .B1(new_n1067), .B2(new_n1070), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  AOI211_X1 g648(.A(new_n1069), .B(G168), .C1(new_n1064), .C2(new_n1066), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  AOI22_X1  g650(.A1(new_n1061), .A2(new_n1062), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(G1981), .B1(new_n586), .B2(new_n592), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n589), .A2(G651), .B1(G48), .B2(new_n516), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1078), .B(new_n802), .C1(new_n557), .C2(new_n585), .ZN(new_n1079));
  OR2_X1    g654(.A1(KEYINPUT117), .A2(KEYINPUT49), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1077), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(KEYINPUT117), .A2(KEYINPUT49), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1069), .B1(new_n1045), .B2(new_n1041), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1077), .A2(new_n1079), .A3(KEYINPUT117), .A4(KEYINPUT49), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(KEYINPUT118), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT118), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1083), .A2(new_n1084), .A3(new_n1088), .A4(new_n1085), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1084), .B1(new_n791), .B2(G288), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT52), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT116), .B(G1976), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT52), .B1(G288), .B2(new_n1093), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1084), .B(new_n1094), .C1(new_n791), .C2(G288), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1090), .A2(new_n1092), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT115), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT55), .ZN(new_n1098));
  NAND4_X1  g673(.A1(G303), .A2(new_n1097), .A3(new_n1098), .A4(G8), .ZN(new_n1099));
  NAND2_X1  g674(.A1(G303), .A2(G8), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g676(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1099), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(G1971), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1045), .B1(new_n1032), .B2(new_n1031), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT114), .B1(new_n1012), .B2(new_n1033), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1105), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  OR2_X1    g683(.A1(new_n1046), .A2(G2090), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1104), .B1(new_n1110), .B2(G8), .ZN(new_n1111));
  AOI211_X1 g686(.A(new_n1069), .B(new_n1103), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n1096), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1059), .A2(new_n1076), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT120), .ZN(new_n1115));
  AOI21_X1  g690(.A(KEYINPUT57), .B1(new_n573), .B2(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n1116), .B(G299), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g693(.A(KEYINPUT56), .B(G2072), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1035), .A2(new_n1037), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1046), .A2(new_n730), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1118), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1045), .A2(new_n1041), .ZN(new_n1124));
  NOR3_X1   g699(.A1(new_n1124), .A2(KEYINPUT122), .A3(G2067), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1125), .B1(new_n844), .B2(new_n1046), .ZN(new_n1126));
  OAI21_X1  g701(.A(KEYINPUT122), .B1(new_n1124), .B2(G2067), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1123), .B1(new_n1128), .B2(new_n842), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1117), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1117), .A2(new_n1120), .A3(KEYINPUT121), .A4(new_n1121), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1129), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(G1996), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1035), .A2(new_n1135), .A3(new_n1037), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(KEYINPUT123), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1035), .A2(new_n1037), .A3(new_n1138), .A4(new_n1135), .ZN(new_n1139));
  XOR2_X1   g714(.A(KEYINPUT58), .B(G1341), .Z(new_n1140));
  NAND2_X1  g715(.A1(new_n1124), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1137), .A2(new_n1139), .A3(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n560), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n1143), .B(KEYINPUT59), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1126), .B(new_n1127), .C1(KEYINPUT60), .C2(new_n609), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n609), .A2(KEYINPUT60), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1145), .B(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1132), .A2(new_n1123), .A3(new_n1133), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT61), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n1130), .A2(KEYINPUT61), .ZN(new_n1150));
  AOI22_X1  g725(.A1(new_n1148), .A2(new_n1149), .B1(new_n1123), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1144), .A2(new_n1147), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1114), .B1(new_n1134), .B2(new_n1152), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1071), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT62), .ZN(new_n1155));
  OAI21_X1  g730(.A(KEYINPUT126), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1040), .A2(new_n1047), .ZN(new_n1157));
  OAI21_X1  g732(.A(G171), .B1(new_n1157), .B2(new_n1056), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1158), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1072), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1067), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1160), .A2(new_n1075), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1162), .A2(new_n1163), .A3(KEYINPUT62), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1156), .A2(new_n1159), .A3(new_n1113), .A4(new_n1164), .ZN(new_n1165));
  AND3_X1   g740(.A1(new_n1090), .A2(new_n1092), .A3(new_n1095), .ZN(new_n1166));
  AOI21_X1  g741(.A(G1971), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1046), .A2(G2090), .ZN(new_n1168));
  OAI21_X1  g743(.A(G8), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n1103), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1110), .A2(G8), .A3(new_n1104), .ZN(new_n1171));
  AOI211_X1 g746(.A(new_n1069), .B(G286), .C1(new_n1064), .C2(new_n1066), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1166), .A2(new_n1170), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT63), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT119), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1096), .A2(new_n1177), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1090), .A2(KEYINPUT119), .A3(new_n1092), .A4(new_n1095), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1176), .A2(KEYINPUT63), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1172), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1175), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  AND2_X1   g757(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1090), .A2(new_n791), .A3(new_n786), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1184), .A2(new_n1079), .ZN(new_n1185));
  AOI22_X1  g760(.A1(new_n1183), .A2(new_n1112), .B1(new_n1084), .B2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1165), .A2(new_n1182), .A3(new_n1186), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1030), .B1(new_n1153), .B2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n714), .A2(G2067), .ZN(new_n1189));
  AND2_X1   g764(.A1(new_n1022), .A2(new_n825), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1189), .B1(new_n1190), .B2(new_n828), .ZN(new_n1191));
  INV_X1    g766(.A(new_n1018), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1018), .A2(new_n832), .A3(new_n598), .ZN(new_n1193));
  XOR2_X1   g768(.A(new_n1193), .B(KEYINPUT48), .Z(new_n1194));
  OAI22_X1  g769(.A1(new_n1191), .A2(new_n1192), .B1(new_n1027), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT46), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1196), .B1(new_n1192), .B2(G1996), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1018), .B1(new_n1020), .B2(new_n748), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1018), .A2(KEYINPUT46), .A3(new_n1135), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g775(.A(KEYINPUT127), .B(KEYINPUT47), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n1200), .B(new_n1201), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1195), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1188), .A2(new_n1203), .ZN(G329));
  assign    G231 = 1'b0;
  OAI211_X1 g779(.A(G319), .B(new_n698), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1206));
  AOI21_X1  g780(.A(G401), .B1(new_n920), .B2(new_n921), .ZN(new_n1207));
  INV_X1    g781(.A(G227), .ZN(new_n1208));
  NAND2_X1  g782(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NOR2_X1   g783(.A1(new_n1206), .A2(new_n1209), .ZN(G308));
  AOI211_X1 g784(.A(G227), .B(G401), .C1(new_n920), .C2(new_n921), .ZN(new_n1211));
  OR2_X1    g785(.A1(new_n988), .A2(new_n997), .ZN(new_n1212));
  OAI21_X1  g786(.A(new_n1000), .B1(new_n1212), .B2(KEYINPUT43), .ZN(new_n1213));
  NAND4_X1  g787(.A1(new_n1211), .A2(new_n1213), .A3(G319), .A4(new_n698), .ZN(G225));
endmodule


