//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 0 0 0 1 0 0 0 1 0 0 0 0 0 0 1 0 0 1 1 1 1 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 1 0 0 1 0 1 0 1 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n612, new_n613, new_n614, new_n615, new_n616, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G469), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(new_n190), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT10), .ZN(new_n194));
  INV_X1    g008(.A(G104), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT3), .B1(new_n195), .B2(G107), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT3), .ZN(new_n197));
  INV_X1    g011(.A(G107), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(G104), .ZN(new_n199));
  INV_X1    g013(.A(G101), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n195), .A2(G107), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n196), .A2(new_n199), .A3(new_n200), .A4(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(G104), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n200), .B1(new_n203), .B2(new_n201), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(KEYINPUT78), .ZN(new_n205));
  XNOR2_X1  g019(.A(G104), .B(G107), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT78), .ZN(new_n207));
  NOR3_X1   g021(.A1(new_n206), .A2(new_n207), .A3(new_n200), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n202), .B1(new_n205), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n211), .A2(KEYINPUT1), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(new_n215), .A3(G128), .ZN(new_n216));
  INV_X1    g030(.A(G128), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n211), .B(new_n213), .C1(KEYINPUT1), .C2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n194), .B1(new_n209), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(G143), .B(G146), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT0), .B(G128), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n224));
  AND2_X1   g038(.A1(KEYINPUT0), .A2(G128), .ZN(new_n225));
  AOI22_X1  g039(.A1(new_n223), .A2(new_n224), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n196), .A2(new_n199), .A3(new_n201), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G101), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(KEYINPUT4), .A3(new_n202), .ZN(new_n229));
  OAI21_X1  g043(.A(KEYINPUT65), .B1(new_n221), .B2(new_n222), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT4), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n227), .A2(new_n231), .A3(G101), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n226), .A2(new_n229), .A3(new_n230), .A4(new_n232), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n216), .A2(new_n218), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n204), .A2(KEYINPUT78), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n207), .B1(new_n206), .B2(new_n200), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n234), .A2(KEYINPUT10), .A3(new_n237), .A4(new_n202), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n220), .A2(new_n233), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT11), .ZN(new_n240));
  INV_X1    g054(.A(G134), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n240), .B1(new_n241), .B2(G137), .ZN(new_n242));
  INV_X1    g056(.A(G137), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(KEYINPUT11), .A3(G134), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n241), .A2(G137), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n242), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G131), .ZN(new_n247));
  INV_X1    g061(.A(G131), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n242), .A2(new_n244), .A3(new_n248), .A4(new_n245), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n247), .A2(KEYINPUT66), .A3(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT66), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n246), .A2(new_n251), .A3(G131), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT68), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n250), .A2(KEYINPUT68), .A3(new_n252), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OR2_X1    g071(.A1(new_n239), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(G110), .B(G140), .ZN(new_n259));
  INV_X1    g073(.A(G953), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n260), .A2(G227), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n259), .B(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n258), .A2(new_n263), .ZN(new_n264));
  AND3_X1   g078(.A1(new_n250), .A2(KEYINPUT68), .A3(new_n252), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT68), .B1(new_n250), .B2(new_n252), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n209), .A2(new_n219), .ZN(new_n267));
  AOI22_X1  g081(.A1(new_n237), .A2(new_n202), .B1(new_n218), .B2(new_n216), .ZN(new_n268));
  OAI22_X1  g082(.A1(new_n265), .A2(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT12), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n209), .A2(new_n219), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n234), .A2(new_n202), .A3(new_n237), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n253), .A2(new_n270), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n269), .A2(new_n270), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  OR2_X1    g089(.A1(new_n264), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT79), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n239), .A2(new_n257), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n277), .B1(new_n239), .B2(new_n257), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n258), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n262), .ZN(new_n281));
  AOI21_X1  g095(.A(G902), .B1(new_n276), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n193), .B1(new_n282), .B2(new_n192), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n258), .B(new_n263), .C1(new_n278), .C2(new_n279), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n239), .A2(new_n257), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n262), .B1(new_n275), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n284), .A2(new_n286), .A3(G469), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n191), .B1(new_n283), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(G214), .B1(G237), .B2(G902), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(G110), .B(G122), .ZN(new_n291));
  XOR2_X1   g105(.A(new_n291), .B(KEYINPUT8), .Z(new_n292));
  XNOR2_X1  g106(.A(G116), .B(G119), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT5), .ZN(new_n294));
  INV_X1    g108(.A(G116), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n295), .A2(KEYINPUT5), .A3(G119), .ZN(new_n296));
  INV_X1    g110(.A(G113), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  XOR2_X1   g112(.A(KEYINPUT2), .B(G113), .Z(new_n299));
  AOI22_X1  g113(.A1(new_n294), .A2(new_n298), .B1(new_n299), .B2(new_n293), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n209), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n300), .A2(new_n237), .A3(new_n202), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n292), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n226), .A2(new_n230), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G125), .ZN(new_n306));
  INV_X1    g120(.A(G125), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n219), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n260), .A2(G224), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT7), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n306), .A2(new_n308), .A3(new_n311), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n304), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n303), .A2(KEYINPUT80), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n299), .B(new_n293), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(new_n229), .A3(new_n232), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT80), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n300), .A2(new_n237), .A3(new_n319), .A4(new_n202), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n316), .A2(new_n318), .A3(new_n320), .A4(new_n291), .ZN(new_n321));
  AOI21_X1  g135(.A(G902), .B1(new_n315), .B2(new_n321), .ZN(new_n322));
  XOR2_X1   g136(.A(new_n310), .B(KEYINPUT82), .Z(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n309), .B(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n316), .A2(new_n318), .A3(new_n320), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n291), .A2(KEYINPUT81), .ZN(new_n327));
  AOI22_X1  g141(.A1(KEYINPUT6), .A2(new_n321), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n326), .A2(KEYINPUT6), .A3(new_n327), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n325), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n322), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(G210), .B1(G237), .B2(G902), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n322), .A2(new_n330), .A3(new_n332), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n290), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(G113), .B(G122), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n337), .B(new_n195), .ZN(new_n338));
  INV_X1    g152(.A(G140), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G125), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n307), .A2(G140), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n340), .A2(new_n341), .A3(KEYINPUT74), .A4(KEYINPUT16), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n340), .A2(new_n341), .A3(KEYINPUT16), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT74), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n344), .B1(new_n340), .B2(KEYINPUT16), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n210), .B(new_n342), .C1(new_n343), .C2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n340), .A2(new_n341), .A3(KEYINPUT16), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n347), .B(new_n344), .C1(KEYINPUT16), .C2(new_n340), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n210), .B1(new_n348), .B2(new_n342), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n346), .B1(new_n349), .B2(KEYINPUT75), .ZN(new_n350));
  INV_X1    g164(.A(G237), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(new_n260), .A3(G214), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n212), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n351), .A2(new_n260), .A3(G143), .A4(G214), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(KEYINPUT17), .A3(G131), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(G131), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n353), .A2(new_n248), .A3(new_n354), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n356), .B1(new_n359), .B2(KEYINPUT17), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n342), .B1(new_n343), .B2(new_n345), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G146), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT75), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NOR3_X1   g178(.A1(new_n350), .A2(new_n360), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(KEYINPUT18), .A2(G131), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n366), .B1(new_n353), .B2(new_n354), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n367), .B(KEYINPUT83), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n340), .A2(new_n341), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n369), .B(new_n210), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n353), .A2(new_n354), .A3(new_n366), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n372), .B(KEYINPUT84), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n338), .B1(new_n365), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n338), .ZN(new_n376));
  XOR2_X1   g190(.A(new_n369), .B(KEYINPUT19), .Z(new_n377));
  OAI211_X1 g191(.A(new_n362), .B(new_n359), .C1(new_n377), .C2(G146), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n376), .B(new_n378), .C1(new_n371), .C2(new_n373), .ZN(new_n379));
  NOR2_X1   g193(.A1(G475), .A2(G902), .ZN(new_n380));
  XOR2_X1   g194(.A(new_n380), .B(KEYINPUT85), .Z(new_n381));
  NAND3_X1  g195(.A1(new_n375), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT20), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT20), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n375), .A2(new_n384), .A3(new_n379), .A4(new_n381), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n365), .A2(new_n374), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n376), .A2(KEYINPUT86), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n190), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n387), .A2(new_n388), .ZN(new_n391));
  OAI21_X1  g205(.A(G475), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n386), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G478), .ZN(new_n394));
  OR2_X1    g208(.A1(new_n394), .A2(KEYINPUT15), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n212), .A2(G128), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n217), .A2(G143), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n397), .A3(new_n241), .ZN(new_n398));
  INV_X1    g212(.A(G122), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G116), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n295), .A2(G122), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n402), .A2(G107), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n198), .B1(new_n400), .B2(new_n401), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n398), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT13), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n396), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n212), .A2(KEYINPUT13), .A3(G128), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(new_n408), .A3(new_n397), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n409), .A2(G134), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n295), .A2(G122), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n401), .B1(new_n413), .B2(KEYINPUT14), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(KEYINPUT87), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT87), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n416), .B(new_n401), .C1(new_n413), .C2(KEYINPUT14), .ZN(new_n417));
  OR2_X1    g231(.A1(new_n401), .A2(KEYINPUT14), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n415), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G107), .ZN(new_n420));
  INV_X1    g234(.A(new_n398), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n241), .B1(new_n396), .B2(new_n397), .ZN(new_n422));
  OAI22_X1  g236(.A1(new_n421), .A2(new_n422), .B1(G107), .B2(new_n402), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n189), .A2(G217), .A3(new_n260), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n412), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n423), .B1(new_n419), .B2(G107), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n426), .B1(new_n429), .B2(new_n411), .ZN(new_n430));
  AOI21_X1  g244(.A(G902), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT88), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n395), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n428), .A2(new_n430), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n190), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT88), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n431), .A2(new_n432), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n433), .B1(new_n438), .B2(new_n395), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  AOI211_X1 g254(.A(new_n190), .B(new_n260), .C1(G234), .C2(G237), .ZN(new_n441));
  XNOR2_X1  g255(.A(KEYINPUT21), .B(G898), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n260), .A2(G952), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n444), .B1(G234), .B2(G237), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n447), .B(KEYINPUT89), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NOR3_X1   g263(.A1(new_n393), .A2(new_n440), .A3(new_n449), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n288), .A2(new_n336), .A3(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(G472), .A2(G902), .ZN(new_n452));
  INV_X1    g266(.A(new_n317), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n241), .A2(G137), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n243), .A2(G134), .ZN(new_n455));
  OAI21_X1  g269(.A(G131), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n249), .A2(new_n456), .ZN(new_n457));
  OR2_X1    g271(.A1(new_n219), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT70), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n458), .B(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n305), .ZN(new_n462));
  AOI21_X1  g276(.A(KEYINPUT69), .B1(new_n257), .B2(new_n462), .ZN(new_n463));
  OAI211_X1 g277(.A(KEYINPUT69), .B(new_n462), .C1(new_n265), .C2(new_n266), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n453), .B(new_n461), .C1(new_n463), .C2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n351), .A2(new_n260), .A3(G210), .ZN(new_n467));
  XOR2_X1   g281(.A(new_n467), .B(KEYINPUT27), .Z(new_n468));
  XNOR2_X1  g282(.A(KEYINPUT26), .B(G101), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n468), .B(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n457), .A2(KEYINPUT67), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n234), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n457), .A2(KEYINPUT67), .ZN(new_n475));
  OAI22_X1  g289(.A1(new_n253), .A2(new_n305), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n317), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n462), .B1(new_n265), .B2(new_n266), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT69), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n460), .B1(new_n482), .B2(new_n464), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n479), .B1(new_n483), .B2(KEYINPUT30), .ZN(new_n484));
  OAI21_X1  g298(.A(KEYINPUT31), .B1(new_n472), .B2(new_n484), .ZN(new_n485));
  OAI211_X1 g299(.A(KEYINPUT30), .B(new_n461), .C1(new_n463), .C2(new_n465), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(new_n317), .A3(new_n478), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT31), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n470), .B1(new_n483), .B2(new_n453), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  XOR2_X1   g305(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n492));
  AOI211_X1 g306(.A(new_n317), .B(new_n460), .C1(new_n482), .C2(new_n464), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n476), .A2(new_n317), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n492), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n458), .A2(new_n453), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(KEYINPUT28), .B1(new_n480), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n471), .B1(new_n496), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n452), .B1(new_n491), .B2(new_n501), .ZN(new_n502));
  XOR2_X1   g316(.A(KEYINPUT72), .B(KEYINPUT32), .Z(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n492), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n506), .B1(new_n466), .B2(new_n494), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n471), .B1(new_n507), .B2(new_n499), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n487), .A2(new_n470), .A3(new_n466), .ZN(new_n509));
  AOI21_X1  g323(.A(KEYINPUT29), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n482), .A2(new_n464), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n453), .B1(new_n511), .B2(new_n461), .ZN(new_n512));
  OAI21_X1  g326(.A(KEYINPUT28), .B1(new_n512), .B2(new_n493), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n471), .A2(KEYINPUT29), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n500), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n190), .ZN(new_n516));
  OAI21_X1  g330(.A(G472), .B1(new_n510), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n470), .B1(new_n507), .B2(new_n499), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(new_n485), .A3(new_n490), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(KEYINPUT32), .A3(new_n452), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n505), .A2(new_n517), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(G234), .ZN(new_n522));
  OAI21_X1  g336(.A(G217), .B1(new_n522), .B2(G902), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n523), .B(KEYINPUT73), .ZN(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT22), .B(G137), .ZN(new_n525));
  NOR3_X1   g339(.A1(new_n187), .A2(new_n522), .A3(G953), .ZN(new_n526));
  XOR2_X1   g340(.A(new_n525), .B(new_n526), .Z(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT23), .ZN(new_n529));
  INV_X1    g343(.A(G119), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n529), .B1(new_n530), .B2(G128), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n217), .A2(KEYINPUT23), .A3(G119), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n531), .B(new_n532), .C1(G119), .C2(new_n217), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(G110), .ZN(new_n534));
  XOR2_X1   g348(.A(KEYINPUT24), .B(G110), .Z(new_n535));
  XNOR2_X1  g349(.A(G119), .B(G128), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n346), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n539), .B1(new_n363), .B2(new_n362), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n349), .A2(KEYINPUT75), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n538), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  XOR2_X1   g356(.A(KEYINPUT76), .B(G110), .Z(new_n543));
  OAI22_X1  g357(.A1(new_n533), .A2(new_n543), .B1(new_n536), .B2(new_n535), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n369), .A2(new_n210), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n362), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT77), .B1(new_n542), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n538), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n549), .B1(new_n350), .B2(new_n364), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT77), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n550), .A2(new_n551), .A3(new_n546), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n528), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n540), .A2(new_n541), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n547), .B1(new_n554), .B2(new_n549), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n527), .B1(new_n555), .B2(new_n551), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(KEYINPUT25), .B1(new_n557), .B2(new_n190), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT25), .ZN(new_n559));
  NOR4_X1   g373(.A1(new_n553), .A2(new_n556), .A3(new_n559), .A4(G902), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n524), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n524), .A2(G902), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n557), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n451), .A2(new_n521), .A3(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(G101), .ZN(G3));
  NAND2_X1  g381(.A1(new_n519), .A2(new_n190), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n568), .A2(G472), .B1(new_n452), .B2(new_n519), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n569), .A2(new_n565), .A3(new_n288), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n334), .A2(KEYINPUT90), .A3(new_n335), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n332), .B1(new_n322), .B2(new_n330), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT90), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n290), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AND2_X1   g388(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n448), .ZN(new_n576));
  INV_X1    g390(.A(new_n393), .ZN(new_n577));
  XOR2_X1   g391(.A(new_n434), .B(KEYINPUT33), .Z(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(G478), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n394), .A2(new_n190), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n580), .B1(new_n431), .B2(new_n394), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n577), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n576), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n570), .A2(new_n585), .ZN(new_n586));
  XOR2_X1   g400(.A(KEYINPUT34), .B(G104), .Z(new_n587));
  XNOR2_X1  g401(.A(new_n586), .B(new_n587), .ZN(G6));
  NAND2_X1  g402(.A1(new_n577), .A2(new_n440), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n576), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n570), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(KEYINPUT91), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(KEYINPUT92), .ZN(new_n593));
  XOR2_X1   g407(.A(KEYINPUT35), .B(G107), .Z(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(G9));
  NOR3_X1   g409(.A1(new_n542), .A2(KEYINPUT93), .A3(new_n547), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT93), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n597), .B1(new_n550), .B2(new_n546), .ZN(new_n598));
  OAI22_X1  g412(.A1(new_n596), .A2(new_n598), .B1(KEYINPUT36), .B2(new_n528), .ZN(new_n599));
  OAI21_X1  g413(.A(KEYINPUT93), .B1(new_n542), .B2(new_n547), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n528), .A2(KEYINPUT36), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n550), .A2(new_n597), .A3(new_n546), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n599), .A2(new_n603), .A3(new_n563), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(KEYINPUT94), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n561), .A2(new_n605), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n606), .A2(new_n450), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n607), .A2(new_n569), .A3(new_n288), .A4(new_n336), .ZN(new_n608));
  XOR2_X1   g422(.A(KEYINPUT37), .B(G110), .Z(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(KEYINPUT95), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n608), .B(new_n610), .ZN(G12));
  AND2_X1   g425(.A1(new_n288), .A2(new_n606), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT96), .B(G900), .Z(new_n613));
  AOI21_X1  g427(.A(new_n445), .B1(new_n441), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n589), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n521), .A2(new_n612), .A3(new_n575), .A4(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(G128), .ZN(G30));
  NAND2_X1  g431(.A1(new_n334), .A2(new_n335), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(KEYINPUT38), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n439), .B1(new_n386), .B2(new_n392), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n289), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n620), .A2(new_n606), .A3(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(new_n614), .B(KEYINPUT39), .Z(new_n624));
  NAND2_X1  g438(.A1(new_n288), .A2(new_n624), .ZN(new_n625));
  OR2_X1    g439(.A1(new_n625), .A2(KEYINPUT40), .ZN(new_n626));
  OR2_X1    g440(.A1(new_n512), .A2(new_n493), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n190), .B1(new_n627), .B2(new_n471), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n470), .B1(new_n487), .B2(new_n466), .ZN(new_n629));
  OAI21_X1  g443(.A(G472), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n505), .A2(new_n520), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n625), .A2(KEYINPUT40), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n623), .A2(new_n626), .A3(new_n631), .A4(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G143), .ZN(G45));
  INV_X1    g448(.A(new_n582), .ZN(new_n635));
  INV_X1    g449(.A(new_n614), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n635), .A2(new_n393), .A3(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n521), .A2(new_n612), .A3(new_n575), .A4(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G146), .ZN(G48));
  OR2_X1    g454(.A1(new_n282), .A2(new_n192), .ZN(new_n641));
  INV_X1    g455(.A(new_n191), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n239), .A2(new_n257), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(KEYINPUT79), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n239), .A2(new_n257), .A3(new_n277), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n263), .B1(new_n646), .B2(new_n258), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n264), .A2(new_n275), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n192), .B(new_n190), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n641), .A2(new_n642), .A3(new_n649), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n650), .A2(new_n562), .A3(new_n564), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n651), .A2(new_n521), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n585), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT41), .B(G113), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT97), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n653), .B(new_n655), .ZN(G15));
  NAND2_X1  g470(.A1(new_n652), .A2(new_n590), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G116), .ZN(G18));
  INV_X1    g472(.A(new_n650), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n521), .A2(new_n575), .A3(new_n607), .A4(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G119), .ZN(G21));
  NAND3_X1  g475(.A1(new_n621), .A2(new_n571), .A3(new_n574), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(KEYINPUT99), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT99), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n621), .A2(new_n571), .A3(new_n664), .A4(new_n574), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n666), .A2(new_n659), .A3(new_n448), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n471), .B1(new_n513), .B2(new_n500), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n452), .B1(new_n491), .B2(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(KEYINPUT98), .B1(new_n568), .B2(G472), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT98), .ZN(new_n671));
  INV_X1    g485(.A(G472), .ZN(new_n672));
  AOI211_X1 g486(.A(new_n671), .B(new_n672), .C1(new_n519), .C2(new_n190), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n565), .B(new_n669), .C1(new_n670), .C2(new_n673), .ZN(new_n674));
  OR2_X1    g488(.A1(new_n667), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G122), .ZN(G24));
  OR2_X1    g490(.A1(new_n670), .A2(new_n673), .ZN(new_n677));
  INV_X1    g491(.A(new_n575), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n678), .A2(new_n637), .A3(new_n650), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n677), .A2(new_n679), .A3(new_n606), .A4(new_n669), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G125), .ZN(G27));
  NOR2_X1   g495(.A1(new_n191), .A2(new_n290), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n334), .A2(new_n335), .A3(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT100), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n287), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n284), .A2(new_n286), .A3(KEYINPUT100), .A4(G469), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(KEYINPUT101), .B1(new_n688), .B2(new_n283), .ZN(new_n689));
  INV_X1    g503(.A(new_n193), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n649), .A2(new_n690), .A3(new_n686), .A4(new_n687), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT101), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n684), .B1(new_n689), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(KEYINPUT102), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n688), .A2(new_n283), .A3(KEYINPUT101), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n691), .A2(new_n692), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT102), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n698), .A2(new_n699), .A3(new_n684), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n695), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT32), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n502), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n703), .A2(new_n517), .A3(new_n520), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n565), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n701), .A2(new_n638), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n521), .A2(new_n565), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n708), .B1(new_n700), .B2(new_n695), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n637), .A2(KEYINPUT42), .ZN(new_n710));
  AOI22_X1  g524(.A1(new_n707), .A2(KEYINPUT42), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G131), .ZN(G33));
  INV_X1    g526(.A(new_n708), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n701), .A2(new_n713), .A3(new_n615), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G134), .ZN(G36));
  NAND2_X1  g529(.A1(new_n577), .A2(new_n635), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(KEYINPUT43), .ZN(new_n717));
  AOI211_X1 g531(.A(new_n569), .B(new_n717), .C1(new_n561), .C2(new_n605), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(KEYINPUT44), .ZN(new_n719));
  XOR2_X1   g533(.A(new_n719), .B(KEYINPUT105), .Z(new_n720));
  NAND2_X1  g534(.A1(new_n718), .A2(KEYINPUT44), .ZN(new_n721));
  XOR2_X1   g535(.A(new_n721), .B(KEYINPUT104), .Z(new_n722));
  AOI21_X1  g536(.A(KEYINPUT45), .B1(new_n284), .B2(new_n286), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n723), .A2(new_n192), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n284), .A2(new_n286), .A3(KEYINPUT45), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n690), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT46), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(KEYINPUT103), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n727), .A2(new_n728), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n730), .A2(new_n649), .A3(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(new_n642), .A3(new_n624), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n733), .A2(new_n290), .A3(new_n618), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n720), .A2(new_n722), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G137), .ZN(G39));
  NAND2_X1  g550(.A1(new_n732), .A2(new_n642), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT47), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n618), .A2(new_n290), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n638), .A2(new_n740), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n521), .A2(new_n565), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G140), .ZN(G42));
  NAND4_X1  g558(.A1(new_n565), .A2(new_n577), .A3(new_n635), .A4(new_n682), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(KEYINPUT106), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n641), .A2(new_n649), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(KEYINPUT49), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n746), .A2(new_n748), .A3(new_n619), .ZN(new_n749));
  INV_X1    g563(.A(new_n631), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n745), .A2(KEYINPUT106), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(G952), .A2(G953), .ZN(new_n753));
  XOR2_X1   g567(.A(new_n753), .B(KEYINPUT117), .Z(new_n754));
  NOR3_X1   g568(.A1(new_n674), .A2(new_n446), .A3(new_n717), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n755), .A2(new_n575), .A3(new_n659), .ZN(new_n756));
  NOR4_X1   g570(.A1(new_n717), .A2(new_n446), .A3(new_n747), .A4(new_n683), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(KEYINPUT113), .ZN(new_n758));
  OR2_X1    g572(.A1(new_n758), .A2(new_n705), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT48), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n759), .A2(new_n760), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n444), .B(KEYINPUT115), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n747), .A2(new_n446), .A3(new_n683), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n750), .A2(new_n565), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n763), .B1(new_n765), .B2(new_n583), .ZN(new_n766));
  AND4_X1   g580(.A1(new_n756), .A2(new_n761), .A3(new_n762), .A4(new_n766), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n747), .A2(KEYINPUT112), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n747), .A2(KEYINPUT112), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n768), .A2(new_n769), .A3(new_n642), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n740), .B(new_n755), .C1(new_n739), .C2(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n755), .A2(new_n290), .A3(new_n620), .A4(new_n659), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(KEYINPUT50), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n765), .A2(new_n577), .A3(new_n582), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n606), .B(new_n669), .C1(new_n670), .C2(new_n673), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n774), .B1(new_n758), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n771), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(KEYINPUT111), .B(KEYINPUT51), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n777), .A2(KEYINPUT114), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n771), .B(KEYINPUT51), .C1(new_n777), .C2(KEYINPUT114), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n767), .B(new_n780), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n561), .A2(new_n605), .A3(new_n636), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(KEYINPUT108), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT108), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n561), .A2(new_n605), .A3(new_n786), .A4(new_n636), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n191), .B1(new_n696), .B2(new_n697), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n788), .A2(new_n631), .A3(new_n666), .A4(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(KEYINPUT109), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n680), .A2(new_n616), .A3(new_n639), .ZN(new_n792));
  OAI21_X1  g606(.A(KEYINPUT52), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT109), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n790), .B(new_n794), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n680), .A2(new_n616), .A3(new_n639), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n393), .A2(new_n440), .A3(new_n614), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n521), .A2(new_n612), .A3(new_n740), .A4(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n802), .B1(new_n709), .B2(new_n615), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n699), .B1(new_n698), .B2(new_n684), .ZN(new_n804));
  AOI211_X1 g618(.A(KEYINPUT102), .B(new_n683), .C1(new_n696), .C2(new_n697), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n638), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(KEYINPUT42), .B1(new_n806), .B2(new_n705), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n709), .A2(new_n710), .ZN(new_n808));
  INV_X1    g622(.A(new_n775), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n701), .A2(new_n809), .A3(new_n638), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n803), .A2(new_n807), .A3(new_n808), .A4(new_n810), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n651), .B(new_n521), .C1(new_n585), .C2(new_n590), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n336), .A2(new_n448), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n813), .B1(new_n584), .B2(new_n589), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n570), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n812), .A2(new_n815), .A3(new_n660), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n608), .B(new_n566), .C1(new_n667), .C2(new_n674), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(KEYINPUT107), .B1(new_n811), .B2(new_n818), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n810), .A2(new_n714), .A3(new_n801), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n816), .A2(new_n817), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT107), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n820), .A2(new_n711), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n799), .B1(new_n819), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(KEYINPUT53), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n680), .A2(new_n616), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT52), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(KEYINPUT53), .ZN(new_n829));
  AOI211_X1 g643(.A(new_n829), .B(new_n799), .C1(new_n819), .C2(new_n823), .ZN(new_n830));
  OAI21_X1  g644(.A(KEYINPUT54), .B1(new_n825), .B2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n811), .A2(new_n818), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n828), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n833), .A2(new_n798), .A3(new_n793), .A4(new_n835), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n832), .B(new_n836), .C1(new_n824), .C2(KEYINPUT53), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n831), .A2(KEYINPUT110), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n819), .A2(new_n823), .ZN(new_n839));
  INV_X1    g653(.A(new_n799), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n834), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT110), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n842), .A2(new_n843), .A3(new_n832), .A4(new_n836), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n783), .B1(new_n838), .B2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n754), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI211_X1 g661(.A(KEYINPUT116), .B(new_n783), .C1(new_n838), .C2(new_n844), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n752), .B1(new_n847), .B2(new_n848), .ZN(G75));
  NOR2_X1   g663(.A1(new_n260), .A2(G952), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n836), .B1(new_n824), .B2(KEYINPUT53), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n851), .A2(G210), .A3(G902), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT56), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n328), .A2(new_n329), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(new_n325), .ZN(new_n856));
  XOR2_X1   g670(.A(new_n856), .B(KEYINPUT55), .Z(new_n857));
  AOI21_X1  g671(.A(new_n850), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n851), .A2(KEYINPUT118), .A3(G902), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT118), .B1(new_n851), .B2(G902), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n859), .A2(new_n860), .A3(new_n332), .ZN(new_n861));
  XNOR2_X1  g675(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n858), .B1(new_n861), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n858), .B(KEYINPUT120), .C1(new_n861), .C2(new_n864), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(G51));
  NAND2_X1  g683(.A1(new_n851), .A2(KEYINPUT54), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n837), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n193), .B(KEYINPUT57), .Z(new_n873));
  OAI22_X1  g687(.A1(new_n872), .A2(new_n873), .B1(new_n647), .B2(new_n648), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n859), .A2(new_n860), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n875), .A2(new_n725), .A3(new_n724), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n850), .B1(new_n874), .B2(new_n876), .ZN(G54));
  NAND3_X1  g691(.A1(new_n875), .A2(KEYINPUT58), .A3(G475), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n375), .A2(new_n379), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n850), .ZN(new_n881));
  INV_X1    g695(.A(new_n879), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n875), .A2(KEYINPUT58), .A3(G475), .A4(new_n882), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n880), .A2(new_n881), .A3(new_n883), .ZN(G60));
  XNOR2_X1  g698(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n885), .B(new_n580), .Z(new_n886));
  OAI21_X1  g700(.A(new_n824), .B1(KEYINPUT53), .B2(new_n828), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n832), .B1(new_n842), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n837), .A2(KEYINPUT110), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n844), .B(new_n886), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n578), .ZN(new_n891));
  INV_X1    g705(.A(new_n886), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n578), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n850), .B1(new_n871), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(KEYINPUT122), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n891), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n896), .A2(new_n898), .ZN(G63));
  AND2_X1   g713(.A1(new_n599), .A2(new_n603), .ZN(new_n900));
  NAND2_X1  g714(.A1(G217), .A2(G902), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT60), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n851), .A2(new_n900), .A3(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n557), .B1(new_n851), .B2(new_n903), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n905), .A2(new_n906), .A3(new_n850), .ZN(new_n907));
  OAI211_X1 g721(.A(KEYINPUT124), .B(KEYINPUT61), .C1(new_n907), .C2(KEYINPUT123), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT124), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n906), .A2(new_n850), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n904), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT123), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n909), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT61), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n914), .B1(new_n911), .B2(new_n909), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n908), .B1(new_n913), .B2(new_n915), .ZN(G66));
  INV_X1    g730(.A(G224), .ZN(new_n917));
  OAI21_X1  g731(.A(G953), .B1(new_n442), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n918), .B1(new_n821), .B2(G953), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n855), .B1(G898), .B2(new_n260), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n919), .B(new_n920), .ZN(G69));
  NAND2_X1  g735(.A1(new_n486), .A2(new_n478), .ZN(new_n922));
  XOR2_X1   g736(.A(KEYINPUT125), .B(KEYINPUT126), .Z(new_n923));
  XNOR2_X1  g737(.A(new_n922), .B(new_n923), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT127), .Z(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(new_n377), .Z(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n927), .B1(G900), .B2(G953), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n735), .A2(new_n796), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n706), .A2(new_n666), .ZN(new_n930));
  OR2_X1    g744(.A1(new_n733), .A2(new_n930), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n743), .A2(new_n714), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n929), .A2(new_n711), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n928), .B1(new_n933), .B2(G953), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n796), .A2(new_n633), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(KEYINPUT62), .ZN(new_n936));
  INV_X1    g750(.A(new_n625), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n584), .A2(new_n589), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n713), .A2(new_n937), .A3(new_n740), .A4(new_n938), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n735), .A2(new_n743), .A3(new_n936), .A4(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n935), .A2(KEYINPUT62), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n260), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n927), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n934), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n260), .B1(G227), .B2(G900), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n944), .B(new_n945), .ZN(G72));
  NAND2_X1  g760(.A1(G472), .A2(G902), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT63), .Z(new_n948));
  OAI21_X1  g762(.A(new_n948), .B1(new_n933), .B2(new_n818), .ZN(new_n949));
  INV_X1    g763(.A(new_n509), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n940), .A2(new_n818), .A3(new_n941), .ZN(new_n952));
  INV_X1    g766(.A(new_n948), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n629), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n951), .A2(new_n881), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n842), .A2(new_n887), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n950), .A2(new_n629), .A3(new_n953), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(G57));
endmodule


