//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 1 0 0 1 0 0 0 0 1 1 1 0 0 1 1 0 0 0 1 1 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 0 1 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1188, new_n1189,
    new_n1190, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n202), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n209), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  XOR2_X1   g0020(.A(KEYINPUT64), .B(G238), .Z(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  XOR2_X1   g0023(.A(KEYINPUT65), .B(G77), .Z(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT66), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n211), .B1(new_n225), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n214), .B(new_n219), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G226), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n246), .B(new_n247), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n217), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT8), .B(G58), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n209), .A2(G33), .ZN(new_n253));
  INV_X1    g0053(.A(G150), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  OAI22_X1  g0056(.A1(new_n252), .A2(new_n253), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G50), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n209), .B1(new_n201), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n251), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(new_n251), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n208), .A2(G20), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G50), .ZN(new_n266));
  XNOR2_X1  g0066(.A(new_n266), .B(KEYINPUT71), .ZN(new_n267));
  OAI221_X1 g0067(.A(new_n260), .B1(G50), .B2(new_n261), .C1(new_n264), .C2(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n268), .B(KEYINPUT9), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G33), .ZN(new_n272));
  INV_X1    g0072(.A(G41), .ZN(new_n273));
  OAI211_X1 g0073(.A(G1), .B(G13), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n271), .A2(new_n274), .A3(G274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n270), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT69), .B(G226), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT3), .B(G33), .ZN(new_n278));
  INV_X1    g0078(.A(G1698), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n278), .A2(G222), .A3(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n280), .B1(new_n224), .B2(new_n278), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT70), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n272), .A2(KEYINPUT3), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT3), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n282), .B1(new_n286), .B2(new_n279), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n278), .A2(KEYINPUT70), .A3(G1698), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n281), .B1(new_n289), .B2(G223), .ZN(new_n290));
  OAI221_X1 g0090(.A(new_n275), .B1(new_n276), .B2(new_n277), .C1(new_n290), .C2(new_n274), .ZN(new_n291));
  XOR2_X1   g0091(.A(KEYINPUT74), .B(G200), .Z(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G190), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n269), .B(new_n293), .C1(new_n294), .C2(new_n291), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT10), .ZN(new_n296));
  INV_X1    g0096(.A(G169), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n291), .A2(new_n297), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n298), .B(new_n268), .C1(G179), .C2(new_n291), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n262), .A2(new_n222), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n301), .B(KEYINPUT12), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n255), .A2(G50), .B1(G20), .B2(new_n222), .ZN(new_n303));
  INV_X1    g0103(.A(G77), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n303), .B1(new_n304), .B2(new_n253), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n305), .A2(KEYINPUT11), .A3(new_n251), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n263), .A2(G68), .A3(new_n265), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n302), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(KEYINPUT11), .B1(new_n305), .B2(new_n251), .ZN(new_n309));
  OR3_X1    g0109(.A1(new_n308), .A2(KEYINPUT75), .A3(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(KEYINPUT75), .B1(new_n308), .B2(new_n309), .ZN(new_n311));
  AND2_X1   g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n278), .A2(G226), .A3(new_n279), .ZN(new_n313));
  NAND2_X1  g0113(.A1(G33), .A2(G97), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n278), .A2(G232), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n313), .B(new_n314), .C1(new_n315), .C2(new_n279), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G274), .ZN(new_n319));
  NOR3_X1   g0119(.A1(new_n317), .A2(new_n319), .A3(new_n270), .ZN(new_n320));
  INV_X1    g0120(.A(new_n276), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n320), .B1(G238), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT13), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT13), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n318), .A2(new_n325), .A3(new_n322), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT14), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n327), .A2(new_n328), .A3(G169), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n324), .A2(G179), .A3(new_n326), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n328), .B1(new_n327), .B2(G169), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n312), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n327), .A2(G200), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n308), .A2(new_n309), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n334), .B(new_n335), .C1(new_n294), .C2(new_n327), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n221), .B1(new_n287), .B2(new_n288), .ZN(new_n338));
  OAI22_X1  g0138(.A1(new_n315), .A2(G1698), .B1(new_n205), .B2(new_n278), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT73), .ZN(new_n340));
  OR3_X1    g0140(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n340), .B1(new_n338), .B2(new_n339), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n341), .A2(new_n342), .A3(new_n317), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n275), .B1(new_n276), .B2(new_n223), .ZN(new_n344));
  XNOR2_X1  g0144(.A(new_n344), .B(KEYINPUT72), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n292), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n263), .A2(G77), .A3(new_n265), .ZN(new_n348));
  INV_X1    g0148(.A(new_n224), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n348), .B1(new_n349), .B2(new_n261), .ZN(new_n350));
  INV_X1    g0150(.A(new_n252), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n255), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT15), .B(G87), .ZN(new_n353));
  OAI221_X1 g0153(.A(new_n352), .B1(new_n209), .B2(new_n224), .C1(new_n253), .C2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n350), .B1(new_n354), .B2(new_n251), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n347), .B(new_n355), .C1(new_n294), .C2(new_n346), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n355), .B1(new_n346), .B2(new_n297), .ZN(new_n357));
  INV_X1    g0157(.A(G179), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n343), .A2(new_n358), .A3(new_n345), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  NOR3_X1   g0161(.A1(new_n300), .A2(new_n337), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n351), .A2(new_n265), .ZN(new_n363));
  OAI22_X1  g0163(.A1(new_n264), .A2(new_n363), .B1(new_n261), .B2(new_n351), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n278), .A2(G226), .A3(G1698), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n278), .A2(G223), .A3(new_n279), .ZN(new_n367));
  INV_X1    g0167(.A(G87), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n366), .B(new_n367), .C1(new_n272), .C2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n317), .ZN(new_n370));
  INV_X1    g0170(.A(G232), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n275), .B1(new_n276), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n370), .A2(new_n373), .A3(new_n294), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n372), .B1(new_n369), .B2(new_n317), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n374), .B1(G200), .B2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(KEYINPUT7), .B1(new_n286), .B2(new_n209), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT7), .ZN(new_n378));
  AOI211_X1 g0178(.A(new_n378), .B(G20), .C1(new_n283), .C2(new_n285), .ZN(new_n379));
  OAI21_X1  g0179(.A(G68), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  AND2_X1   g0180(.A1(G58), .A2(G68), .ZN(new_n381));
  OAI21_X1  g0181(.A(G20), .B1(new_n381), .B2(new_n201), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT76), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI211_X1 g0184(.A(KEYINPUT76), .B(G20), .C1(new_n381), .C2(new_n201), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n384), .A2(new_n385), .B1(G159), .B2(new_n255), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n380), .A2(KEYINPUT16), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT16), .B1(new_n380), .B2(new_n386), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT77), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n251), .B(new_n387), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  AOI211_X1 g0190(.A(KEYINPUT77), .B(KEYINPUT16), .C1(new_n380), .C2(new_n386), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n365), .B(new_n376), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  XOR2_X1   g0192(.A(new_n392), .B(KEYINPUT17), .Z(new_n393));
  OAI21_X1  g0193(.A(new_n365), .B1(new_n390), .B2(new_n391), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n375), .A2(G179), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n375), .A2(new_n297), .ZN(new_n396));
  OR2_X1    g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT18), .ZN(new_n398));
  AND3_X1   g0198(.A1(new_n394), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n398), .B1(new_n394), .B2(new_n397), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT78), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n380), .A2(new_n386), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT16), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n389), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n387), .A2(new_n251), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n391), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n364), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n395), .A2(new_n396), .ZN(new_n409));
  OAI21_X1  g0209(.A(KEYINPUT18), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT78), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n394), .A2(new_n397), .A3(new_n398), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n393), .B1(new_n401), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n362), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n262), .A2(KEYINPUT25), .A3(new_n205), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(KEYINPUT25), .B1(new_n262), .B2(new_n205), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n208), .A2(G33), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n261), .A2(new_n420), .A3(new_n217), .A4(new_n250), .ZN(new_n421));
  OAI22_X1  g0221(.A1(new_n418), .A2(new_n419), .B1(new_n205), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT23), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(new_n209), .B2(G107), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n205), .A2(KEYINPUT23), .A3(G20), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G33), .A2(G116), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n426), .B1(G20), .B2(new_n427), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n283), .A2(new_n285), .A3(new_n209), .A4(G87), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT22), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT22), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n278), .A2(new_n431), .A3(new_n209), .A4(G87), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n428), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n433), .A2(KEYINPUT85), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n433), .A2(KEYINPUT85), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(KEYINPUT24), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n251), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT24), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n438), .B1(new_n434), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n422), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n278), .A2(G257), .A3(G1698), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n278), .A2(G250), .A3(new_n279), .ZN(new_n443));
  NAND2_X1  g0243(.A1(G33), .A2(G294), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT87), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT87), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n442), .A2(new_n443), .A3(new_n447), .A4(new_n444), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n446), .A2(new_n317), .A3(new_n448), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n208), .B(G45), .C1(new_n273), .C2(KEYINPUT5), .ZN(new_n450));
  OR2_X1    g0250(.A1(new_n450), .A2(KEYINPUT79), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n317), .A2(new_n319), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(KEYINPUT79), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n273), .A2(KEYINPUT5), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n451), .A2(new_n452), .A3(new_n453), .A4(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n453), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n454), .B1(new_n450), .B2(KEYINPUT79), .ZN(new_n457));
  OAI211_X1 g0257(.A(G264), .B(new_n274), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n449), .A2(new_n455), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(G200), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n449), .A2(new_n294), .A3(new_n455), .A4(new_n458), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n441), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT88), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n441), .A2(new_n463), .A3(KEYINPUT88), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n436), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT24), .B1(new_n433), .B2(KEYINPUT85), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n440), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n422), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(KEYINPUT86), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT86), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n441), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n459), .A2(G169), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n477), .B1(new_n358), .B2(new_n459), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n474), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  AND2_X1   g0279(.A1(new_n468), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g0280(.A(G270), .B(new_n274), .C1(new_n456), .C2(new_n457), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n455), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n278), .A2(G264), .A3(G1698), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n278), .A2(G257), .A3(new_n279), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n286), .A2(G303), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT84), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n274), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT84), .A4(new_n485), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n482), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(G33), .A2(G283), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n491), .B(new_n209), .C1(G33), .C2(new_n204), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n492), .B(new_n251), .C1(new_n209), .C2(G116), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT20), .ZN(new_n494));
  XNOR2_X1  g0294(.A(new_n493), .B(new_n494), .ZN(new_n495));
  MUX2_X1   g0295(.A(new_n261), .B(new_n421), .S(G116), .Z(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n490), .A2(G179), .A3(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n490), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT21), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n499), .A2(new_n500), .A3(G169), .A4(new_n497), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n497), .A2(G169), .ZN(new_n502));
  OAI21_X1  g0302(.A(KEYINPUT21), .B1(new_n502), .B2(new_n490), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n498), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n278), .A2(G244), .A3(new_n279), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT4), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n278), .A2(KEYINPUT4), .A3(G244), .A4(new_n279), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n278), .A2(G250), .A3(G1698), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n507), .A2(new_n491), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n317), .ZN(new_n511));
  OAI211_X1 g0311(.A(G257), .B(new_n274), .C1(new_n456), .C2(new_n457), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n511), .A2(new_n455), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n297), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n205), .A2(KEYINPUT6), .A3(G97), .ZN(new_n515));
  XOR2_X1   g0315(.A(G97), .B(G107), .Z(new_n516));
  OAI21_X1  g0316(.A(new_n515), .B1(new_n516), .B2(KEYINPUT6), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n517), .A2(G20), .B1(G77), .B2(new_n255), .ZN(new_n518));
  OAI21_X1  g0318(.A(G107), .B1(new_n377), .B2(new_n379), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n438), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n262), .A2(new_n204), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(new_n421), .B2(new_n204), .ZN(new_n522));
  OR2_X1    g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n511), .A2(new_n358), .A3(new_n455), .A4(new_n512), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n514), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n520), .A2(new_n522), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n511), .A2(G190), .A3(new_n455), .A4(new_n512), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n512), .A2(new_n455), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n528), .B1(new_n317), .B2(new_n510), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n526), .B(new_n527), .C1(new_n460), .C2(new_n529), .ZN(new_n530));
  AND2_X1   g0330(.A1(new_n525), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n497), .B1(new_n499), .B2(G200), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(new_n294), .B2(new_n499), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n278), .A2(new_n209), .A3(G68), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT19), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n209), .B1(new_n314), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(G87), .B2(new_n206), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n535), .B1(new_n253), .B2(new_n204), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n534), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT81), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n438), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n534), .A2(new_n537), .A3(KEYINPUT81), .A4(new_n538), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n421), .A2(new_n353), .ZN(new_n544));
  XNOR2_X1  g0344(.A(new_n544), .B(KEYINPUT82), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n353), .A2(new_n262), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n543), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(G45), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n548), .A2(G1), .ZN(new_n549));
  INV_X1    g0349(.A(G250), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n274), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT80), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n551), .A2(KEYINPUT80), .A3(new_n274), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n554), .A2(new_n555), .B1(new_n452), .B2(new_n549), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n278), .A2(G244), .A3(G1698), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n278), .A2(G238), .A3(new_n279), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n557), .A2(new_n558), .A3(new_n427), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n317), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n556), .A2(G179), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n297), .B1(new_n556), .B2(new_n560), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n547), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n556), .A2(new_n560), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n292), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n541), .A2(new_n542), .B1(new_n262), .B2(new_n353), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n421), .A2(new_n368), .ZN(new_n567));
  XNOR2_X1  g0367(.A(new_n567), .B(KEYINPUT83), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n556), .A2(G190), .A3(new_n560), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n565), .A2(new_n566), .A3(new_n568), .A4(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n563), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  AND4_X1   g0372(.A1(new_n504), .A2(new_n531), .A3(new_n533), .A4(new_n572), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n416), .A2(new_n480), .A3(new_n573), .ZN(G372));
  NOR2_X1   g0374(.A1(new_n399), .A2(new_n400), .ZN(new_n575));
  INV_X1    g0375(.A(new_n333), .ZN(new_n576));
  INV_X1    g0376(.A(new_n360), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n576), .B1(new_n336), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n575), .B1(new_n578), .B2(new_n393), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n296), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n580), .A2(new_n299), .ZN(new_n581));
  AND4_X1   g0381(.A1(new_n563), .A2(new_n525), .A3(new_n570), .A4(new_n530), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n473), .A2(new_n478), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n504), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n468), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT89), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n526), .B1(new_n297), .B2(new_n513), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n587), .A2(new_n563), .A3(new_n570), .A4(new_n524), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT26), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n586), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n525), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n572), .A2(new_n591), .A3(KEYINPUT89), .A4(KEYINPUT26), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n588), .A2(new_n589), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n590), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n585), .A2(new_n594), .A3(new_n563), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n581), .B1(new_n415), .B2(new_n596), .ZN(G369));
  NAND3_X1  g0397(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n598));
  OR2_X1    g0398(.A1(new_n598), .A2(KEYINPUT27), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(KEYINPUT27), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n599), .A2(G213), .A3(new_n600), .ZN(new_n601));
  XOR2_X1   g0401(.A(KEYINPUT90), .B(G343), .Z(new_n602));
  NOR2_X1   g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n474), .A2(new_n476), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n480), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n603), .ZN(new_n606));
  OR2_X1    g0406(.A1(new_n479), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n504), .A2(new_n533), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n497), .A2(new_n603), .ZN(new_n610));
  MUX2_X1   g0410(.A(new_n504), .B(new_n609), .S(new_n610), .Z(new_n611));
  INV_X1    g0411(.A(G330), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g0414(.A(new_n614), .B(KEYINPUT91), .Z(new_n615));
  NOR2_X1   g0415(.A1(new_n504), .A2(new_n603), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n480), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n473), .A2(new_n478), .A3(new_n606), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OR2_X1    g0419(.A1(new_n615), .A2(new_n619), .ZN(G399));
  INV_X1    g0420(.A(KEYINPUT92), .ZN(new_n621));
  INV_X1    g0421(.A(new_n212), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n621), .B1(new_n622), .B2(G41), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n212), .A2(KEYINPUT92), .A3(new_n273), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(G1), .A3(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n627), .B1(new_n215), .B2(new_n625), .ZN(new_n628));
  XNOR2_X1  g0428(.A(new_n628), .B(KEYINPUT28), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n573), .A2(new_n468), .A3(new_n479), .A4(new_n606), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n449), .A2(new_n458), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n631), .A2(new_n490), .A3(new_n561), .A4(new_n529), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT93), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(KEYINPUT30), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT30), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n632), .A2(new_n633), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(G179), .B1(new_n556), .B2(new_n560), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n499), .A2(new_n459), .A3(new_n513), .A4(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n635), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n603), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT31), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n640), .A2(KEYINPUT31), .A3(new_n603), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n630), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(G330), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n479), .A2(new_n504), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n648), .A2(new_n468), .A3(new_n582), .ZN(new_n649));
  INV_X1    g0449(.A(new_n563), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n572), .A2(KEYINPUT26), .A3(new_n591), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n650), .B1(new_n651), .B2(new_n593), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n603), .B1(new_n649), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT29), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n595), .A2(new_n606), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n656), .A2(KEYINPUT29), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n647), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n629), .B1(new_n658), .B2(G1), .ZN(G364));
  INV_X1    g0459(.A(new_n625), .ZN(new_n660));
  INV_X1    g0460(.A(G13), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n661), .A2(new_n548), .A3(G20), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n662), .A2(KEYINPUT94), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(KEYINPUT94), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(G1), .A3(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n613), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n611), .A2(new_n612), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(G13), .A2(G33), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(G20), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n217), .B1(G20), .B2(new_n297), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n212), .A2(new_n286), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n676), .B1(new_n548), .B2(new_n216), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n248), .B2(new_n548), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n622), .A2(new_n286), .ZN(new_n679));
  INV_X1    g0479(.A(G116), .ZN(new_n680));
  AOI22_X1  g0480(.A1(new_n679), .A2(G355), .B1(new_n680), .B2(new_n622), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n675), .B1(new_n678), .B2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(G283), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n209), .A2(G190), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n292), .A2(new_n358), .A3(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n209), .A2(new_n294), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n292), .A2(new_n358), .A3(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(G303), .ZN(new_n688));
  OAI22_X1  g0488(.A1(new_n683), .A2(new_n685), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(G179), .A2(G200), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT96), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n691), .A2(new_n209), .A3(G190), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n689), .B1(G329), .B2(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n209), .A2(new_n358), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n694), .A2(G190), .A3(G200), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT95), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n695), .A2(new_n696), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(G326), .ZN(new_n701));
  OAI21_X1  g0501(.A(G20), .B1(new_n691), .B2(new_n294), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(G294), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n358), .A2(G200), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n684), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(G311), .ZN(new_n706));
  INV_X1    g0506(.A(G322), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n686), .A2(new_n704), .ZN(new_n708));
  OAI221_X1 g0508(.A(new_n286), .B1(new_n705), .B2(new_n706), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n694), .A2(new_n294), .A3(G200), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  XNOR2_X1  g0511(.A(KEYINPUT33), .B(G317), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n709), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n693), .A2(new_n701), .A3(new_n703), .A4(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n700), .A2(G50), .ZN(new_n715));
  INV_X1    g0515(.A(G58), .ZN(new_n716));
  OAI221_X1 g0516(.A(new_n278), .B1(new_n708), .B2(new_n716), .C1(new_n224), .C2(new_n705), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n717), .B1(G68), .B2(new_n711), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n687), .A2(new_n368), .ZN(new_n719));
  INV_X1    g0519(.A(new_n685), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n719), .B1(G107), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n702), .A2(G97), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n715), .A2(new_n718), .A3(new_n721), .A4(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n692), .A2(G159), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT32), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n714), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n682), .B1(new_n726), .B2(new_n673), .ZN(new_n727));
  INV_X1    g0527(.A(new_n611), .ZN(new_n728));
  INV_X1    g0528(.A(new_n672), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n669), .B1(new_n666), .B2(new_n730), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n731), .B(KEYINPUT97), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(G396));
  AND3_X1   g0533(.A1(new_n357), .A2(new_n359), .A3(new_n606), .ZN(new_n734));
  OR2_X1    g0534(.A1(new_n355), .A2(new_n606), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n356), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n734), .B1(new_n736), .B2(new_n360), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n656), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n595), .A2(new_n606), .A3(new_n737), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n666), .B1(new_n741), .B2(new_n646), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n742), .B1(new_n646), .B2(new_n741), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n673), .A2(new_n670), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n744), .B(KEYINPUT98), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n666), .B1(new_n745), .B2(G77), .ZN(new_n746));
  INV_X1    g0546(.A(new_n708), .ZN(new_n747));
  INV_X1    g0547(.A(new_n705), .ZN(new_n748));
  AOI22_X1  g0548(.A1(G143), .A2(new_n747), .B1(new_n748), .B2(G159), .ZN(new_n749));
  INV_X1    g0549(.A(G137), .ZN(new_n750));
  OAI221_X1 g0550(.A(new_n749), .B1(new_n254), .B2(new_n710), .C1(new_n699), .C2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT34), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n692), .ZN(new_n754));
  INV_X1    g0554(.A(G132), .ZN(new_n755));
  OAI22_X1  g0555(.A1(new_n754), .A2(new_n755), .B1(new_n258), .B2(new_n687), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n685), .A2(new_n222), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n756), .A2(new_n286), .A3(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n702), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n753), .B(new_n758), .C1(new_n716), .C2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n751), .A2(new_n752), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n685), .A2(new_n368), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n762), .B1(G311), .B2(new_n692), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n763), .B1(new_n205), .B2(new_n687), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n700), .A2(G303), .ZN(new_n765));
  INV_X1    g0565(.A(G294), .ZN(new_n766));
  OAI221_X1 g0566(.A(new_n286), .B1(new_n705), .B2(new_n680), .C1(new_n766), .C2(new_n708), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n767), .B1(G283), .B2(new_n711), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n765), .A2(new_n722), .A3(new_n768), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n760), .A2(new_n761), .B1(new_n764), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n746), .B1(new_n770), .B2(new_n673), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(new_n737), .B2(new_n671), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n743), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(G384));
  OR2_X1    g0574(.A1(new_n517), .A2(KEYINPUT35), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n517), .A2(KEYINPUT35), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n775), .A2(G116), .A3(new_n218), .A4(new_n776), .ZN(new_n777));
  XOR2_X1   g0577(.A(new_n777), .B(KEYINPUT36), .Z(new_n778));
  OR3_X1    g0578(.A1(new_n224), .A2(new_n215), .A3(new_n381), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n258), .A2(G68), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n208), .B(G13), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(KEYINPUT38), .ZN(new_n783));
  INV_X1    g0583(.A(new_n601), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT100), .ZN(new_n785));
  AOI21_X1  g0585(.A(KEYINPUT16), .B1(new_n402), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n380), .A2(KEYINPUT100), .A3(new_n386), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n405), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n784), .B1(new_n788), .B2(new_n364), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n401), .A2(new_n413), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n392), .B(KEYINPUT17), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n384), .A2(new_n385), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n255), .A2(G159), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n378), .B1(new_n278), .B2(G20), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n286), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n222), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n785), .B1(new_n795), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n799), .A2(new_n403), .A3(new_n787), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n387), .A2(new_n251), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n364), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n392), .B1(new_n601), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n802), .A2(new_n409), .ZN(new_n804));
  OAI211_X1 g0604(.A(KEYINPUT101), .B(KEYINPUT37), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n394), .A2(new_n397), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n394), .A2(new_n784), .ZN(new_n807));
  XOR2_X1   g0607(.A(KEYINPUT102), .B(KEYINPUT37), .Z(new_n808));
  NAND4_X1  g0608(.A1(new_n806), .A2(new_n807), .A3(new_n392), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n805), .A2(new_n809), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n789), .B(new_n392), .C1(new_n409), .C2(new_n802), .ZN(new_n811));
  AOI21_X1  g0611(.A(KEYINPUT101), .B1(new_n811), .B2(KEYINPUT37), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n783), .B1(new_n792), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(KEYINPUT37), .B1(new_n803), .B2(new_n804), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT101), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n817), .A2(new_n809), .A3(new_n805), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n818), .B(KEYINPUT38), .C1(new_n414), .C2(new_n789), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n814), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(KEYINPUT39), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT39), .ZN(new_n822));
  XOR2_X1   g0622(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n823));
  NAND3_X1  g0623(.A1(new_n806), .A2(new_n807), .A3(new_n392), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(new_n808), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n807), .B1(new_n575), .B2(new_n791), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n823), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n819), .A2(new_n822), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n821), .A2(KEYINPUT104), .A3(new_n828), .ZN(new_n829));
  AOI211_X1 g0629(.A(KEYINPUT104), .B(new_n822), .C1(new_n814), .C2(new_n819), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n576), .A2(new_n606), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n829), .A2(new_n831), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n575), .A2(new_n784), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n820), .ZN(new_n837));
  INV_X1    g0637(.A(new_n734), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n740), .A2(new_n838), .ZN(new_n839));
  AND3_X1   g0639(.A1(new_n310), .A2(new_n311), .A3(new_n603), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT99), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n841), .B1(new_n337), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n333), .A2(new_n842), .A3(new_n336), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n336), .A2(new_n840), .ZN(new_n845));
  INV_X1    g0645(.A(new_n332), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n846), .A2(new_n330), .A3(new_n329), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n844), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n843), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n839), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n836), .B1(new_n837), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(KEYINPUT103), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n850), .B1(new_n740), .B2(new_n838), .ZN(new_n855));
  AOI211_X1 g0655(.A(KEYINPUT103), .B(new_n835), .C1(new_n855), .C2(new_n820), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n834), .A2(new_n854), .A3(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n416), .B1(new_n655), .B2(new_n657), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n859), .A2(new_n581), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n858), .B(new_n860), .Z(new_n861));
  NAND3_X1  g0661(.A1(new_n843), .A2(new_n849), .A3(new_n737), .ZN(new_n862));
  INV_X1    g0662(.A(new_n644), .ZN(new_n863));
  AOI21_X1  g0663(.A(KEYINPUT31), .B1(new_n640), .B2(new_n603), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n862), .B1(new_n630), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(KEYINPUT40), .B1(new_n820), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT106), .ZN(new_n868));
  AND3_X1   g0668(.A1(new_n819), .A2(new_n868), .A3(new_n827), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n868), .B1(new_n819), .B2(new_n827), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AND3_X1   g0671(.A1(new_n843), .A2(new_n849), .A3(new_n737), .ZN(new_n872));
  AND3_X1   g0672(.A1(new_n872), .A2(new_n645), .A3(KEYINPUT40), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n867), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n874), .A2(new_n416), .A3(new_n645), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n874), .B1(new_n416), .B2(new_n645), .ZN(new_n876));
  OR3_X1    g0676(.A1(new_n875), .A2(new_n876), .A3(new_n612), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n861), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(G1), .B1(new_n661), .B2(G20), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n861), .A2(new_n877), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n782), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  XOR2_X1   g0682(.A(new_n882), .B(KEYINPUT107), .Z(G367));
  INV_X1    g0683(.A(new_n615), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n531), .B1(new_n526), .B2(new_n606), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n591), .A2(new_n603), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT42), .B1(new_n617), .B2(new_n888), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT109), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n525), .B1(new_n885), .B2(new_n479), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n892), .A2(KEYINPUT108), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n606), .B1(new_n892), .B2(KEYINPUT108), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n890), .B(new_n891), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  OR3_X1    g0695(.A1(new_n617), .A2(KEYINPUT42), .A3(new_n888), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n566), .A2(new_n568), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n603), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n572), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n563), .B2(new_n899), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n901), .A2(KEYINPUT43), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n890), .B1(new_n893), .B2(new_n894), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(KEYINPUT109), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n897), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n897), .A2(new_n904), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n901), .B(KEYINPUT43), .Z(new_n907));
  AOI22_X1  g0707(.A1(new_n905), .A2(KEYINPUT110), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT110), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n897), .A2(new_n909), .A3(new_n902), .A4(new_n904), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n889), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n905), .A2(KEYINPUT110), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n906), .A2(new_n907), .ZN(new_n913));
  AND4_X1   g0713(.A1(new_n889), .A2(new_n912), .A3(new_n910), .A4(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n625), .B(KEYINPUT41), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT111), .B1(new_n619), .B2(new_n888), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT111), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n617), .A2(new_n918), .A3(new_n618), .A4(new_n887), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT45), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n619), .A2(new_n888), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT44), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n619), .A2(KEYINPUT44), .A3(new_n888), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n924), .A2(KEYINPUT112), .A3(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT112), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n922), .A2(new_n927), .A3(new_n923), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n921), .B(new_n929), .C1(new_n884), .C2(KEYINPUT113), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n920), .A2(KEYINPUT45), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT45), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n917), .B2(new_n919), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n926), .B(new_n928), .C1(new_n931), .C2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT113), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n934), .A2(new_n935), .A3(new_n615), .ZN(new_n936));
  INV_X1    g0736(.A(new_n658), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n617), .B1(new_n608), .B2(new_n616), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(new_n667), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n930), .A2(new_n936), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n916), .B1(new_n941), .B2(new_n658), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n915), .B1(new_n942), .B2(new_n665), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n674), .B1(new_n212), .B2(new_n353), .C1(new_n240), .C2(new_n676), .ZN(new_n944));
  AND2_X1   g0744(.A1(new_n666), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n687), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(G116), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT46), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n947), .A2(new_n948), .B1(G107), .B2(new_n702), .ZN(new_n949));
  OAI221_X1 g0749(.A(new_n949), .B1(new_n948), .B2(new_n947), .C1(new_n706), .C2(new_n699), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n685), .A2(new_n204), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(G317), .B2(new_n692), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n286), .B1(new_n705), .B2(new_n683), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(G303), .B2(new_n747), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n952), .B(new_n954), .C1(new_n766), .C2(new_n710), .ZN(new_n955));
  AOI22_X1  g0755(.A1(G58), .A2(new_n946), .B1(new_n720), .B2(new_n349), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n750), .B2(new_n754), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n278), .B1(new_n705), .B2(new_n258), .C1(new_n254), .C2(new_n708), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(G159), .B2(new_n711), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n702), .A2(G68), .ZN(new_n960));
  INV_X1    g0760(.A(G143), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n959), .B(new_n960), .C1(new_n961), .C2(new_n699), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n950), .A2(new_n955), .B1(new_n957), .B2(new_n962), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n963), .B(KEYINPUT47), .Z(new_n964));
  INV_X1    g0764(.A(new_n673), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n945), .B1(new_n901), .B2(new_n729), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n943), .A2(new_n966), .ZN(G387));
  INV_X1    g0767(.A(new_n940), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n937), .A2(new_n939), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n968), .A2(new_n969), .A3(new_n660), .ZN(new_n970));
  INV_X1    g0770(.A(new_n626), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n679), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(G107), .B2(new_n212), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n237), .A2(new_n548), .ZN(new_n974));
  AOI211_X1 g0774(.A(G45), .B(new_n971), .C1(G68), .C2(G77), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n252), .A2(G50), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT50), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n676), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n973), .B1(new_n974), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n666), .B1(new_n979), .B2(new_n675), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n687), .A2(new_n224), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n951), .B(new_n981), .C1(G150), .C2(new_n692), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n759), .A2(new_n353), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n700), .A2(G159), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n278), .B1(new_n705), .B2(new_n222), .C1(new_n258), .C2(new_n708), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(new_n351), .B2(new_n711), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n982), .A2(new_n983), .A3(new_n984), .A4(new_n986), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n759), .A2(new_n683), .B1(new_n766), .B2(new_n687), .ZN(new_n988));
  AOI22_X1  g0788(.A1(G317), .A2(new_n747), .B1(new_n748), .B2(G303), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n706), .B2(new_n710), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(G322), .B2(new_n700), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n988), .B1(new_n991), .B2(KEYINPUT48), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT114), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(KEYINPUT48), .B2(new_n991), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT49), .Z(new_n995));
  AOI21_X1  g0795(.A(new_n278), .B1(new_n692), .B2(G326), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n680), .B2(new_n685), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n987), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n980), .B1(new_n998), .B2(new_n673), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n605), .A2(new_n607), .A3(new_n672), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n665), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n970), .B(new_n1001), .C1(new_n1002), .C2(new_n939), .ZN(G393));
  NOR2_X1   g0803(.A1(new_n934), .A2(new_n615), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n884), .B1(new_n921), .B2(new_n929), .ZN(new_n1005));
  OAI21_X1  g0805(.A(KEYINPUT115), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n934), .A2(new_n615), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n921), .A2(new_n884), .A3(new_n929), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT115), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1006), .A2(new_n665), .A3(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n968), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1012), .A2(new_n941), .A3(new_n660), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n245), .A2(new_n676), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n674), .B1(new_n204), .B2(new_n212), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n666), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(G159), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n699), .A2(new_n254), .B1(new_n1017), .B2(new_n708), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT51), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n702), .A2(G77), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n754), .A2(new_n961), .B1(new_n222), .B2(new_n687), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n278), .B1(new_n705), .B2(new_n252), .C1(new_n710), .C2(new_n258), .ZN(new_n1022));
  NOR3_X1   g0822(.A1(new_n1021), .A2(new_n762), .A3(new_n1022), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1019), .A2(new_n1020), .A3(new_n1023), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n700), .A2(G317), .B1(G311), .B2(new_n747), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT116), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(KEYINPUT52), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n278), .B1(new_n748), .B2(G294), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n688), .B2(new_n710), .C1(new_n205), .C2(new_n685), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n754), .A2(new_n707), .B1(new_n683), .B2(new_n687), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n1029), .B(new_n1030), .C1(G116), .C2(new_n702), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1027), .A2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1026), .A2(KEYINPUT52), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1024), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1016), .B1(new_n1034), .B2(new_n673), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n729), .B2(new_n887), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1011), .A2(new_n1013), .A3(new_n1036), .ZN(G390));
  NAND3_X1  g0837(.A1(new_n647), .A2(new_n737), .A3(new_n851), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n855), .A2(new_n833), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n829), .B2(new_n831), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n819), .A2(new_n827), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(KEYINPUT106), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n819), .A2(new_n868), .A3(new_n827), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n736), .A2(new_n360), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n734), .B1(new_n653), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n832), .B1(new_n1047), .B2(new_n850), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1039), .B1(new_n1041), .B2(new_n1049), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT104), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n820), .B2(KEYINPUT39), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n830), .B1(new_n1053), .B2(new_n828), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1051), .B(new_n1038), .C1(new_n1054), .C2(new_n1040), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1050), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n647), .A2(new_n416), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n859), .A2(new_n1057), .A3(new_n581), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n850), .B1(new_n646), .B2(new_n738), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1038), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n839), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1038), .A2(new_n1047), .A3(new_n1059), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1058), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n625), .B1(new_n1056), .B2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1050), .A2(new_n1055), .A3(new_n1063), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n666), .B1(new_n745), .B2(new_n351), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n719), .B(new_n757), .C1(G294), .C2(new_n692), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n700), .A2(G283), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n286), .B1(new_n705), .B2(new_n204), .C1(new_n680), .C2(new_n708), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(G107), .B2(new_n711), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1069), .A2(new_n1020), .A3(new_n1070), .A4(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(KEYINPUT54), .B(G143), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(G132), .A2(new_n747), .B1(new_n748), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n750), .B2(new_n710), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(G125), .B2(new_n692), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n278), .B1(new_n685), .B2(new_n258), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(KEYINPUT117), .ZN(new_n1080));
  OR2_X1    g0880(.A1(new_n1079), .A2(KEYINPUT117), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n700), .A2(G128), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1078), .A2(new_n1080), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  OR3_X1    g0883(.A1(new_n687), .A2(KEYINPUT53), .A3(new_n254), .ZN(new_n1084));
  OAI21_X1  g0884(.A(KEYINPUT53), .B1(new_n687), .B2(new_n254), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1084), .B(new_n1085), .C1(new_n759), .C2(new_n1017), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1073), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1068), .B1(new_n1087), .B2(new_n673), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n1054), .B2(new_n671), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n1056), .B2(new_n1002), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n1067), .A2(new_n1090), .ZN(G378));
  NAND2_X1  g0891(.A1(new_n268), .A2(new_n784), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n300), .B(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1093), .B(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n874), .B2(G330), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n820), .A2(new_n866), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT40), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1043), .A2(new_n1044), .A3(new_n873), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1095), .A2(new_n1099), .A3(new_n1100), .A4(G330), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n858), .B1(new_n1096), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n856), .B1(new_n1054), .B2(new_n833), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1099), .A2(new_n1100), .A3(G330), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1095), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1104), .A2(new_n1107), .A3(new_n854), .A4(new_n1101), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1103), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1106), .A2(new_n670), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n744), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n666), .B1(G50), .B2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n278), .A2(G41), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1113), .B1(new_n353), .B2(new_n705), .C1(new_n205), .C2(new_n708), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(G97), .B2(new_n711), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n685), .A2(new_n716), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n981), .B(new_n1116), .C1(G283), .C2(new_n692), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n960), .B1(new_n699), .B2(new_n680), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n1118), .A2(KEYINPUT118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1118), .A2(KEYINPUT118), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1115), .B(new_n1117), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1121));
  XOR2_X1   g0921(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1113), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1124), .B(new_n258), .C1(G33), .C2(G41), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(G128), .A2(new_n747), .B1(new_n748), .B2(G137), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n755), .B2(new_n710), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(new_n946), .B2(new_n1075), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n700), .A2(G125), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1129), .B(new_n1130), .C1(new_n254), .C2(new_n759), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1131), .A2(KEYINPUT59), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(KEYINPUT59), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n720), .A2(G159), .ZN(new_n1134));
  AOI211_X1 g0934(.A(G33), .B(G41), .C1(new_n692), .C2(G124), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n1126), .B1(new_n1122), .B2(new_n1121), .C1(new_n1132), .C2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1112), .B1(new_n1137), .B2(new_n673), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n1109), .A2(new_n665), .B1(new_n1110), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT57), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n1103), .B2(new_n1108), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1058), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1066), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1144), .A2(KEYINPUT120), .A3(new_n660), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1143), .A2(new_n1109), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n1140), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(KEYINPUT120), .B1(new_n1144), .B2(new_n660), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1139), .B1(new_n1148), .B2(new_n1149), .ZN(G375));
  NAND3_X1  g0950(.A1(new_n1061), .A2(new_n1058), .A3(new_n1062), .ZN(new_n1151));
  OR2_X1    g0951(.A1(new_n1151), .A2(KEYINPUT121), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(KEYINPUT121), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1063), .A2(new_n916), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n665), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n666), .B1(new_n745), .B2(G68), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n687), .A2(new_n1017), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n1116), .B(new_n1159), .C1(G128), .C2(new_n692), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n700), .A2(G132), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n702), .A2(G50), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n278), .B1(new_n705), .B2(new_n254), .C1(new_n750), .C2(new_n708), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n711), .B2(new_n1075), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .A4(new_n1164), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(G283), .A2(new_n747), .B1(new_n748), .B2(G107), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n680), .B2(new_n710), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(G97), .B2(new_n946), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n692), .A2(G303), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n700), .A2(G294), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1168), .A2(new_n983), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n286), .B1(new_n685), .B2(new_n304), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT122), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1165), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT123), .ZN(new_n1175));
  OR2_X1    g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n965), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1158), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n851), .B2(new_n671), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1157), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1155), .A2(new_n1181), .ZN(G381));
  OR3_X1    g0982(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1183));
  NOR4_X1   g0983(.A1(G387), .A2(new_n1183), .A3(G390), .A4(G381), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1184), .B(KEYINPUT124), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(G375), .A2(G378), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(G407));
  NAND2_X1  g0987(.A1(new_n602), .A2(G213), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1186), .A2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(G407), .A2(G213), .A3(new_n1190), .ZN(G409));
  OAI211_X1 g0991(.A(G378), .B(new_n1139), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1067), .A2(new_n1090), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1139), .B1(new_n1146), .B2(new_n916), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1189), .B1(new_n1192), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1064), .A2(KEYINPUT60), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1197), .A2(new_n1153), .A3(new_n1152), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1151), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n625), .B1(new_n1199), .B2(KEYINPUT60), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(G384), .B1(new_n1201), .B2(new_n1181), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n773), .B(new_n1180), .C1(new_n1198), .C2(new_n1200), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1196), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT63), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1189), .A2(G2897), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1204), .A2(new_n1208), .ZN(new_n1209));
  OAI211_X1 g1009(.A(G2897), .B(new_n1189), .C1(new_n1202), .C2(new_n1203), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  OR2_X1    g1011(.A1(new_n1196), .A2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1196), .A2(KEYINPUT63), .A3(new_n1204), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n943), .A2(G390), .A3(new_n966), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(G390), .B1(new_n943), .B2(new_n966), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(G393), .B(new_n732), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NOR3_X1   g1018(.A1(new_n1215), .A2(new_n1216), .A3(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(G390), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(G387), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1217), .B1(new_n1221), .B2(new_n1214), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(new_n1219), .A2(new_n1222), .A3(KEYINPUT61), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1207), .A2(new_n1212), .A3(new_n1213), .A4(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT62), .ZN(new_n1225));
  AND3_X1   g1025(.A1(new_n1196), .A2(new_n1225), .A3(new_n1204), .ZN(new_n1226));
  XOR2_X1   g1026(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n1196), .B2(new_n1211), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1225), .B1(new_n1196), .B2(new_n1204), .ZN(new_n1229));
  NOR3_X1   g1029(.A1(new_n1226), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT126), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n1219), .B2(new_n1222), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1218), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1221), .A2(new_n1217), .A3(new_n1214), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1233), .A2(new_n1234), .A3(KEYINPUT126), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1232), .A2(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1224), .B1(new_n1230), .B2(new_n1236), .ZN(G405));
  NOR2_X1   g1037(.A1(new_n1204), .A2(KEYINPUT127), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  AND3_X1   g1039(.A1(new_n1232), .A2(new_n1235), .A3(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1239), .B1(new_n1232), .B2(new_n1235), .ZN(new_n1241));
  AND2_X1   g1041(.A1(G375), .A2(new_n1193), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1204), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT127), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1192), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n1240), .A2(new_n1241), .B1(new_n1242), .B2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1236), .A2(new_n1238), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1245), .A2(new_n1242), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1232), .A2(new_n1235), .A3(new_n1239), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1247), .A2(new_n1248), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1246), .A2(new_n1250), .ZN(G402));
endmodule


