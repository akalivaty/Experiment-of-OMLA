//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 0 0 1 0 1 1 1 0 1 0 1 1 0 1 0 0 0 1 1 0 0 1 1 1 1 1 0 1 0 1 1 1 1 0 0 0 1 0 0 0 1 0 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n780,
    new_n781, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT23), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G128), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT23), .A3(G119), .ZN(new_n192));
  OAI211_X1 g006(.A(new_n190), .B(new_n192), .C1(G119), .C2(new_n191), .ZN(new_n193));
  XNOR2_X1  g007(.A(G119), .B(G128), .ZN(new_n194));
  XOR2_X1   g008(.A(KEYINPUT24), .B(G110), .Z(new_n195));
  AOI22_X1  g009(.A1(new_n193), .A2(G110), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G140), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G125), .ZN(new_n198));
  INV_X1    g012(.A(G125), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G140), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n198), .A2(new_n200), .A3(KEYINPUT16), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n199), .A2(G140), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT16), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  AND3_X1   g018(.A1(new_n201), .A2(G146), .A3(new_n204), .ZN(new_n205));
  AOI21_X1  g019(.A(G146), .B1(new_n201), .B2(new_n204), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n196), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  OAI22_X1  g021(.A1(new_n193), .A2(G110), .B1(new_n194), .B2(new_n195), .ZN(new_n208));
  NOR3_X1   g022(.A1(new_n199), .A2(KEYINPUT16), .A3(G140), .ZN(new_n209));
  XNOR2_X1  g023(.A(G125), .B(G140), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n209), .B1(new_n210), .B2(KEYINPUT16), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G146), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n198), .A2(new_n200), .A3(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n208), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n207), .A2(new_n215), .A3(KEYINPUT73), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT22), .B(G137), .ZN(new_n217));
  INV_X1    g031(.A(G953), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(G221), .A3(G234), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n217), .B(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n216), .A2(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(KEYINPUT73), .B1(new_n207), .B2(new_n215), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n207), .A2(new_n215), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT73), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n226), .A3(new_n220), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n187), .B1(new_n224), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT25), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n225), .A2(new_n226), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(new_n216), .A3(new_n221), .ZN(new_n232));
  AOI21_X1  g046(.A(G902), .B1(new_n232), .B2(new_n227), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT25), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G217), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n236), .B1(G234), .B2(new_n187), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n230), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n232), .A2(new_n227), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n237), .A2(G902), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n242), .B(KEYINPUT74), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n239), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  OR2_X1    g059(.A1(KEYINPUT67), .A2(G137), .ZN(new_n246));
  NAND2_X1  g060(.A1(KEYINPUT67), .A2(G137), .ZN(new_n247));
  AOI21_X1  g061(.A(G134), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G137), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G134), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(G131), .B1(new_n248), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT11), .ZN(new_n253));
  INV_X1    g067(.A(G134), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n255), .A2(new_n246), .A3(new_n247), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(G137), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT66), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n258), .B1(new_n250), .B2(new_n253), .ZN(new_n259));
  AOI211_X1 g073(.A(KEYINPUT66), .B(KEYINPUT11), .C1(new_n249), .C2(G134), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n256), .B(new_n257), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n252), .B1(new_n261), .B2(G131), .ZN(new_n262));
  INV_X1    g076(.A(G143), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT1), .B1(new_n263), .B2(G146), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT68), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n213), .A2(G143), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT68), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(new_n267), .A3(KEYINPUT1), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n265), .A2(G128), .A3(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT64), .B1(new_n263), .B2(G146), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT64), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(new_n213), .A3(G143), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n213), .A2(G143), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n263), .A2(G146), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT65), .B1(new_n213), .B2(G143), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT65), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n279), .A2(new_n263), .A3(G146), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n277), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n191), .A2(KEYINPUT1), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n269), .A2(new_n276), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n262), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n279), .B1(new_n263), .B2(G146), .ZN(new_n285));
  NOR3_X1   g099(.A1(new_n213), .A2(KEYINPUT65), .A3(G143), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n266), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(KEYINPUT0), .A2(G128), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n274), .B1(new_n270), .B2(new_n272), .ZN(new_n289));
  INV_X1    g103(.A(new_n288), .ZN(new_n290));
  NOR2_X1   g104(.A1(KEYINPUT0), .A2(G128), .ZN(new_n291));
  OR2_X1    g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI22_X1  g106(.A1(new_n287), .A2(new_n288), .B1(new_n289), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n261), .A2(G131), .ZN(new_n294));
  AND2_X1   g108(.A1(KEYINPUT67), .A2(G137), .ZN(new_n295));
  NOR2_X1   g109(.A1(KEYINPUT67), .A2(G137), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n297), .A2(new_n255), .B1(new_n254), .B2(G137), .ZN(new_n298));
  INV_X1    g112(.A(G131), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n253), .B1(new_n254), .B2(G137), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT66), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n250), .A2(new_n258), .A3(new_n253), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n298), .A2(new_n299), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n293), .B1(new_n294), .B2(new_n304), .ZN(new_n305));
  OAI211_X1 g119(.A(KEYINPUT70), .B(KEYINPUT30), .C1(new_n284), .C2(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n290), .A2(new_n291), .ZN(new_n307));
  AOI22_X1  g121(.A1(new_n276), .A2(new_n307), .B1(new_n281), .B2(new_n290), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n261), .A2(G131), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n299), .B1(new_n298), .B2(new_n303), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT1), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n312), .B1(G143), .B2(new_n213), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n191), .B1(new_n313), .B2(new_n267), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n289), .B1(new_n314), .B2(new_n265), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n266), .B(new_n282), .C1(new_n285), .C2(new_n286), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n304), .B(new_n252), .C1(new_n315), .C2(new_n317), .ZN(new_n318));
  OR2_X1    g132(.A1(KEYINPUT70), .A2(KEYINPUT30), .ZN(new_n319));
  NAND2_X1  g133(.A1(KEYINPUT70), .A2(KEYINPUT30), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n311), .A2(new_n318), .A3(new_n319), .A4(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n306), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n189), .A2(G116), .ZN(new_n323));
  INV_X1    g137(.A(G116), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G119), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT69), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT69), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n323), .A2(new_n325), .A3(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT2), .B(G113), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n327), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  OR2_X1    g145(.A1(new_n326), .A2(new_n330), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n322), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT31), .ZN(new_n335));
  INV_X1    g149(.A(new_n333), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n311), .A2(new_n336), .A3(new_n318), .ZN(new_n337));
  NOR2_X1   g151(.A1(G237), .A2(G953), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G210), .ZN(new_n339));
  XOR2_X1   g153(.A(new_n339), .B(KEYINPUT27), .Z(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT26), .B(G101), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n340), .B(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n334), .A2(new_n335), .A3(new_n337), .A4(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT71), .ZN(new_n345));
  NOR3_X1   g159(.A1(new_n284), .A2(new_n305), .A3(new_n333), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n346), .B1(new_n322), .B2(new_n333), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT71), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n347), .A2(new_n348), .A3(new_n335), .A4(new_n343), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n336), .B1(new_n311), .B2(new_n318), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT28), .B1(new_n346), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT28), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n337), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(KEYINPUT72), .B1(new_n355), .B2(new_n342), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n333), .B1(new_n284), .B2(new_n305), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n353), .B1(new_n357), .B2(new_n337), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n337), .A2(new_n353), .ZN(new_n359));
  OAI211_X1 g173(.A(KEYINPUT72), .B(new_n342), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n356), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n347), .A2(new_n343), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT31), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n350), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(G472), .A2(G902), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT32), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n366), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n370), .A2(new_n368), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT29), .ZN(new_n372));
  AOI211_X1 g186(.A(new_n346), .B(new_n343), .C1(new_n322), .C2(new_n333), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n342), .B1(new_n352), .B2(new_n354), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n355), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n342), .A2(new_n372), .ZN(new_n377));
  AOI21_X1  g191(.A(G902), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  AOI22_X1  g193(.A1(new_n365), .A2(new_n371), .B1(G472), .B2(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n245), .B1(new_n369), .B2(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n197), .A2(G125), .ZN(new_n382));
  OAI21_X1  g196(.A(G146), .B1(new_n202), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n214), .ZN(new_n384));
  NAND2_X1  g198(.A1(KEYINPUT18), .A2(G131), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G237), .ZN(new_n387));
  AND4_X1   g201(.A1(G143), .A2(new_n387), .A3(new_n218), .A4(G214), .ZN(new_n388));
  AOI21_X1  g202(.A(G143), .B1(new_n338), .B2(G214), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n386), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n387), .A2(new_n218), .A3(G214), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n263), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n338), .A2(G143), .A3(G214), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n393), .A3(new_n385), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n384), .A2(new_n390), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(KEYINPUT84), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT84), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n384), .A2(new_n390), .A3(new_n397), .A4(new_n394), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n205), .A2(new_n206), .ZN(new_n400));
  OAI211_X1 g214(.A(KEYINPUT17), .B(G131), .C1(new_n388), .C2(new_n389), .ZN(new_n401));
  OAI21_X1  g215(.A(G131), .B1(new_n388), .B2(new_n389), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n392), .A2(new_n299), .A3(new_n393), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n400), .B(new_n401), .C1(KEYINPUT17), .C2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n399), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(G113), .B(G122), .ZN(new_n407));
  INV_X1    g221(.A(G104), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n407), .B(new_n408), .ZN(new_n409));
  XOR2_X1   g223(.A(new_n409), .B(KEYINPUT88), .Z(new_n410));
  NOR2_X1   g224(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT87), .ZN(new_n412));
  AOI22_X1  g226(.A1(new_n402), .A2(new_n403), .B1(new_n211), .B2(G146), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT85), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n210), .A2(new_n414), .A3(KEYINPUT19), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT19), .B1(new_n210), .B2(new_n414), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n213), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n388), .A2(new_n389), .ZN(new_n419));
  AOI22_X1  g233(.A1(new_n419), .A2(new_n385), .B1(new_n214), .B2(new_n383), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n397), .B1(new_n420), .B2(new_n390), .ZN(new_n421));
  INV_X1    g235(.A(new_n398), .ZN(new_n422));
  OAI211_X1 g236(.A(KEYINPUT86), .B(new_n418), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n409), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(KEYINPUT86), .B1(new_n399), .B2(new_n418), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n412), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI22_X1  g241(.A1(new_n396), .A2(new_n398), .B1(new_n417), .B2(new_n413), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n409), .B1(new_n428), .B2(KEYINPUT86), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n418), .B1(new_n421), .B2(new_n422), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT86), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n429), .A2(KEYINPUT87), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n411), .B1(new_n427), .B2(new_n433), .ZN(new_n434));
  NOR2_X1   g248(.A1(G475), .A2(G902), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(KEYINPUT20), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n411), .ZN(new_n438));
  NOR3_X1   g252(.A1(new_n425), .A2(new_n412), .A3(new_n426), .ZN(new_n439));
  AOI21_X1  g253(.A(KEYINPUT87), .B1(new_n429), .B2(new_n432), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT20), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n441), .A2(new_n442), .A3(new_n435), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n437), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n406), .A2(new_n424), .ZN(new_n445));
  AOI21_X1  g259(.A(G902), .B1(new_n438), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(G475), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n444), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(KEYINPUT89), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT91), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n324), .A2(G122), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n324), .A2(G122), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n452), .B(new_n453), .C1(new_n454), .C2(KEYINPUT14), .ZN(new_n455));
  INV_X1    g269(.A(new_n453), .ZN(new_n456));
  INV_X1    g270(.A(new_n454), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT14), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(KEYINPUT91), .B1(new_n453), .B2(KEYINPUT14), .ZN(new_n460));
  OAI211_X1 g274(.A(G107), .B(new_n455), .C1(new_n459), .C2(new_n460), .ZN(new_n461));
  NOR3_X1   g275(.A1(new_n456), .A2(G107), .A3(new_n454), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n191), .A2(G143), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n263), .A2(G128), .ZN(new_n464));
  OR3_X1    g278(.A1(new_n463), .A2(new_n464), .A3(G134), .ZN(new_n465));
  OAI21_X1  g279(.A(G134), .B1(new_n463), .B2(new_n464), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n461), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(KEYINPUT13), .B1(new_n263), .B2(G128), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n469), .B1(new_n191), .B2(G143), .ZN(new_n470));
  OR2_X1    g284(.A1(new_n470), .A2(KEYINPUT90), .ZN(new_n471));
  AOI22_X1  g285(.A1(new_n470), .A2(KEYINPUT90), .B1(KEYINPUT13), .B2(new_n463), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n254), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(G107), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n474), .B1(new_n457), .B2(new_n453), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n465), .B1(new_n475), .B2(new_n462), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n468), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(KEYINPUT9), .B(G234), .ZN(new_n478));
  NOR3_X1   g292(.A1(new_n478), .A2(new_n236), .A3(G953), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n468), .B(new_n479), .C1(new_n473), .C2(new_n476), .ZN(new_n482));
  AOI21_X1  g296(.A(G902), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  XOR2_X1   g297(.A(new_n483), .B(KEYINPUT92), .Z(new_n484));
  INV_X1    g298(.A(G478), .ZN(new_n485));
  AOI211_X1 g299(.A(KEYINPUT15), .B(new_n485), .C1(new_n483), .C2(KEYINPUT93), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n485), .A2(KEYINPUT15), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT93), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n488), .B1(new_n483), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(G234), .A2(G237), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n493), .A2(G952), .A3(new_n218), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n493), .A2(G902), .A3(G953), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  XOR2_X1   g311(.A(KEYINPUT21), .B(G898), .Z(new_n498));
  OAI21_X1  g312(.A(new_n495), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n492), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT89), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n444), .A2(new_n501), .A3(new_n449), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n451), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(G214), .B1(G237), .B2(G902), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(G110), .B(G122), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT5), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n507), .B1(new_n327), .B2(new_n329), .ZN(new_n508));
  OAI21_X1  g322(.A(G113), .B1(new_n323), .B2(KEYINPUT5), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n332), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT3), .ZN(new_n511));
  NOR3_X1   g325(.A1(new_n408), .A2(KEYINPUT77), .A3(G107), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n511), .B1(new_n512), .B2(KEYINPUT76), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n474), .A2(KEYINPUT76), .A3(G104), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n408), .A2(G107), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(G101), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT76), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n474), .A2(G104), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n519), .B(KEYINPUT3), .C1(new_n520), .C2(KEYINPUT77), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n513), .A2(new_n517), .A3(new_n518), .A4(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n515), .A2(new_n520), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G101), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n522), .A2(KEYINPUT4), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n519), .B1(new_n520), .B2(KEYINPUT77), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n516), .B1(new_n527), .B2(new_n511), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n518), .B1(new_n528), .B2(new_n521), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n513), .A2(new_n517), .A3(new_n521), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT4), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n532), .A3(G101), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n333), .ZN(new_n534));
  OAI221_X1 g348(.A(new_n506), .B1(new_n510), .B2(new_n525), .C1(new_n530), .C2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT80), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n536), .B1(new_n308), .B2(new_n199), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n283), .A2(new_n199), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n293), .A2(KEYINPUT80), .A3(G125), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n218), .A2(G224), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(KEYINPUT7), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n537), .A2(new_n538), .A3(new_n539), .A4(new_n542), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n522), .A2(new_n524), .ZN(new_n544));
  OAI22_X1  g358(.A1(new_n509), .A2(KEYINPUT82), .B1(new_n326), .B2(new_n507), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n509), .A2(KEYINPUT82), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n332), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n506), .B(KEYINPUT8), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n548), .B(new_n549), .C1(new_n544), .C2(new_n510), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n535), .A2(new_n543), .A3(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n537), .A2(new_n539), .A3(new_n538), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n552), .A2(KEYINPUT83), .A3(new_n541), .ZN(new_n553));
  AOI21_X1  g367(.A(KEYINPUT83), .B1(new_n552), .B2(new_n541), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(G902), .B1(new_n551), .B2(new_n555), .ZN(new_n556));
  OAI22_X1  g370(.A1(new_n530), .A2(new_n534), .B1(new_n525), .B2(new_n510), .ZN(new_n557));
  INV_X1    g371(.A(new_n506), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n559), .A2(KEYINPUT6), .A3(new_n535), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n540), .B(KEYINPUT81), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n552), .B(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT6), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n557), .A2(new_n563), .A3(new_n558), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n560), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n556), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(G210), .B1(G237), .B2(G902), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n556), .A2(new_n567), .A3(new_n565), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n505), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(G221), .B1(new_n478), .B2(G902), .ZN(new_n572));
  XOR2_X1   g386(.A(new_n572), .B(KEYINPUT75), .Z(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(G469), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT78), .ZN(new_n576));
  OAI21_X1  g390(.A(KEYINPUT10), .B1(new_n315), .B2(new_n317), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n576), .B1(new_n577), .B2(new_n525), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT10), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n269), .A2(new_n276), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n579), .B1(new_n580), .B2(new_n316), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n544), .A2(new_n581), .A3(KEYINPUT78), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n293), .B1(new_n529), .B2(new_n532), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n531), .A2(G101), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n585), .A2(KEYINPUT4), .A3(new_n522), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n313), .A2(new_n191), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n316), .B1(new_n281), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n588), .A2(new_n524), .A3(new_n522), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n584), .A2(new_n586), .B1(new_n579), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n309), .A2(new_n310), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n583), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n525), .A2(new_n283), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n589), .ZN(new_n594));
  INV_X1    g408(.A(new_n591), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(KEYINPUT12), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT12), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n594), .A2(new_n595), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n592), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(G110), .B(G140), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n218), .A2(G227), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n583), .A2(new_n590), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n595), .ZN(new_n606));
  INV_X1    g420(.A(new_n603), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n606), .A2(new_n592), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(KEYINPUT79), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT79), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n604), .A2(new_n611), .A3(new_n608), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n575), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n607), .B1(new_n606), .B2(new_n592), .ZN(new_n614));
  AND4_X1   g428(.A1(new_n592), .A2(new_n607), .A3(new_n597), .A4(new_n599), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n575), .B(new_n187), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n575), .A2(new_n187), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n571), .B(new_n574), .C1(new_n613), .C2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n381), .A2(new_n503), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(G101), .ZN(G3));
  NOR2_X1   g437(.A1(new_n484), .A2(G478), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n481), .A2(new_n482), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(KEYINPUT33), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n485), .A2(G902), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n624), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n628), .B1(new_n451), .B2(new_n502), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n244), .B(new_n574), .C1(new_n613), .C2(new_n619), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n335), .B1(new_n347), .B2(new_n343), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n356), .A2(new_n632), .A3(new_n361), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n370), .B1(new_n633), .B2(new_n350), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n365), .A2(new_n187), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n634), .B1(new_n635), .B2(G472), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n556), .A2(new_n567), .A3(new_n565), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n567), .B1(new_n556), .B2(new_n565), .ZN(new_n638));
  OAI211_X1 g452(.A(new_n499), .B(new_n504), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n629), .A2(new_n631), .A3(new_n636), .A4(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT34), .B(G104), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G6));
  NAND2_X1  g457(.A1(new_n448), .A2(KEYINPUT94), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT94), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n645), .B1(new_n446), .B2(new_n447), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n490), .B1(new_n484), .B2(new_n486), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n444), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n631), .A2(new_n636), .A3(new_n640), .A4(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT35), .B(G107), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G9));
  NOR2_X1   g467(.A1(new_n221), .A2(KEYINPUT36), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n225), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n241), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n238), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n503), .A2(new_n621), .A3(new_n636), .A4(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT37), .B(G110), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G12));
  AND2_X1   g474(.A1(new_n345), .A2(new_n349), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n342), .B1(new_n358), .B2(new_n359), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT72), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n364), .A2(new_n360), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n371), .B1(new_n661), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n379), .A2(G472), .ZN(new_n667));
  OAI211_X1 g481(.A(new_n666), .B(new_n667), .C1(new_n634), .C2(KEYINPUT32), .ZN(new_n668));
  OR2_X1    g482(.A1(new_n497), .A2(G900), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n495), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n649), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n621), .A2(new_n668), .A3(new_n657), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  XNOR2_X1  g488(.A(new_n670), .B(KEYINPUT39), .ZN(new_n675));
  OAI211_X1 g489(.A(new_n574), .B(new_n675), .C1(new_n613), .C2(new_n619), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT40), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT98), .ZN(new_n678));
  OR2_X1    g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n501), .B1(new_n444), .B2(new_n449), .ZN(new_n681));
  AOI211_X1 g495(.A(KEYINPUT89), .B(new_n448), .C1(new_n437), .C2(new_n443), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n648), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(G472), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n187), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n347), .A2(new_n343), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n343), .B1(new_n357), .B2(new_n337), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n685), .B1(new_n689), .B2(KEYINPUT96), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n342), .B1(new_n346), .B2(new_n351), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT96), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n687), .B1(new_n688), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(KEYINPUT97), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT97), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n697), .B(new_n687), .C1(new_n688), .C2(new_n694), .ZN(new_n698));
  AOI22_X1  g512(.A1(new_n365), .A2(new_n371), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n369), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n569), .A2(new_n570), .ZN(new_n701));
  XOR2_X1   g515(.A(KEYINPUT95), .B(KEYINPUT38), .Z(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NOR4_X1   g517(.A1(new_n700), .A2(new_n505), .A3(new_n703), .A4(new_n657), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n679), .A2(new_n680), .A3(new_n684), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G143), .ZN(G45));
  AOI211_X1 g520(.A(new_n671), .B(new_n628), .C1(new_n451), .C2(new_n502), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n707), .A2(new_n668), .A3(new_n621), .A4(new_n657), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G146), .ZN(G48));
  NAND2_X1  g523(.A1(new_n451), .A2(new_n502), .ZN(new_n710));
  INV_X1    g524(.A(new_n628), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n710), .A2(new_n711), .A3(new_n640), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n187), .B1(new_n614), .B2(new_n615), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(G469), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(new_n574), .A3(new_n616), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n666), .A2(new_n667), .ZN(new_n717));
  AOI21_X1  g531(.A(KEYINPUT32), .B1(new_n365), .B2(new_n366), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n244), .B(new_n716), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n712), .A2(new_n719), .ZN(new_n720));
  XOR2_X1   g534(.A(KEYINPUT41), .B(G113), .Z(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G15));
  NOR2_X1   g536(.A1(new_n649), .A2(new_n639), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n668), .A2(new_n244), .A3(new_n716), .A4(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(KEYINPUT99), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT99), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n381), .A2(new_n726), .A3(new_n716), .A4(new_n723), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G116), .ZN(G18));
  NAND2_X1  g543(.A1(new_n668), .A2(new_n657), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n504), .B1(new_n637), .B2(new_n638), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n715), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n732), .A2(new_n502), .A3(new_n451), .A4(new_n500), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(new_n189), .ZN(G21));
  INV_X1    g549(.A(KEYINPUT100), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n355), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n352), .A2(KEYINPUT100), .A3(new_n354), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n342), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n364), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n366), .B1(new_n661), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(G902), .B1(new_n633), .B2(new_n350), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n741), .B(new_n244), .C1(new_n742), .C2(new_n685), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n714), .A2(new_n616), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n744), .A2(new_n499), .A3(new_n571), .A4(new_n574), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n683), .A2(KEYINPUT101), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT101), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n748), .B(new_n648), .C1(new_n681), .C2(new_n682), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n746), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(KEYINPUT102), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT102), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n746), .A2(new_n747), .A3(new_n752), .A4(new_n749), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G122), .ZN(G24));
  INV_X1    g569(.A(new_n732), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n741), .B(new_n657), .C1(new_n742), .C2(new_n685), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT103), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(new_n707), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n635), .A2(G472), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n761), .A2(new_n732), .A3(new_n657), .A4(new_n741), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n711), .B(new_n670), .C1(new_n681), .C2(new_n682), .ZN(new_n763));
  OAI21_X1  g577(.A(KEYINPUT103), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G125), .ZN(G27));
  NOR3_X1   g580(.A1(new_n637), .A2(new_n638), .A3(new_n505), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n608), .A2(KEYINPUT104), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT104), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n606), .A2(new_n769), .A3(new_n592), .A4(new_n607), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n768), .A2(G469), .A3(new_n604), .A4(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n616), .A3(new_n618), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n767), .A2(new_n574), .A3(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n707), .A2(new_n381), .A3(KEYINPUT42), .A4(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT42), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n668), .A2(new_n773), .A3(new_n244), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n775), .B1(new_n776), .B2(new_n763), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G131), .ZN(G33));
  INV_X1    g593(.A(new_n672), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  XOR2_X1   g595(.A(KEYINPUT105), .B(G134), .Z(new_n782));
  XNOR2_X1  g596(.A(new_n781), .B(new_n782), .ZN(G36));
  INV_X1    g597(.A(new_n636), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n710), .A2(new_n628), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(KEYINPUT43), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n784), .B(new_n657), .C1(new_n786), .C2(KEYINPUT106), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n787), .B1(KEYINPUT106), .B2(new_n786), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n788), .A2(KEYINPUT44), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(KEYINPUT44), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT46), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n610), .A2(new_n612), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(KEYINPUT45), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n768), .A2(KEYINPUT45), .A3(new_n604), .A4(new_n770), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(G469), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n791), .B1(new_n797), .B2(new_n617), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n796), .A2(KEYINPUT46), .A3(new_n618), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n616), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n574), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n802), .A2(new_n675), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n767), .B(KEYINPUT107), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n789), .A2(new_n790), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G137), .ZN(G39));
  AND2_X1   g620(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n807));
  NOR2_X1   g621(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n802), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n801), .A2(new_n807), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n767), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n668), .A2(new_n244), .A3(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n812), .A2(new_n707), .A3(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G140), .ZN(G42));
  AND2_X1   g630(.A1(new_n786), .A2(new_n494), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n813), .A2(new_n715), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n817), .A2(new_n381), .A3(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(KEYINPUT48), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n700), .A2(new_n244), .A3(new_n494), .A4(new_n818), .ZN(new_n821));
  INV_X1    g635(.A(new_n629), .ZN(new_n822));
  OAI211_X1 g636(.A(G952), .B(new_n218), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n743), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n817), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n823), .B1(new_n825), .B2(new_n732), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n820), .A2(new_n826), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n827), .A2(KEYINPUT118), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(KEYINPUT118), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n817), .A2(new_n818), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n830), .A2(new_n757), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n821), .A2(new_n710), .A3(new_n711), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n703), .A2(new_n505), .A3(new_n716), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n825), .A2(KEYINPUT50), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT50), .B1(new_n825), .B2(new_n834), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n833), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n744), .A2(KEYINPUT115), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n744), .A2(KEYINPUT115), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n838), .A2(new_n573), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n840), .B1(new_n810), .B2(new_n811), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n825), .A2(new_n804), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n837), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n828), .B(new_n829), .C1(new_n843), .C2(KEYINPUT51), .ZN(new_n844));
  OR2_X1    g658(.A1(new_n841), .A2(KEYINPUT116), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n841), .A2(KEYINPUT116), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n845), .A2(new_n842), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n837), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n847), .A2(KEYINPUT51), .A3(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT117), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n847), .A2(new_n848), .A3(KEYINPUT117), .A4(KEYINPUT51), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n844), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n854));
  OAI22_X1  g668(.A1(new_n712), .A2(new_n719), .B1(new_n730), .B2(new_n733), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n855), .B1(new_n727), .B2(new_n725), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n781), .B1(new_n774), .B2(new_n777), .ZN(new_n857));
  AND4_X1   g671(.A1(new_n761), .A2(new_n773), .A3(new_n657), .A4(new_n741), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n574), .B1(new_n613), .B2(new_n619), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n492), .A2(new_n657), .A3(new_n670), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n444), .A2(new_n647), .ZN(new_n861));
  NOR4_X1   g675(.A1(new_n859), .A2(new_n813), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  AOI22_X1  g676(.A1(new_n858), .A2(new_n707), .B1(new_n862), .B2(new_n668), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n856), .A2(new_n754), .A3(new_n857), .A4(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT109), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n865), .B1(new_n622), .B2(new_n641), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n681), .A2(new_n682), .A3(new_n492), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n867), .A2(new_n631), .A3(new_n640), .A4(new_n636), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n658), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n622), .A2(new_n865), .A3(new_n641), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT53), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n864), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT52), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n759), .B1(new_n758), .B2(new_n707), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n762), .A2(new_n763), .A3(KEYINPUT103), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n673), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n237), .B1(new_n233), .B2(new_n234), .ZN(new_n880));
  AOI211_X1 g694(.A(KEYINPUT25), .B(G902), .C1(new_n232), .C2(new_n227), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n656), .B(new_n670), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(KEYINPUT111), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT111), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n238), .A2(new_n884), .A3(new_n656), .A4(new_n670), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(new_n574), .A3(new_n772), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n887), .B1(new_n369), .B2(new_n699), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n747), .A2(new_n888), .A3(new_n571), .A4(new_n749), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n708), .A2(new_n889), .ZN(new_n890));
  OAI211_X1 g704(.A(KEYINPUT112), .B(new_n876), .C1(new_n879), .C2(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n876), .B1(new_n879), .B2(new_n890), .ZN(new_n892));
  INV_X1    g706(.A(new_n673), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n893), .B1(new_n760), .B2(new_n764), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n708), .A2(new_n889), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n894), .A2(new_n895), .A3(KEYINPUT52), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT112), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n892), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n875), .A2(new_n891), .A3(new_n898), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n892), .A2(new_n896), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT110), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n901), .B1(new_n864), .B2(new_n873), .ZN(new_n902));
  AOI221_X4 g716(.A(new_n855), .B1(new_n727), .B2(new_n725), .C1(new_n751), .C2(new_n753), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n871), .A2(new_n866), .A3(new_n869), .ZN(new_n904));
  INV_X1    g718(.A(new_n781), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n778), .A2(new_n905), .A3(new_n863), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n903), .A2(KEYINPUT110), .A3(new_n904), .A4(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n900), .B1(new_n902), .B2(new_n907), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n854), .B(new_n899), .C1(new_n908), .C2(KEYINPUT53), .ZN(new_n909));
  OR2_X1    g723(.A1(new_n909), .A2(KEYINPUT113), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT114), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n909), .A2(KEYINPUT113), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n902), .A2(new_n907), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n874), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n898), .A2(new_n891), .ZN(new_n915));
  OAI221_X1 g729(.A(KEYINPUT54), .B1(new_n908), .B2(new_n874), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n910), .A2(new_n911), .A3(new_n912), .A4(new_n916), .ZN(new_n917));
  OAI22_X1  g731(.A1(new_n914), .A2(new_n915), .B1(new_n908), .B2(new_n874), .ZN(new_n918));
  OAI22_X1  g732(.A1(new_n918), .A2(new_n854), .B1(new_n909), .B2(KEYINPUT113), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n909), .A2(KEYINPUT113), .ZN(new_n920));
  OAI21_X1  g734(.A(KEYINPUT114), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n853), .A2(new_n917), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n922), .B1(G952), .B2(G953), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n714), .A2(new_n616), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n924), .A2(KEYINPUT49), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n924), .A2(KEYINPUT49), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n244), .A2(new_n504), .A3(new_n574), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n785), .A2(new_n700), .A3(new_n928), .A4(new_n703), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n923), .A2(new_n929), .ZN(G75));
  NOR2_X1   g744(.A1(new_n218), .A2(G952), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n560), .A2(new_n564), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(new_n562), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT55), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n899), .B1(new_n908), .B2(KEYINPUT53), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n935), .A2(G902), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(G210), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT56), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n934), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n936), .B(KEYINPUT119), .Z(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n568), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n934), .A2(new_n938), .ZN(new_n942));
  AOI211_X1 g756(.A(new_n931), .B(new_n939), .C1(new_n941), .C2(new_n942), .ZN(G51));
  INV_X1    g757(.A(KEYINPUT121), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n935), .A2(KEYINPUT54), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n909), .ZN(new_n946));
  XNOR2_X1  g760(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(new_n617), .ZN(new_n948));
  INV_X1    g762(.A(new_n592), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n591), .B1(new_n583), .B2(new_n590), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n603), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n592), .A2(new_n607), .A3(new_n597), .A4(new_n599), .ZN(new_n952));
  AOI22_X1  g766(.A1(new_n946), .A2(new_n948), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AOI22_X1  g767(.A1(new_n940), .A2(new_n797), .B1(new_n944), .B2(new_n953), .ZN(new_n954));
  OR2_X1    g768(.A1(new_n953), .A2(new_n944), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n931), .B1(new_n954), .B2(new_n955), .ZN(G54));
  AND2_X1   g770(.A1(KEYINPUT58), .A2(G475), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n940), .A2(new_n441), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n441), .B1(new_n940), .B2(new_n957), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n958), .A2(new_n959), .A3(new_n931), .ZN(G60));
  INV_X1    g774(.A(new_n626), .ZN(new_n961));
  NAND2_X1  g775(.A1(G478), .A2(G902), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT59), .Z(new_n963));
  NOR2_X1   g777(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n931), .B1(new_n946), .B2(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n963), .B1(new_n921), .B2(new_n917), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n965), .B1(new_n966), .B2(new_n626), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(KEYINPUT122), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT122), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n969), .B(new_n965), .C1(new_n966), .C2(new_n626), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n968), .A2(new_n970), .ZN(G63));
  NAND2_X1  g785(.A1(G217), .A2(G902), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT124), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT60), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n935), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n931), .B1(new_n975), .B2(new_n655), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n976), .B1(new_n240), .B2(new_n975), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(KEYINPUT123), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT61), .ZN(G66));
  AOI21_X1  g793(.A(new_n218), .B1(new_n498), .B2(G224), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n903), .A2(new_n904), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n980), .B1(new_n981), .B2(new_n218), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n932), .B1(G898), .B2(new_n218), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT125), .Z(new_n984));
  XNOR2_X1  g798(.A(new_n982), .B(new_n984), .ZN(G69));
  NOR2_X1   g799(.A1(new_n415), .A2(new_n416), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n322), .B(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n987), .B1(G900), .B2(G953), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n894), .A2(new_n708), .ZN(new_n989));
  AND3_X1   g803(.A1(new_n747), .A2(new_n571), .A3(new_n749), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n803), .A2(new_n381), .A3(new_n990), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n991), .A2(new_n857), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n805), .A2(new_n815), .A3(new_n989), .A4(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n988), .B1(new_n993), .B2(G953), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(KEYINPUT126), .ZN(new_n995));
  INV_X1    g809(.A(new_n987), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n989), .A2(new_n705), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT62), .Z(new_n998));
  NOR2_X1   g812(.A1(new_n676), .A2(new_n813), .ZN(new_n999));
  OAI211_X1 g813(.A(new_n381), .B(new_n999), .C1(new_n629), .C2(new_n867), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n805), .A2(new_n815), .A3(new_n998), .A4(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n996), .B1(new_n1001), .B2(new_n218), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n995), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n218), .B1(G227), .B2(G900), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1003), .B(new_n1004), .Z(G72));
  XNOR2_X1  g819(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1006), .B(new_n686), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1007), .B1(new_n1001), .B2(new_n981), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n347), .A2(new_n342), .ZN(new_n1009));
  AND2_X1   g823(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1007), .B1(new_n993), .B2(new_n981), .ZN(new_n1011));
  AND2_X1   g825(.A1(new_n1011), .A2(new_n373), .ZN(new_n1012));
  INV_X1    g826(.A(new_n373), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1013), .A2(new_n1007), .ZN(new_n1014));
  NOR3_X1   g828(.A1(new_n918), .A2(new_n1009), .A3(new_n1014), .ZN(new_n1015));
  NOR4_X1   g829(.A1(new_n1010), .A2(new_n1012), .A3(new_n931), .A4(new_n1015), .ZN(G57));
endmodule


