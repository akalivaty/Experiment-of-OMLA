

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U548 ( .A1(G1966), .A2(n791), .ZN(n732) );
  OR2_X1 U549 ( .A1(n791), .A2(n790), .ZN(n513) );
  AND2_X1 U550 ( .A1(n925), .A2(n756), .ZN(n514) );
  OR2_X1 U551 ( .A1(n754), .A2(KEYINPUT33), .ZN(n515) );
  AND2_X1 U552 ( .A1(n792), .A2(n513), .ZN(n516) );
  XOR2_X1 U553 ( .A(KEYINPUT29), .B(n714), .Z(n517) );
  XNOR2_X1 U554 ( .A(n692), .B(KEYINPUT26), .ZN(n693) );
  INV_X1 U555 ( .A(KEYINPUT31), .ZN(n727) );
  BUF_X1 U556 ( .A(n691), .Z(n737) );
  AND2_X1 U557 ( .A1(n744), .A2(n743), .ZN(n745) );
  INV_X1 U558 ( .A(KEYINPUT12), .ZN(n567) );
  XNOR2_X1 U559 ( .A(n567), .B(KEYINPUT71), .ZN(n568) );
  XNOR2_X1 U560 ( .A(n569), .B(n568), .ZN(n571) );
  NOR2_X1 U561 ( .A1(G651), .A2(G543), .ZN(n530) );
  AND2_X1 U562 ( .A1(n522), .A2(G2104), .ZN(n871) );
  NOR2_X1 U563 ( .A1(G651), .A2(n650), .ZN(n642) );
  NOR2_X1 U564 ( .A1(n574), .A2(n573), .ZN(n576) );
  NAND2_X1 U565 ( .A1(n576), .A2(n575), .ZN(n912) );
  AND2_X1 U566 ( .A1(G2105), .A2(G2104), .ZN(n875) );
  NAND2_X1 U567 ( .A1(G113), .A2(n875), .ZN(n518) );
  XNOR2_X1 U568 ( .A(n518), .B(KEYINPUT66), .ZN(n521) );
  INV_X1 U569 ( .A(G2105), .ZN(n522) );
  NAND2_X1 U570 ( .A1(G101), .A2(n871), .ZN(n519) );
  XOR2_X1 U571 ( .A(KEYINPUT23), .B(n519), .Z(n520) );
  NAND2_X1 U572 ( .A1(n521), .A2(n520), .ZN(n527) );
  NOR2_X1 U573 ( .A1(G2104), .A2(n522), .ZN(n877) );
  NAND2_X1 U574 ( .A1(G125), .A2(n877), .ZN(n525) );
  NOR2_X1 U575 ( .A1(G2104), .A2(G2105), .ZN(n523) );
  XOR2_X2 U576 ( .A(KEYINPUT17), .B(n523), .Z(n872) );
  NAND2_X1 U577 ( .A1(G137), .A2(n872), .ZN(n524) );
  NAND2_X1 U578 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X1 U579 ( .A1(n527), .A2(n526), .ZN(G160) );
  INV_X1 U580 ( .A(G651), .ZN(n533) );
  NOR2_X1 U581 ( .A1(G543), .A2(n533), .ZN(n529) );
  XNOR2_X1 U582 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n528) );
  XNOR2_X1 U583 ( .A(n529), .B(n528), .ZN(n648) );
  NAND2_X1 U584 ( .A1(G60), .A2(n648), .ZN(n532) );
  XOR2_X1 U585 ( .A(KEYINPUT65), .B(n530), .Z(n634) );
  NAND2_X1 U586 ( .A1(G85), .A2(n634), .ZN(n531) );
  NAND2_X1 U587 ( .A1(n532), .A2(n531), .ZN(n537) );
  XOR2_X1 U588 ( .A(KEYINPUT0), .B(G543), .Z(n650) );
  NAND2_X1 U589 ( .A1(G47), .A2(n642), .ZN(n535) );
  NOR2_X1 U590 ( .A1(n650), .A2(n533), .ZN(n631) );
  NAND2_X1 U591 ( .A1(G72), .A2(n631), .ZN(n534) );
  NAND2_X1 U592 ( .A1(n535), .A2(n534), .ZN(n536) );
  OR2_X1 U593 ( .A1(n537), .A2(n536), .ZN(G290) );
  AND2_X1 U594 ( .A1(G452), .A2(G94), .ZN(G173) );
  AND2_X1 U595 ( .A1(G138), .A2(n872), .ZN(n543) );
  NAND2_X1 U596 ( .A1(G114), .A2(n875), .ZN(n539) );
  NAND2_X1 U597 ( .A1(G126), .A2(n877), .ZN(n538) );
  AND2_X1 U598 ( .A1(n539), .A2(n538), .ZN(n541) );
  NAND2_X1 U599 ( .A1(G102), .A2(n871), .ZN(n540) );
  NAND2_X1 U600 ( .A1(n541), .A2(n540), .ZN(n542) );
  NOR2_X1 U601 ( .A1(n543), .A2(n542), .ZN(G164) );
  INV_X1 U602 ( .A(G57), .ZN(G237) );
  INV_X1 U603 ( .A(G132), .ZN(G219) );
  INV_X1 U604 ( .A(G82), .ZN(G220) );
  NAND2_X1 U605 ( .A1(n642), .A2(G52), .ZN(n545) );
  NAND2_X1 U606 ( .A1(n648), .A2(G64), .ZN(n544) );
  NAND2_X1 U607 ( .A1(n545), .A2(n544), .ZN(n551) );
  NAND2_X1 U608 ( .A1(G90), .A2(n634), .ZN(n547) );
  NAND2_X1 U609 ( .A1(G77), .A2(n631), .ZN(n546) );
  NAND2_X1 U610 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U611 ( .A(KEYINPUT9), .B(n548), .Z(n549) );
  XNOR2_X1 U612 ( .A(KEYINPUT68), .B(n549), .ZN(n550) );
  NOR2_X1 U613 ( .A1(n551), .A2(n550), .ZN(G171) );
  NAND2_X1 U614 ( .A1(n648), .A2(G63), .ZN(n552) );
  XNOR2_X1 U615 ( .A(KEYINPUT75), .B(n552), .ZN(n555) );
  NAND2_X1 U616 ( .A1(n642), .A2(G51), .ZN(n553) );
  XOR2_X1 U617 ( .A(KEYINPUT76), .B(n553), .Z(n554) );
  NOR2_X1 U618 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U619 ( .A(n556), .B(KEYINPUT6), .ZN(n562) );
  NAND2_X1 U620 ( .A1(n634), .A2(G89), .ZN(n557) );
  XNOR2_X1 U621 ( .A(n557), .B(KEYINPUT4), .ZN(n559) );
  NAND2_X1 U622 ( .A1(G76), .A2(n631), .ZN(n558) );
  NAND2_X1 U623 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U624 ( .A(KEYINPUT5), .B(n560), .ZN(n561) );
  NAND2_X1 U625 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U626 ( .A(n563), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U627 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U628 ( .A1(G7), .A2(G661), .ZN(n564) );
  XNOR2_X1 U629 ( .A(n564), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U630 ( .A(G223), .B(KEYINPUT70), .Z(n820) );
  NAND2_X1 U631 ( .A1(n820), .A2(G567), .ZN(n565) );
  XOR2_X1 U632 ( .A(KEYINPUT11), .B(n565), .Z(G234) );
  NAND2_X1 U633 ( .A1(G56), .A2(n648), .ZN(n566) );
  XOR2_X1 U634 ( .A(KEYINPUT14), .B(n566), .Z(n574) );
  NAND2_X1 U635 ( .A1(G81), .A2(n634), .ZN(n569) );
  NAND2_X1 U636 ( .A1(G68), .A2(n631), .ZN(n570) );
  AND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(KEYINPUT13), .B(n572), .ZN(n573) );
  NAND2_X1 U639 ( .A1(n642), .A2(G43), .ZN(n575) );
  INV_X1 U640 ( .A(G860), .ZN(n614) );
  OR2_X1 U641 ( .A1(n912), .A2(n614), .ZN(G153) );
  INV_X1 U642 ( .A(G171), .ZN(G301) );
  NAND2_X1 U643 ( .A1(G66), .A2(n648), .ZN(n578) );
  NAND2_X1 U644 ( .A1(G92), .A2(n634), .ZN(n577) );
  NAND2_X1 U645 ( .A1(n578), .A2(n577), .ZN(n582) );
  NAND2_X1 U646 ( .A1(G54), .A2(n642), .ZN(n580) );
  NAND2_X1 U647 ( .A1(G79), .A2(n631), .ZN(n579) );
  NAND2_X1 U648 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U649 ( .A1(n582), .A2(n581), .ZN(n584) );
  XNOR2_X1 U650 ( .A(KEYINPUT72), .B(KEYINPUT15), .ZN(n583) );
  XOR2_X1 U651 ( .A(n584), .B(n583), .Z(n917) );
  NOR2_X1 U652 ( .A1(G868), .A2(n917), .ZN(n585) );
  XNOR2_X1 U653 ( .A(n585), .B(KEYINPUT73), .ZN(n587) );
  NAND2_X1 U654 ( .A1(G868), .A2(G301), .ZN(n586) );
  NAND2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U656 ( .A(KEYINPUT74), .B(n588), .ZN(G284) );
  NAND2_X1 U657 ( .A1(G65), .A2(n648), .ZN(n590) );
  NAND2_X1 U658 ( .A1(G78), .A2(n631), .ZN(n589) );
  NAND2_X1 U659 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U660 ( .A1(G91), .A2(n634), .ZN(n591) );
  XNOR2_X1 U661 ( .A(KEYINPUT69), .B(n591), .ZN(n592) );
  NOR2_X1 U662 ( .A1(n593), .A2(n592), .ZN(n595) );
  NAND2_X1 U663 ( .A1(n642), .A2(G53), .ZN(n594) );
  NAND2_X1 U664 ( .A1(n595), .A2(n594), .ZN(G299) );
  INV_X1 U665 ( .A(G868), .ZN(n663) );
  NOR2_X1 U666 ( .A1(G286), .A2(n663), .ZN(n597) );
  NOR2_X1 U667 ( .A1(G868), .A2(G299), .ZN(n596) );
  NOR2_X1 U668 ( .A1(n597), .A2(n596), .ZN(G297) );
  NAND2_X1 U669 ( .A1(n614), .A2(G559), .ZN(n598) );
  NAND2_X1 U670 ( .A1(n598), .A2(n917), .ZN(n599) );
  XNOR2_X1 U671 ( .A(n599), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U672 ( .A1(G868), .A2(n912), .ZN(n602) );
  NAND2_X1 U673 ( .A1(n917), .A2(G868), .ZN(n600) );
  NOR2_X1 U674 ( .A1(G559), .A2(n600), .ZN(n601) );
  NOR2_X1 U675 ( .A1(n602), .A2(n601), .ZN(G282) );
  XOR2_X1 U676 ( .A(G2100), .B(KEYINPUT78), .Z(n612) );
  NAND2_X1 U677 ( .A1(G123), .A2(n877), .ZN(n603) );
  XNOR2_X1 U678 ( .A(n603), .B(KEYINPUT18), .ZN(n606) );
  NAND2_X1 U679 ( .A1(G111), .A2(n875), .ZN(n604) );
  XOR2_X1 U680 ( .A(KEYINPUT77), .B(n604), .Z(n605) );
  NAND2_X1 U681 ( .A1(n606), .A2(n605), .ZN(n610) );
  NAND2_X1 U682 ( .A1(G99), .A2(n871), .ZN(n608) );
  NAND2_X1 U683 ( .A1(G135), .A2(n872), .ZN(n607) );
  NAND2_X1 U684 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U685 ( .A1(n610), .A2(n609), .ZN(n993) );
  XNOR2_X1 U686 ( .A(n993), .B(G2096), .ZN(n611) );
  NAND2_X1 U687 ( .A1(n612), .A2(n611), .ZN(G156) );
  NAND2_X1 U688 ( .A1(n917), .A2(G559), .ZN(n613) );
  XOR2_X1 U689 ( .A(n912), .B(n613), .Z(n660) );
  NAND2_X1 U690 ( .A1(n614), .A2(n660), .ZN(n622) );
  NAND2_X1 U691 ( .A1(G67), .A2(n648), .ZN(n616) );
  NAND2_X1 U692 ( .A1(G93), .A2(n634), .ZN(n615) );
  NAND2_X1 U693 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U694 ( .A1(G80), .A2(n631), .ZN(n617) );
  XNOR2_X1 U695 ( .A(KEYINPUT79), .B(n617), .ZN(n618) );
  NOR2_X1 U696 ( .A1(n619), .A2(n618), .ZN(n621) );
  NAND2_X1 U697 ( .A1(n642), .A2(G55), .ZN(n620) );
  NAND2_X1 U698 ( .A1(n621), .A2(n620), .ZN(n664) );
  XNOR2_X1 U699 ( .A(n622), .B(n664), .ZN(G145) );
  NAND2_X1 U700 ( .A1(G88), .A2(n634), .ZN(n629) );
  NAND2_X1 U701 ( .A1(G62), .A2(n648), .ZN(n624) );
  NAND2_X1 U702 ( .A1(G50), .A2(n642), .ZN(n623) );
  NAND2_X1 U703 ( .A1(n624), .A2(n623), .ZN(n627) );
  NAND2_X1 U704 ( .A1(G75), .A2(n631), .ZN(n625) );
  XNOR2_X1 U705 ( .A(KEYINPUT85), .B(n625), .ZN(n626) );
  NOR2_X1 U706 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U707 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U708 ( .A(n630), .B(KEYINPUT86), .Z(G166) );
  XOR2_X1 U709 ( .A(KEYINPUT84), .B(KEYINPUT2), .Z(n633) );
  NAND2_X1 U710 ( .A1(G73), .A2(n631), .ZN(n632) );
  XNOR2_X1 U711 ( .A(n633), .B(n632), .ZN(n639) );
  NAND2_X1 U712 ( .A1(G61), .A2(n648), .ZN(n636) );
  NAND2_X1 U713 ( .A1(G86), .A2(n634), .ZN(n635) );
  NAND2_X1 U714 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U715 ( .A(KEYINPUT83), .B(n637), .Z(n638) );
  NOR2_X1 U716 ( .A1(n639), .A2(n638), .ZN(n641) );
  NAND2_X1 U717 ( .A1(n642), .A2(G48), .ZN(n640) );
  NAND2_X1 U718 ( .A1(n641), .A2(n640), .ZN(G305) );
  NAND2_X1 U719 ( .A1(n642), .A2(G49), .ZN(n643) );
  XNOR2_X1 U720 ( .A(n643), .B(KEYINPUT80), .ZN(n645) );
  NAND2_X1 U721 ( .A1(G74), .A2(G651), .ZN(n644) );
  NAND2_X1 U722 ( .A1(n645), .A2(n644), .ZN(n646) );
  XOR2_X1 U723 ( .A(KEYINPUT81), .B(n646), .Z(n647) );
  NOR2_X1 U724 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U725 ( .A(n649), .B(KEYINPUT82), .ZN(n652) );
  NAND2_X1 U726 ( .A1(G87), .A2(n650), .ZN(n651) );
  NAND2_X1 U727 ( .A1(n652), .A2(n651), .ZN(G288) );
  XOR2_X1 U728 ( .A(G299), .B(n664), .Z(n657) );
  XNOR2_X1 U729 ( .A(KEYINPUT87), .B(KEYINPUT88), .ZN(n654) );
  XNOR2_X1 U730 ( .A(G290), .B(KEYINPUT19), .ZN(n653) );
  XNOR2_X1 U731 ( .A(n654), .B(n653), .ZN(n655) );
  XOR2_X1 U732 ( .A(G166), .B(n655), .Z(n656) );
  XNOR2_X1 U733 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U734 ( .A(n658), .B(G305), .ZN(n659) );
  XNOR2_X1 U735 ( .A(n659), .B(G288), .ZN(n888) );
  XNOR2_X1 U736 ( .A(n888), .B(n660), .ZN(n661) );
  NAND2_X1 U737 ( .A1(n661), .A2(G868), .ZN(n662) );
  XOR2_X1 U738 ( .A(KEYINPUT89), .B(n662), .Z(n666) );
  NAND2_X1 U739 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U740 ( .A1(n666), .A2(n665), .ZN(G295) );
  XNOR2_X1 U741 ( .A(KEYINPUT20), .B(KEYINPUT91), .ZN(n669) );
  NAND2_X1 U742 ( .A1(G2078), .A2(G2084), .ZN(n667) );
  XNOR2_X1 U743 ( .A(n667), .B(KEYINPUT90), .ZN(n668) );
  XNOR2_X1 U744 ( .A(n669), .B(n668), .ZN(n670) );
  NAND2_X1 U745 ( .A1(G2090), .A2(n670), .ZN(n671) );
  XNOR2_X1 U746 ( .A(KEYINPUT21), .B(n671), .ZN(n672) );
  NAND2_X1 U747 ( .A1(n672), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U748 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U749 ( .A1(G220), .A2(G219), .ZN(n673) );
  XNOR2_X1 U750 ( .A(KEYINPUT22), .B(n673), .ZN(n674) );
  NAND2_X1 U751 ( .A1(n674), .A2(G96), .ZN(n675) );
  NOR2_X1 U752 ( .A1(G218), .A2(n675), .ZN(n676) );
  XOR2_X1 U753 ( .A(KEYINPUT92), .B(n676), .Z(n910) );
  NAND2_X1 U754 ( .A1(n910), .A2(G2106), .ZN(n680) );
  NAND2_X1 U755 ( .A1(G120), .A2(G108), .ZN(n677) );
  NOR2_X1 U756 ( .A1(G237), .A2(n677), .ZN(n678) );
  NAND2_X1 U757 ( .A1(G69), .A2(n678), .ZN(n909) );
  NAND2_X1 U758 ( .A1(G567), .A2(n909), .ZN(n679) );
  NAND2_X1 U759 ( .A1(n680), .A2(n679), .ZN(n825) );
  NAND2_X1 U760 ( .A1(G483), .A2(G661), .ZN(n681) );
  NOR2_X1 U761 ( .A1(n825), .A2(n681), .ZN(n822) );
  NAND2_X1 U762 ( .A1(n822), .A2(G36), .ZN(G176) );
  INV_X1 U763 ( .A(G166), .ZN(G303) );
  NAND2_X1 U764 ( .A1(G160), .A2(G40), .ZN(n784) );
  NOR2_X2 U765 ( .A1(G164), .A2(G1384), .ZN(n785) );
  INV_X1 U766 ( .A(n785), .ZN(n684) );
  NOR2_X4 U767 ( .A1(n784), .A2(n684), .ZN(n715) );
  INV_X1 U768 ( .A(n715), .ZN(n691) );
  NAND2_X1 U769 ( .A1(n691), .A2(G8), .ZN(n685) );
  XNOR2_X1 U770 ( .A(KEYINPUT97), .B(n685), .ZN(n686) );
  NAND2_X1 U771 ( .A1(G1976), .A2(G288), .ZN(n928) );
  NAND2_X1 U772 ( .A1(n686), .A2(n928), .ZN(n752) );
  NOR2_X1 U773 ( .A1(G303), .A2(G1971), .ZN(n750) );
  NOR2_X1 U774 ( .A1(G2084), .A2(n737), .ZN(n721) );
  NAND2_X1 U775 ( .A1(G8), .A2(n721), .ZN(n734) );
  INV_X1 U776 ( .A(n686), .ZN(n791) );
  NAND2_X1 U777 ( .A1(G1348), .A2(n691), .ZN(n688) );
  NAND2_X1 U778 ( .A1(n715), .A2(G2067), .ZN(n687) );
  NAND2_X1 U779 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U780 ( .A(n689), .B(KEYINPUT100), .Z(n690) );
  NAND2_X1 U781 ( .A1(n917), .A2(n690), .ZN(n700) );
  OR2_X1 U782 ( .A1(n917), .A2(n690), .ZN(n698) );
  INV_X1 U783 ( .A(G1996), .ZN(n940) );
  NOR2_X1 U784 ( .A1(n691), .A2(n940), .ZN(n692) );
  INV_X1 U785 ( .A(n693), .ZN(n695) );
  NAND2_X1 U786 ( .A1(n737), .A2(G1341), .ZN(n694) );
  NAND2_X1 U787 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U788 ( .A1(n912), .A2(n696), .ZN(n697) );
  NAND2_X1 U789 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U790 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U791 ( .A(n701), .B(KEYINPUT101), .ZN(n707) );
  INV_X1 U792 ( .A(G299), .ZN(n709) );
  NAND2_X1 U793 ( .A1(G1956), .A2(n737), .ZN(n704) );
  NAND2_X1 U794 ( .A1(n715), .A2(G2072), .ZN(n702) );
  XOR2_X1 U795 ( .A(KEYINPUT27), .B(n702), .Z(n703) );
  NAND2_X1 U796 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U797 ( .A(KEYINPUT98), .B(n705), .Z(n708) );
  NAND2_X1 U798 ( .A1(n709), .A2(n708), .ZN(n706) );
  NAND2_X1 U799 ( .A1(n707), .A2(n706), .ZN(n713) );
  NOR2_X1 U800 ( .A1(n709), .A2(n708), .ZN(n711) );
  XNOR2_X1 U801 ( .A(KEYINPUT99), .B(KEYINPUT28), .ZN(n710) );
  XNOR2_X1 U802 ( .A(n711), .B(n710), .ZN(n712) );
  NAND2_X1 U803 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U804 ( .A1(G1961), .A2(n737), .ZN(n717) );
  XOR2_X1 U805 ( .A(KEYINPUT25), .B(G2078), .Z(n939) );
  NAND2_X1 U806 ( .A1(n715), .A2(n939), .ZN(n716) );
  NAND2_X1 U807 ( .A1(n717), .A2(n716), .ZN(n719) );
  OR2_X1 U808 ( .A1(G301), .A2(n719), .ZN(n718) );
  NAND2_X1 U809 ( .A1(n517), .A2(n718), .ZN(n730) );
  NAND2_X1 U810 ( .A1(G301), .A2(n719), .ZN(n720) );
  XOR2_X1 U811 ( .A(KEYINPUT102), .B(n720), .Z(n726) );
  NOR2_X1 U812 ( .A1(n732), .A2(n721), .ZN(n722) );
  NAND2_X1 U813 ( .A1(G8), .A2(n722), .ZN(n723) );
  XNOR2_X1 U814 ( .A(KEYINPUT30), .B(n723), .ZN(n724) );
  NOR2_X1 U815 ( .A1(G168), .A2(n724), .ZN(n725) );
  NOR2_X1 U816 ( .A1(n726), .A2(n725), .ZN(n728) );
  XNOR2_X1 U817 ( .A(n728), .B(n727), .ZN(n729) );
  NAND2_X1 U818 ( .A1(n730), .A2(n729), .ZN(n736) );
  INV_X1 U819 ( .A(n736), .ZN(n731) );
  NOR2_X1 U820 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U821 ( .A1(n734), .A2(n733), .ZN(n747) );
  AND2_X1 U822 ( .A1(G286), .A2(G8), .ZN(n735) );
  NAND2_X1 U823 ( .A1(n736), .A2(n735), .ZN(n744) );
  INV_X1 U824 ( .A(G8), .ZN(n742) );
  NOR2_X1 U825 ( .A1(G1971), .A2(n791), .ZN(n739) );
  NOR2_X1 U826 ( .A1(G2090), .A2(n737), .ZN(n738) );
  NOR2_X1 U827 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U828 ( .A1(n740), .A2(G303), .ZN(n741) );
  OR2_X1 U829 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U830 ( .A(n745), .B(KEYINPUT32), .ZN(n746) );
  NAND2_X1 U831 ( .A1(n747), .A2(n746), .ZN(n759) );
  NOR2_X1 U832 ( .A1(G288), .A2(G1976), .ZN(n748) );
  XNOR2_X1 U833 ( .A(n748), .B(KEYINPUT103), .ZN(n932) );
  NAND2_X1 U834 ( .A1(n759), .A2(n932), .ZN(n749) );
  NOR2_X1 U835 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U836 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U837 ( .A(n753), .B(KEYINPUT64), .ZN(n754) );
  XOR2_X1 U838 ( .A(G1981), .B(G305), .Z(n925) );
  NOR2_X1 U839 ( .A1(n791), .A2(n932), .ZN(n755) );
  NAND2_X1 U840 ( .A1(KEYINPUT33), .A2(n755), .ZN(n756) );
  NAND2_X1 U841 ( .A1(n515), .A2(n514), .ZN(n793) );
  NOR2_X1 U842 ( .A1(G303), .A2(G2090), .ZN(n757) );
  XNOR2_X1 U843 ( .A(KEYINPUT104), .B(n757), .ZN(n758) );
  NAND2_X1 U844 ( .A1(n758), .A2(G8), .ZN(n760) );
  NAND2_X1 U845 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U846 ( .A1(n761), .A2(n791), .ZN(n788) );
  NAND2_X1 U847 ( .A1(G105), .A2(n871), .ZN(n762) );
  XNOR2_X1 U848 ( .A(n762), .B(KEYINPUT38), .ZN(n763) );
  XNOR2_X1 U849 ( .A(n763), .B(KEYINPUT96), .ZN(n765) );
  NAND2_X1 U850 ( .A1(G117), .A2(n875), .ZN(n764) );
  NAND2_X1 U851 ( .A1(n765), .A2(n764), .ZN(n769) );
  NAND2_X1 U852 ( .A1(G129), .A2(n877), .ZN(n767) );
  NAND2_X1 U853 ( .A1(G141), .A2(n872), .ZN(n766) );
  NAND2_X1 U854 ( .A1(n767), .A2(n766), .ZN(n768) );
  NOR2_X1 U855 ( .A1(n769), .A2(n768), .ZN(n864) );
  AND2_X1 U856 ( .A1(n940), .A2(n864), .ZN(n987) );
  NOR2_X1 U857 ( .A1(G1986), .A2(G290), .ZN(n776) );
  NAND2_X1 U858 ( .A1(G107), .A2(n875), .ZN(n771) );
  NAND2_X1 U859 ( .A1(G119), .A2(n877), .ZN(n770) );
  NAND2_X1 U860 ( .A1(n771), .A2(n770), .ZN(n775) );
  NAND2_X1 U861 ( .A1(G95), .A2(n871), .ZN(n773) );
  NAND2_X1 U862 ( .A1(G131), .A2(n872), .ZN(n772) );
  NAND2_X1 U863 ( .A1(n773), .A2(n772), .ZN(n774) );
  OR2_X1 U864 ( .A1(n775), .A2(n774), .ZN(n863) );
  NOR2_X1 U865 ( .A1(G1991), .A2(n863), .ZN(n994) );
  NOR2_X1 U866 ( .A1(n776), .A2(n994), .ZN(n780) );
  NAND2_X1 U867 ( .A1(G1991), .A2(n863), .ZN(n777) );
  XNOR2_X1 U868 ( .A(n777), .B(KEYINPUT95), .ZN(n779) );
  NOR2_X1 U869 ( .A1(n940), .A2(n864), .ZN(n778) );
  NOR2_X1 U870 ( .A1(n779), .A2(n778), .ZN(n795) );
  INV_X1 U871 ( .A(n795), .ZN(n1000) );
  NOR2_X1 U872 ( .A1(n780), .A2(n1000), .ZN(n781) );
  NOR2_X1 U873 ( .A1(n987), .A2(n781), .ZN(n782) );
  XOR2_X1 U874 ( .A(n782), .B(KEYINPUT105), .Z(n783) );
  XNOR2_X1 U875 ( .A(KEYINPUT39), .B(n783), .ZN(n787) );
  NOR2_X1 U876 ( .A1(n785), .A2(n784), .ZN(n786) );
  XOR2_X1 U877 ( .A(KEYINPUT93), .B(n786), .Z(n815) );
  NAND2_X1 U878 ( .A1(n787), .A2(n815), .ZN(n794) );
  AND2_X1 U879 ( .A1(n788), .A2(n794), .ZN(n792) );
  NOR2_X1 U880 ( .A1(G1981), .A2(G305), .ZN(n789) );
  XOR2_X1 U881 ( .A(n789), .B(KEYINPUT24), .Z(n790) );
  NAND2_X1 U882 ( .A1(n793), .A2(n516), .ZN(n800) );
  INV_X1 U883 ( .A(n794), .ZN(n798) );
  XOR2_X1 U884 ( .A(G1986), .B(G290), .Z(n915) );
  NAND2_X1 U885 ( .A1(n915), .A2(n795), .ZN(n796) );
  NAND2_X1 U886 ( .A1(n796), .A2(n815), .ZN(n797) );
  OR2_X1 U887 ( .A1(n798), .A2(n797), .ZN(n799) );
  AND2_X1 U888 ( .A1(n800), .A2(n799), .ZN(n812) );
  NAND2_X1 U889 ( .A1(G104), .A2(n871), .ZN(n802) );
  NAND2_X1 U890 ( .A1(G140), .A2(n872), .ZN(n801) );
  NAND2_X1 U891 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U892 ( .A(KEYINPUT34), .B(n803), .ZN(n809) );
  NAND2_X1 U893 ( .A1(G116), .A2(n875), .ZN(n805) );
  NAND2_X1 U894 ( .A1(G128), .A2(n877), .ZN(n804) );
  NAND2_X1 U895 ( .A1(n805), .A2(n804), .ZN(n806) );
  XOR2_X1 U896 ( .A(KEYINPUT94), .B(n806), .Z(n807) );
  XNOR2_X1 U897 ( .A(KEYINPUT35), .B(n807), .ZN(n808) );
  NOR2_X1 U898 ( .A1(n809), .A2(n808), .ZN(n810) );
  XOR2_X1 U899 ( .A(KEYINPUT36), .B(n810), .Z(n884) );
  XOR2_X1 U900 ( .A(G2067), .B(KEYINPUT37), .Z(n813) );
  AND2_X1 U901 ( .A1(n884), .A2(n813), .ZN(n996) );
  NAND2_X1 U902 ( .A1(n996), .A2(n815), .ZN(n811) );
  NAND2_X1 U903 ( .A1(n812), .A2(n811), .ZN(n817) );
  NOR2_X1 U904 ( .A1(n813), .A2(n884), .ZN(n814) );
  XNOR2_X1 U905 ( .A(n814), .B(KEYINPUT106), .ZN(n992) );
  NAND2_X1 U906 ( .A1(n992), .A2(n815), .ZN(n816) );
  NAND2_X1 U907 ( .A1(n817), .A2(n816), .ZN(n819) );
  XOR2_X1 U908 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n818) );
  XNOR2_X1 U909 ( .A(n819), .B(n818), .ZN(G329) );
  NAND2_X1 U910 ( .A1(G2106), .A2(n820), .ZN(G217) );
  AND2_X1 U911 ( .A1(G15), .A2(G2), .ZN(n821) );
  NAND2_X1 U912 ( .A1(G661), .A2(n821), .ZN(G259) );
  NAND2_X1 U913 ( .A1(G1), .A2(G3), .ZN(n823) );
  NAND2_X1 U914 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U915 ( .A(n824), .B(KEYINPUT110), .ZN(G188) );
  XNOR2_X1 U916 ( .A(KEYINPUT111), .B(n825), .ZN(G319) );
  XOR2_X1 U917 ( .A(G2100), .B(KEYINPUT43), .Z(n827) );
  XNOR2_X1 U918 ( .A(G2090), .B(G2678), .ZN(n826) );
  XNOR2_X1 U919 ( .A(n827), .B(n826), .ZN(n828) );
  XOR2_X1 U920 ( .A(n828), .B(KEYINPUT42), .Z(n830) );
  XNOR2_X1 U921 ( .A(G2072), .B(G2067), .ZN(n829) );
  XNOR2_X1 U922 ( .A(n830), .B(n829), .ZN(n834) );
  XOR2_X1 U923 ( .A(KEYINPUT112), .B(G2096), .Z(n832) );
  XNOR2_X1 U924 ( .A(G2078), .B(G2084), .ZN(n831) );
  XNOR2_X1 U925 ( .A(n832), .B(n831), .ZN(n833) );
  XNOR2_X1 U926 ( .A(n834), .B(n833), .ZN(G227) );
  XOR2_X1 U927 ( .A(G1986), .B(G1976), .Z(n836) );
  XNOR2_X1 U928 ( .A(G1966), .B(G1981), .ZN(n835) );
  XNOR2_X1 U929 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U930 ( .A(n837), .B(KEYINPUT41), .Z(n839) );
  XNOR2_X1 U931 ( .A(G1961), .B(G1971), .ZN(n838) );
  XNOR2_X1 U932 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U933 ( .A(G2474), .B(G1991), .Z(n841) );
  XOR2_X1 U934 ( .A(G1956), .B(n940), .Z(n840) );
  XNOR2_X1 U935 ( .A(n841), .B(n840), .ZN(n842) );
  XNOR2_X1 U936 ( .A(n843), .B(n842), .ZN(G229) );
  NAND2_X1 U937 ( .A1(G112), .A2(n875), .ZN(n845) );
  NAND2_X1 U938 ( .A1(G100), .A2(n871), .ZN(n844) );
  NAND2_X1 U939 ( .A1(n845), .A2(n844), .ZN(n851) );
  NAND2_X1 U940 ( .A1(n877), .A2(G124), .ZN(n846) );
  XNOR2_X1 U941 ( .A(n846), .B(KEYINPUT44), .ZN(n848) );
  NAND2_X1 U942 ( .A1(G136), .A2(n872), .ZN(n847) );
  NAND2_X1 U943 ( .A1(n848), .A2(n847), .ZN(n849) );
  XOR2_X1 U944 ( .A(KEYINPUT113), .B(n849), .Z(n850) );
  NOR2_X1 U945 ( .A1(n851), .A2(n850), .ZN(G162) );
  NAND2_X1 U946 ( .A1(G106), .A2(n871), .ZN(n853) );
  NAND2_X1 U947 ( .A1(G142), .A2(n872), .ZN(n852) );
  NAND2_X1 U948 ( .A1(n853), .A2(n852), .ZN(n854) );
  XNOR2_X1 U949 ( .A(n854), .B(KEYINPUT45), .ZN(n856) );
  NAND2_X1 U950 ( .A1(G118), .A2(n875), .ZN(n855) );
  NAND2_X1 U951 ( .A1(n856), .A2(n855), .ZN(n859) );
  NAND2_X1 U952 ( .A1(n877), .A2(G130), .ZN(n857) );
  XOR2_X1 U953 ( .A(KEYINPUT114), .B(n857), .Z(n858) );
  NOR2_X1 U954 ( .A1(n859), .A2(n858), .ZN(n868) );
  XOR2_X1 U955 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n861) );
  XNOR2_X1 U956 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n860) );
  XNOR2_X1 U957 ( .A(n861), .B(n860), .ZN(n862) );
  XNOR2_X1 U958 ( .A(n863), .B(n862), .ZN(n866) );
  XNOR2_X1 U959 ( .A(G164), .B(n864), .ZN(n865) );
  XNOR2_X1 U960 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U961 ( .A(n868), .B(n867), .Z(n870) );
  XNOR2_X1 U962 ( .A(G160), .B(n993), .ZN(n869) );
  XNOR2_X1 U963 ( .A(n870), .B(n869), .ZN(n883) );
  NAND2_X1 U964 ( .A1(G103), .A2(n871), .ZN(n874) );
  NAND2_X1 U965 ( .A1(G139), .A2(n872), .ZN(n873) );
  NAND2_X1 U966 ( .A1(n874), .A2(n873), .ZN(n882) );
  NAND2_X1 U967 ( .A1(n875), .A2(G115), .ZN(n876) );
  XOR2_X1 U968 ( .A(KEYINPUT115), .B(n876), .Z(n879) );
  NAND2_X1 U969 ( .A1(n877), .A2(G127), .ZN(n878) );
  NAND2_X1 U970 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U971 ( .A(KEYINPUT47), .B(n880), .Z(n881) );
  NOR2_X1 U972 ( .A1(n882), .A2(n881), .ZN(n981) );
  XOR2_X1 U973 ( .A(n883), .B(n981), .Z(n886) );
  XNOR2_X1 U974 ( .A(n884), .B(G162), .ZN(n885) );
  XNOR2_X1 U975 ( .A(n886), .B(n885), .ZN(n887) );
  NOR2_X1 U976 ( .A1(G37), .A2(n887), .ZN(G395) );
  XOR2_X1 U977 ( .A(n888), .B(G286), .Z(n890) );
  XOR2_X1 U978 ( .A(G171), .B(n917), .Z(n889) );
  XNOR2_X1 U979 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U980 ( .A(n891), .B(n912), .ZN(n892) );
  NOR2_X1 U981 ( .A1(G37), .A2(n892), .ZN(G397) );
  XNOR2_X1 U982 ( .A(KEYINPUT108), .B(G2454), .ZN(n901) );
  XNOR2_X1 U983 ( .A(G2430), .B(G2435), .ZN(n899) );
  XOR2_X1 U984 ( .A(G2451), .B(G2427), .Z(n894) );
  XNOR2_X1 U985 ( .A(G2438), .B(G2446), .ZN(n893) );
  XNOR2_X1 U986 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U987 ( .A(n895), .B(G2443), .Z(n897) );
  XNOR2_X1 U988 ( .A(G1341), .B(G1348), .ZN(n896) );
  XNOR2_X1 U989 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U990 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U991 ( .A(n901), .B(n900), .ZN(n902) );
  NAND2_X1 U992 ( .A1(n902), .A2(G14), .ZN(n903) );
  XOR2_X1 U993 ( .A(KEYINPUT109), .B(n903), .Z(n911) );
  NAND2_X1 U994 ( .A1(G319), .A2(n911), .ZN(n906) );
  NOR2_X1 U995 ( .A1(G227), .A2(G229), .ZN(n904) );
  XNOR2_X1 U996 ( .A(KEYINPUT49), .B(n904), .ZN(n905) );
  NOR2_X1 U997 ( .A1(n906), .A2(n905), .ZN(n908) );
  NOR2_X1 U998 ( .A1(G395), .A2(G397), .ZN(n907) );
  NAND2_X1 U999 ( .A1(n908), .A2(n907), .ZN(G225) );
  XOR2_X1 U1000 ( .A(KEYINPUT118), .B(G225), .Z(G308) );
  XNOR2_X1 U1001 ( .A(G108), .B(KEYINPUT119), .ZN(G238) );
  INV_X1 U1003 ( .A(G120), .ZN(G236) );
  INV_X1 U1004 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1005 ( .A1(n910), .A2(n909), .ZN(G325) );
  INV_X1 U1006 ( .A(G325), .ZN(G261) );
  INV_X1 U1007 ( .A(G69), .ZN(G235) );
  INV_X1 U1008 ( .A(n911), .ZN(G401) );
  XNOR2_X1 U1009 ( .A(KEYINPUT56), .B(G16), .ZN(n935) );
  XNOR2_X1 U1010 ( .A(n912), .B(G1341), .ZN(n914) );
  XOR2_X1 U1011 ( .A(G166), .B(G1971), .Z(n913) );
  NOR2_X1 U1012 ( .A1(n914), .A2(n913), .ZN(n924) );
  XOR2_X1 U1013 ( .A(G299), .B(G1956), .Z(n916) );
  NAND2_X1 U1014 ( .A1(n916), .A2(n915), .ZN(n922) );
  XOR2_X1 U1015 ( .A(G171), .B(G1961), .Z(n919) );
  XOR2_X1 U1016 ( .A(n917), .B(G1348), .Z(n918) );
  NOR2_X1 U1017 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1018 ( .A(KEYINPUT124), .B(n920), .Z(n921) );
  NOR2_X1 U1019 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(n931) );
  XNOR2_X1 U1021 ( .A(G1966), .B(G168), .ZN(n926) );
  NAND2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1023 ( .A(n927), .B(KEYINPUT57), .ZN(n929) );
  NAND2_X1 U1024 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1025 ( .A1(n931), .A2(n930), .ZN(n933) );
  NAND2_X1 U1026 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1027 ( .A1(n935), .A2(n934), .ZN(n1013) );
  XOR2_X1 U1028 ( .A(G1991), .B(G25), .Z(n936) );
  NAND2_X1 U1029 ( .A1(n936), .A2(G28), .ZN(n946) );
  XNOR2_X1 U1030 ( .A(G2072), .B(G33), .ZN(n938) );
  XNOR2_X1 U1031 ( .A(G2067), .B(G26), .ZN(n937) );
  NOR2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n944) );
  XNOR2_X1 U1033 ( .A(n939), .B(G27), .ZN(n942) );
  XOR2_X1 U1034 ( .A(n940), .B(G32), .Z(n941) );
  NOR2_X1 U1035 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1036 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1037 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1038 ( .A(KEYINPUT53), .B(n947), .Z(n951) );
  XNOR2_X1 U1039 ( .A(KEYINPUT54), .B(G34), .ZN(n948) );
  XNOR2_X1 U1040 ( .A(n948), .B(KEYINPUT123), .ZN(n949) );
  XNOR2_X1 U1041 ( .A(G2084), .B(n949), .ZN(n950) );
  NAND2_X1 U1042 ( .A1(n951), .A2(n950), .ZN(n953) );
  XNOR2_X1 U1043 ( .A(G35), .B(G2090), .ZN(n952) );
  OR2_X1 U1044 ( .A1(n953), .A2(n952), .ZN(n977) );
  XOR2_X1 U1045 ( .A(KEYINPUT55), .B(KEYINPUT122), .Z(n1005) );
  OR2_X1 U1046 ( .A1(n977), .A2(n1005), .ZN(n954) );
  NAND2_X1 U1047 ( .A1(G11), .A2(n954), .ZN(n1011) );
  XOR2_X1 U1048 ( .A(G1986), .B(G24), .Z(n958) );
  XNOR2_X1 U1049 ( .A(G1971), .B(G22), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(G23), .B(G1976), .ZN(n955) );
  NOR2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n960) );
  XNOR2_X1 U1053 ( .A(KEYINPUT125), .B(KEYINPUT58), .ZN(n959) );
  XNOR2_X1 U1054 ( .A(n960), .B(n959), .ZN(n964) );
  XNOR2_X1 U1055 ( .A(G1966), .B(G21), .ZN(n962) );
  XNOR2_X1 U1056 ( .A(G5), .B(G1961), .ZN(n961) );
  NOR2_X1 U1057 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n974) );
  XOR2_X1 U1059 ( .A(G1348), .B(KEYINPUT59), .Z(n965) );
  XNOR2_X1 U1060 ( .A(G4), .B(n965), .ZN(n967) );
  XNOR2_X1 U1061 ( .A(G20), .B(G1956), .ZN(n966) );
  NOR2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n971) );
  XNOR2_X1 U1063 ( .A(G1341), .B(G19), .ZN(n969) );
  XNOR2_X1 U1064 ( .A(G6), .B(G1981), .ZN(n968) );
  NOR2_X1 U1065 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1067 ( .A(KEYINPUT60), .B(n972), .ZN(n973) );
  NOR2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n975) );
  XOR2_X1 U1069 ( .A(KEYINPUT61), .B(n975), .Z(n976) );
  NOR2_X1 U1070 ( .A1(G16), .A2(n976), .ZN(n980) );
  NAND2_X1 U1071 ( .A1(n1005), .A2(n977), .ZN(n978) );
  NOR2_X1 U1072 ( .A1(G29), .A2(n978), .ZN(n979) );
  NOR2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n1009) );
  XOR2_X1 U1074 ( .A(G164), .B(G2078), .Z(n984) );
  XOR2_X1 U1075 ( .A(n981), .B(KEYINPUT120), .Z(n982) );
  XNOR2_X1 U1076 ( .A(G2072), .B(n982), .ZN(n983) );
  NOR2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1078 ( .A(KEYINPUT50), .B(n985), .ZN(n990) );
  XOR2_X1 U1079 ( .A(G2090), .B(G162), .Z(n986) );
  NOR2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1081 ( .A(KEYINPUT51), .B(n988), .Z(n989) );
  NAND2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n991) );
  NOR2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n1002) );
  NOR2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n998) );
  XOR2_X1 U1085 ( .A(G2084), .B(G160), .Z(n995) );
  NOR2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1090 ( .A(KEYINPUT121), .B(n1003), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(KEYINPUT52), .B(n1004), .ZN(n1006) );
  NAND2_X1 U1092 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1093 ( .A1(n1007), .A2(G29), .ZN(n1008) );
  NAND2_X1 U1094 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NOR2_X1 U1095 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1096 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1097 ( .A(n1014), .B(KEYINPUT126), .ZN(n1015) );
  XOR2_X1 U1098 ( .A(KEYINPUT62), .B(n1015), .Z(G311) );
  INV_X1 U1099 ( .A(G311), .ZN(G150) );
endmodule

