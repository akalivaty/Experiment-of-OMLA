

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U550 ( .A1(G651), .A2(n625), .ZN(n643) );
  NOR2_X1 U551 ( .A1(G2104), .A2(G2105), .ZN(n534) );
  OR2_X1 U552 ( .A1(n719), .A2(n718), .ZN(n517) );
  NAND2_X2 U553 ( .A1(n762), .A2(n760), .ZN(n687) );
  OR2_X1 U554 ( .A1(n726), .A2(n725), .ZN(n732) );
  BUF_X1 U555 ( .A(n693), .Z(n570) );
  AND2_X1 U556 ( .A1(G160), .A2(G40), .ZN(n760) );
  NOR2_X4 U557 ( .A1(n536), .A2(G2105), .ZN(n1000) );
  XOR2_X1 U558 ( .A(G543), .B(KEYINPUT0), .Z(n518) );
  XOR2_X1 U559 ( .A(KEYINPUT30), .B(n720), .Z(n519) );
  INV_X1 U560 ( .A(KEYINPUT26), .ZN(n688) );
  XNOR2_X1 U561 ( .A(KEYINPUT100), .B(KEYINPUT28), .ZN(n707) );
  XNOR2_X1 U562 ( .A(n708), .B(n707), .ZN(n709) );
  INV_X1 U563 ( .A(KEYINPUT103), .ZN(n733) );
  XNOR2_X1 U564 ( .A(n734), .B(n733), .ZN(n740) );
  INV_X1 U565 ( .A(KEYINPUT107), .ZN(n758) );
  XOR2_X1 U566 ( .A(KEYINPUT1), .B(n520), .Z(n644) );
  XNOR2_X1 U567 ( .A(n518), .B(KEYINPUT66), .ZN(n625) );
  NAND2_X1 U568 ( .A1(G53), .A2(n643), .ZN(n522) );
  INV_X1 U569 ( .A(G651), .ZN(n523) );
  NOR2_X1 U570 ( .A1(G543), .A2(n523), .ZN(n520) );
  NAND2_X1 U571 ( .A1(G65), .A2(n644), .ZN(n521) );
  NAND2_X1 U572 ( .A1(n522), .A2(n521), .ZN(n528) );
  NOR2_X2 U573 ( .A1(n625), .A2(n523), .ZN(n642) );
  NAND2_X1 U574 ( .A1(n642), .A2(G78), .ZN(n526) );
  NOR2_X1 U575 ( .A1(G651), .A2(G543), .ZN(n524) );
  XNOR2_X1 U576 ( .A(n524), .B(KEYINPUT64), .ZN(n647) );
  NAND2_X1 U577 ( .A1(G91), .A2(n647), .ZN(n525) );
  NAND2_X1 U578 ( .A1(n526), .A2(n525), .ZN(n527) );
  OR2_X1 U579 ( .A1(n528), .A2(n527), .ZN(G299) );
  INV_X1 U580 ( .A(G2105), .ZN(n535) );
  NOR2_X2 U581 ( .A1(n535), .A2(G2104), .ZN(n997) );
  NAND2_X1 U582 ( .A1(n997), .A2(G125), .ZN(n532) );
  INV_X1 U583 ( .A(G2104), .ZN(n536) );
  NAND2_X1 U584 ( .A1(n1000), .A2(G101), .ZN(n530) );
  INV_X1 U585 ( .A(KEYINPUT23), .ZN(n529) );
  XNOR2_X1 U586 ( .A(n530), .B(n529), .ZN(n531) );
  NAND2_X1 U587 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U588 ( .A(n533), .B(KEYINPUT65), .ZN(n540) );
  XOR2_X2 U589 ( .A(KEYINPUT17), .B(n534), .Z(n1001) );
  NAND2_X1 U590 ( .A1(G137), .A2(n1001), .ZN(n538) );
  NOR2_X1 U591 ( .A1(n536), .A2(n535), .ZN(n544) );
  NAND2_X1 U592 ( .A1(G113), .A2(n544), .ZN(n537) );
  AND2_X1 U593 ( .A1(n538), .A2(n537), .ZN(n539) );
  AND2_X1 U594 ( .A1(n540), .A2(n539), .ZN(G160) );
  AND2_X1 U595 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U596 ( .A1(n1001), .A2(G138), .ZN(n543) );
  NAND2_X1 U597 ( .A1(G102), .A2(n1000), .ZN(n541) );
  XOR2_X1 U598 ( .A(KEYINPUT91), .B(n541), .Z(n542) );
  NAND2_X1 U599 ( .A1(n543), .A2(n542), .ZN(n548) );
  NAND2_X1 U600 ( .A1(G114), .A2(n544), .ZN(n546) );
  NAND2_X1 U601 ( .A1(G126), .A2(n997), .ZN(n545) );
  NAND2_X1 U602 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U603 ( .A1(n548), .A2(n547), .ZN(G164) );
  INV_X1 U604 ( .A(G82), .ZN(G220) );
  INV_X1 U605 ( .A(G120), .ZN(G236) );
  INV_X1 U606 ( .A(G69), .ZN(G235) );
  NAND2_X1 U607 ( .A1(G64), .A2(n644), .ZN(n549) );
  XNOR2_X1 U608 ( .A(n549), .B(KEYINPUT67), .ZN(n556) );
  NAND2_X1 U609 ( .A1(n642), .A2(G77), .ZN(n551) );
  NAND2_X1 U610 ( .A1(G90), .A2(n647), .ZN(n550) );
  NAND2_X1 U611 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U612 ( .A(n552), .B(KEYINPUT9), .ZN(n554) );
  NAND2_X1 U613 ( .A1(G52), .A2(n643), .ZN(n553) );
  NAND2_X1 U614 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U615 ( .A1(n556), .A2(n555), .ZN(G171) );
  INV_X1 U616 ( .A(G171), .ZN(G301) );
  NAND2_X1 U617 ( .A1(G7), .A2(G661), .ZN(n557) );
  XNOR2_X1 U618 ( .A(n557), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U619 ( .A(G223), .B(KEYINPUT70), .Z(n830) );
  NAND2_X1 U620 ( .A1(n830), .A2(G567), .ZN(n558) );
  XOR2_X1 U621 ( .A(KEYINPUT11), .B(n558), .Z(G234) );
  INV_X1 U622 ( .A(G860), .ZN(n953) );
  NAND2_X1 U623 ( .A1(G43), .A2(n643), .ZN(n568) );
  NAND2_X1 U624 ( .A1(n644), .A2(G56), .ZN(n559) );
  XNOR2_X1 U625 ( .A(KEYINPUT14), .B(n559), .ZN(n565) );
  NAND2_X1 U626 ( .A1(G81), .A2(n647), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n560), .B(KEYINPUT12), .ZN(n562) );
  NAND2_X1 U628 ( .A1(G68), .A2(n642), .ZN(n561) );
  NAND2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(KEYINPUT13), .ZN(n564) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(KEYINPUT71), .ZN(n567) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(n569), .B(KEYINPUT72), .ZN(n693) );
  NOR2_X1 U635 ( .A1(n953), .A2(n570), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n571), .B(KEYINPUT73), .ZN(G153) );
  NAND2_X1 U637 ( .A1(G868), .A2(G301), .ZN(n581) );
  NAND2_X1 U638 ( .A1(G66), .A2(n644), .ZN(n573) );
  NAND2_X1 U639 ( .A1(G92), .A2(n647), .ZN(n572) );
  NAND2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n578) );
  NAND2_X1 U641 ( .A1(G54), .A2(n643), .ZN(n575) );
  NAND2_X1 U642 ( .A1(G79), .A2(n642), .ZN(n574) );
  NAND2_X1 U643 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U644 ( .A(KEYINPUT74), .B(n576), .ZN(n577) );
  NOR2_X1 U645 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n579), .B(KEYINPUT15), .ZN(n697) );
  INV_X1 U647 ( .A(G868), .ZN(n594) );
  NAND2_X1 U648 ( .A1(n697), .A2(n594), .ZN(n580) );
  NAND2_X1 U649 ( .A1(n581), .A2(n580), .ZN(G284) );
  NAND2_X1 U650 ( .A1(n642), .A2(G76), .ZN(n582) );
  XNOR2_X1 U651 ( .A(KEYINPUT76), .B(n582), .ZN(n586) );
  XOR2_X1 U652 ( .A(KEYINPUT75), .B(KEYINPUT4), .Z(n584) );
  NAND2_X1 U653 ( .A1(G89), .A2(n647), .ZN(n583) );
  XNOR2_X1 U654 ( .A(n584), .B(n583), .ZN(n585) );
  NAND2_X1 U655 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U656 ( .A(n587), .B(KEYINPUT5), .ZN(n592) );
  NAND2_X1 U657 ( .A1(G51), .A2(n643), .ZN(n589) );
  NAND2_X1 U658 ( .A1(G63), .A2(n644), .ZN(n588) );
  NAND2_X1 U659 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U660 ( .A(KEYINPUT6), .B(n590), .Z(n591) );
  NAND2_X1 U661 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U662 ( .A(n593), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U663 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U664 ( .A1(G286), .A2(n594), .ZN(n596) );
  NOR2_X1 U665 ( .A1(G868), .A2(G299), .ZN(n595) );
  NOR2_X1 U666 ( .A1(n596), .A2(n595), .ZN(G297) );
  NAND2_X1 U667 ( .A1(n953), .A2(G559), .ZN(n597) );
  INV_X1 U668 ( .A(n697), .ZN(n978) );
  NAND2_X1 U669 ( .A1(n597), .A2(n978), .ZN(n598) );
  XNOR2_X1 U670 ( .A(n598), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U671 ( .A1(n570), .A2(G868), .ZN(n601) );
  NAND2_X1 U672 ( .A1(G868), .A2(n978), .ZN(n599) );
  NOR2_X1 U673 ( .A1(G559), .A2(n599), .ZN(n600) );
  NOR2_X1 U674 ( .A1(n601), .A2(n600), .ZN(G282) );
  NAND2_X1 U675 ( .A1(G111), .A2(n544), .ZN(n608) );
  NAND2_X1 U676 ( .A1(G99), .A2(n1000), .ZN(n603) );
  NAND2_X1 U677 ( .A1(G135), .A2(n1001), .ZN(n602) );
  NAND2_X1 U678 ( .A1(n603), .A2(n602), .ZN(n606) );
  NAND2_X1 U679 ( .A1(n997), .A2(G123), .ZN(n604) );
  XOR2_X1 U680 ( .A(KEYINPUT18), .B(n604), .Z(n605) );
  NOR2_X1 U681 ( .A1(n606), .A2(n605), .ZN(n607) );
  NAND2_X1 U682 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U683 ( .A(n609), .B(KEYINPUT77), .ZN(n984) );
  XNOR2_X1 U684 ( .A(G2096), .B(n984), .ZN(n611) );
  INV_X1 U685 ( .A(G2100), .ZN(n610) );
  NAND2_X1 U686 ( .A1(n611), .A2(n610), .ZN(G156) );
  NAND2_X1 U687 ( .A1(G50), .A2(n643), .ZN(n613) );
  NAND2_X1 U688 ( .A1(G62), .A2(n644), .ZN(n612) );
  NAND2_X1 U689 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U690 ( .A(KEYINPUT84), .B(n614), .ZN(n619) );
  NAND2_X1 U691 ( .A1(n642), .A2(G75), .ZN(n616) );
  NAND2_X1 U692 ( .A1(G88), .A2(n647), .ZN(n615) );
  NAND2_X1 U693 ( .A1(n616), .A2(n615), .ZN(n617) );
  XOR2_X1 U694 ( .A(KEYINPUT85), .B(n617), .Z(n618) );
  NOR2_X1 U695 ( .A1(n619), .A2(n618), .ZN(G166) );
  NAND2_X1 U696 ( .A1(G49), .A2(n643), .ZN(n621) );
  NAND2_X1 U697 ( .A1(G74), .A2(G651), .ZN(n620) );
  NAND2_X1 U698 ( .A1(n621), .A2(n620), .ZN(n622) );
  XOR2_X1 U699 ( .A(KEYINPUT81), .B(n622), .Z(n623) );
  NOR2_X1 U700 ( .A1(n644), .A2(n623), .ZN(n624) );
  XNOR2_X1 U701 ( .A(n624), .B(KEYINPUT82), .ZN(n627) );
  NAND2_X1 U702 ( .A1(G87), .A2(n625), .ZN(n626) );
  NAND2_X1 U703 ( .A1(n627), .A2(n626), .ZN(n628) );
  XOR2_X1 U704 ( .A(KEYINPUT83), .B(n628), .Z(G288) );
  NAND2_X1 U705 ( .A1(G61), .A2(n644), .ZN(n630) );
  NAND2_X1 U706 ( .A1(G86), .A2(n647), .ZN(n629) );
  NAND2_X1 U707 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U708 ( .A1(n642), .A2(G73), .ZN(n631) );
  XOR2_X1 U709 ( .A(KEYINPUT2), .B(n631), .Z(n632) );
  NOR2_X1 U710 ( .A1(n633), .A2(n632), .ZN(n635) );
  NAND2_X1 U711 ( .A1(n643), .A2(G48), .ZN(n634) );
  NAND2_X1 U712 ( .A1(n635), .A2(n634), .ZN(G305) );
  AND2_X1 U713 ( .A1(n644), .A2(G60), .ZN(n639) );
  NAND2_X1 U714 ( .A1(G47), .A2(n643), .ZN(n637) );
  NAND2_X1 U715 ( .A1(G85), .A2(n647), .ZN(n636) );
  NAND2_X1 U716 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U717 ( .A1(n639), .A2(n638), .ZN(n641) );
  NAND2_X1 U718 ( .A1(n642), .A2(G72), .ZN(n640) );
  NAND2_X1 U719 ( .A1(n641), .A2(n640), .ZN(G290) );
  NAND2_X1 U720 ( .A1(n642), .A2(G80), .ZN(n652) );
  NAND2_X1 U721 ( .A1(G55), .A2(n643), .ZN(n646) );
  NAND2_X1 U722 ( .A1(G67), .A2(n644), .ZN(n645) );
  NAND2_X1 U723 ( .A1(n646), .A2(n645), .ZN(n650) );
  NAND2_X1 U724 ( .A1(G93), .A2(n647), .ZN(n648) );
  XNOR2_X1 U725 ( .A(KEYINPUT79), .B(n648), .ZN(n649) );
  NOR2_X1 U726 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U727 ( .A1(n652), .A2(n651), .ZN(n653) );
  XOR2_X1 U728 ( .A(KEYINPUT80), .B(n653), .Z(n956) );
  NOR2_X1 U729 ( .A1(G868), .A2(n956), .ZN(n654) );
  XOR2_X1 U730 ( .A(KEYINPUT88), .B(n654), .Z(n665) );
  XNOR2_X1 U731 ( .A(G166), .B(G288), .ZN(n660) );
  XOR2_X1 U732 ( .A(KEYINPUT19), .B(n956), .Z(n656) );
  XNOR2_X1 U733 ( .A(G299), .B(KEYINPUT86), .ZN(n655) );
  XNOR2_X1 U734 ( .A(n656), .B(n655), .ZN(n657) );
  XOR2_X1 U735 ( .A(n657), .B(G290), .Z(n658) );
  XNOR2_X1 U736 ( .A(G305), .B(n658), .ZN(n659) );
  XNOR2_X1 U737 ( .A(n660), .B(n659), .ZN(n977) );
  NAND2_X1 U738 ( .A1(G559), .A2(n978), .ZN(n661) );
  XOR2_X1 U739 ( .A(n570), .B(n661), .Z(n952) );
  XNOR2_X1 U740 ( .A(n977), .B(n952), .ZN(n662) );
  NAND2_X1 U741 ( .A1(n662), .A2(G868), .ZN(n663) );
  XOR2_X1 U742 ( .A(KEYINPUT87), .B(n663), .Z(n664) );
  NAND2_X1 U743 ( .A1(n665), .A2(n664), .ZN(G295) );
  NAND2_X1 U744 ( .A1(G2078), .A2(G2084), .ZN(n666) );
  XNOR2_X1 U745 ( .A(n666), .B(KEYINPUT89), .ZN(n667) );
  XNOR2_X1 U746 ( .A(n667), .B(KEYINPUT20), .ZN(n668) );
  NAND2_X1 U747 ( .A1(n668), .A2(G2090), .ZN(n669) );
  XNOR2_X1 U748 ( .A(KEYINPUT21), .B(n669), .ZN(n670) );
  NAND2_X1 U749 ( .A1(n670), .A2(G2072), .ZN(G158) );
  XOR2_X1 U750 ( .A(KEYINPUT68), .B(G57), .Z(G237) );
  XNOR2_X1 U751 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U752 ( .A(KEYINPUT69), .B(G132), .ZN(G219) );
  NOR2_X1 U753 ( .A1(G235), .A2(G236), .ZN(n671) );
  XOR2_X1 U754 ( .A(KEYINPUT90), .B(n671), .Z(n672) );
  NOR2_X1 U755 ( .A1(G237), .A2(n672), .ZN(n673) );
  NAND2_X1 U756 ( .A1(G108), .A2(n673), .ZN(n950) );
  NAND2_X1 U757 ( .A1(n950), .A2(G567), .ZN(n678) );
  NOR2_X1 U758 ( .A1(G220), .A2(G219), .ZN(n674) );
  XOR2_X1 U759 ( .A(KEYINPUT22), .B(n674), .Z(n675) );
  NOR2_X1 U760 ( .A1(G218), .A2(n675), .ZN(n676) );
  NAND2_X1 U761 ( .A1(G96), .A2(n676), .ZN(n951) );
  NAND2_X1 U762 ( .A1(n951), .A2(G2106), .ZN(n677) );
  NAND2_X1 U763 ( .A1(n678), .A2(n677), .ZN(n957) );
  NAND2_X1 U764 ( .A1(G483), .A2(G661), .ZN(n679) );
  NOR2_X1 U765 ( .A1(n957), .A2(n679), .ZN(n833) );
  NAND2_X1 U766 ( .A1(n833), .A2(G36), .ZN(G176) );
  INV_X1 U767 ( .A(G166), .ZN(G303) );
  NOR2_X1 U768 ( .A1(G164), .A2(G1384), .ZN(n762) );
  NOR2_X1 U769 ( .A1(G2084), .A2(n687), .ZN(n682) );
  XOR2_X1 U770 ( .A(KEYINPUT97), .B(n682), .Z(n718) );
  NAND2_X1 U771 ( .A1(G8), .A2(n718), .ZN(n683) );
  XOR2_X1 U772 ( .A(KEYINPUT98), .B(n683), .Z(n731) );
  NAND2_X1 U773 ( .A1(G8), .A2(n687), .ZN(n803) );
  NOR2_X1 U774 ( .A1(G1966), .A2(n803), .ZN(n728) );
  NAND2_X1 U775 ( .A1(G1348), .A2(n687), .ZN(n685) );
  INV_X1 U776 ( .A(n687), .ZN(n713) );
  NAND2_X1 U777 ( .A1(G2067), .A2(n713), .ZN(n684) );
  NAND2_X1 U778 ( .A1(n685), .A2(n684), .ZN(n696) );
  NOR2_X1 U779 ( .A1(n697), .A2(n696), .ZN(n695) );
  INV_X1 U780 ( .A(G1996), .ZN(n686) );
  NOR2_X1 U781 ( .A1(n687), .A2(n686), .ZN(n689) );
  XNOR2_X1 U782 ( .A(n689), .B(n688), .ZN(n691) );
  NAND2_X1 U783 ( .A1(n687), .A2(G1341), .ZN(n690) );
  NAND2_X1 U784 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U785 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U786 ( .A1(n695), .A2(n694), .ZN(n699) );
  AND2_X1 U787 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U788 ( .A1(n699), .A2(n698), .ZN(n704) );
  NAND2_X1 U789 ( .A1(n713), .A2(G2072), .ZN(n700) );
  XOR2_X1 U790 ( .A(KEYINPUT27), .B(n700), .Z(n702) );
  NAND2_X1 U791 ( .A1(G1956), .A2(n687), .ZN(n701) );
  NAND2_X1 U792 ( .A1(n702), .A2(n701), .ZN(n706) );
  NOR2_X1 U793 ( .A1(n706), .A2(G299), .ZN(n703) );
  NOR2_X1 U794 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U795 ( .A(n705), .B(KEYINPUT101), .ZN(n710) );
  NAND2_X1 U796 ( .A1(n706), .A2(G299), .ZN(n708) );
  NAND2_X1 U797 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U798 ( .A(n711), .B(KEYINPUT29), .ZN(n717) );
  XNOR2_X1 U799 ( .A(G2078), .B(KEYINPUT25), .ZN(n712) );
  XNOR2_X1 U800 ( .A(n712), .B(KEYINPUT99), .ZN(n873) );
  NOR2_X1 U801 ( .A1(n873), .A2(n687), .ZN(n715) );
  NOR2_X1 U802 ( .A1(n713), .A2(G1961), .ZN(n714) );
  NOR2_X1 U803 ( .A1(n715), .A2(n714), .ZN(n721) );
  NOR2_X1 U804 ( .A1(G301), .A2(n721), .ZN(n716) );
  NOR2_X1 U805 ( .A1(n717), .A2(n716), .ZN(n726) );
  INV_X1 U806 ( .A(G8), .ZN(n719) );
  NOR2_X1 U807 ( .A1(n728), .A2(n517), .ZN(n720) );
  NOR2_X1 U808 ( .A1(G168), .A2(n519), .ZN(n723) );
  AND2_X1 U809 ( .A1(G301), .A2(n721), .ZN(n722) );
  NOR2_X1 U810 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U811 ( .A(n724), .B(KEYINPUT31), .ZN(n725) );
  INV_X1 U812 ( .A(n732), .ZN(n727) );
  NOR2_X1 U813 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U814 ( .A(KEYINPUT102), .B(n729), .Z(n730) );
  NOR2_X1 U815 ( .A1(n731), .A2(n730), .ZN(n744) );
  NAND2_X1 U816 ( .A1(n732), .A2(G286), .ZN(n734) );
  NOR2_X1 U817 ( .A1(G1971), .A2(n803), .ZN(n736) );
  NOR2_X1 U818 ( .A1(G2090), .A2(n687), .ZN(n735) );
  NOR2_X1 U819 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U820 ( .A1(n737), .A2(G303), .ZN(n738) );
  XNOR2_X1 U821 ( .A(KEYINPUT104), .B(n738), .ZN(n739) );
  NAND2_X1 U822 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U823 ( .A1(n741), .A2(G8), .ZN(n742) );
  XOR2_X1 U824 ( .A(KEYINPUT32), .B(n742), .Z(n743) );
  NOR2_X1 U825 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U826 ( .A(KEYINPUT105), .B(n745), .ZN(n798) );
  NOR2_X1 U827 ( .A1(G1976), .A2(G288), .ZN(n751) );
  NOR2_X1 U828 ( .A1(G1971), .A2(G303), .ZN(n746) );
  NOR2_X1 U829 ( .A1(n751), .A2(n746), .ZN(n916) );
  INV_X1 U830 ( .A(KEYINPUT33), .ZN(n747) );
  AND2_X1 U831 ( .A1(n916), .A2(n747), .ZN(n748) );
  AND2_X1 U832 ( .A1(n798), .A2(n748), .ZN(n757) );
  NAND2_X1 U833 ( .A1(G1976), .A2(G288), .ZN(n907) );
  INV_X1 U834 ( .A(n907), .ZN(n749) );
  NOR2_X1 U835 ( .A1(n749), .A2(n803), .ZN(n750) );
  OR2_X1 U836 ( .A1(KEYINPUT33), .A2(n750), .ZN(n755) );
  NAND2_X1 U837 ( .A1(KEYINPUT33), .A2(n751), .ZN(n752) );
  NOR2_X1 U838 ( .A1(n803), .A2(n752), .ZN(n753) );
  XOR2_X1 U839 ( .A(n753), .B(KEYINPUT106), .Z(n754) );
  NAND2_X1 U840 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U841 ( .A1(n757), .A2(n756), .ZN(n759) );
  XNOR2_X1 U842 ( .A(n759), .B(n758), .ZN(n795) );
  XOR2_X1 U843 ( .A(G1981), .B(G305), .Z(n897) );
  INV_X1 U844 ( .A(n760), .ZN(n761) );
  NOR2_X1 U845 ( .A1(n762), .A2(n761), .ZN(n816) );
  NAND2_X1 U846 ( .A1(G104), .A2(n1000), .ZN(n764) );
  NAND2_X1 U847 ( .A1(G140), .A2(n1001), .ZN(n763) );
  NAND2_X1 U848 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U849 ( .A(KEYINPUT34), .B(n765), .ZN(n772) );
  NAND2_X1 U850 ( .A1(n997), .A2(G128), .ZN(n766) );
  XNOR2_X1 U851 ( .A(n766), .B(KEYINPUT92), .ZN(n768) );
  NAND2_X1 U852 ( .A1(G116), .A2(n544), .ZN(n767) );
  NAND2_X1 U853 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U854 ( .A(KEYINPUT35), .B(n769), .ZN(n770) );
  XNOR2_X1 U855 ( .A(KEYINPUT93), .B(n770), .ZN(n771) );
  NOR2_X1 U856 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U857 ( .A(KEYINPUT36), .B(n773), .ZN(n1010) );
  XNOR2_X1 U858 ( .A(G2067), .B(KEYINPUT37), .ZN(n806) );
  NOR2_X1 U859 ( .A1(n1010), .A2(n806), .ZN(n868) );
  NAND2_X1 U860 ( .A1(n816), .A2(n868), .ZN(n813) );
  NAND2_X1 U861 ( .A1(G107), .A2(n544), .ZN(n775) );
  NAND2_X1 U862 ( .A1(G119), .A2(n997), .ZN(n774) );
  NAND2_X1 U863 ( .A1(n775), .A2(n774), .ZN(n778) );
  NAND2_X1 U864 ( .A1(n1001), .A2(G131), .ZN(n776) );
  XOR2_X1 U865 ( .A(KEYINPUT94), .B(n776), .Z(n777) );
  NOR2_X1 U866 ( .A1(n778), .A2(n777), .ZN(n780) );
  NAND2_X1 U867 ( .A1(n1000), .A2(G95), .ZN(n779) );
  NAND2_X1 U868 ( .A1(n780), .A2(n779), .ZN(n992) );
  NAND2_X1 U869 ( .A1(G1991), .A2(n992), .ZN(n789) );
  NAND2_X1 U870 ( .A1(G141), .A2(n1001), .ZN(n782) );
  NAND2_X1 U871 ( .A1(G117), .A2(n544), .ZN(n781) );
  NAND2_X1 U872 ( .A1(n782), .A2(n781), .ZN(n785) );
  NAND2_X1 U873 ( .A1(n1000), .A2(G105), .ZN(n783) );
  XOR2_X1 U874 ( .A(KEYINPUT38), .B(n783), .Z(n784) );
  NOR2_X1 U875 ( .A1(n785), .A2(n784), .ZN(n787) );
  NAND2_X1 U876 ( .A1(n997), .A2(G129), .ZN(n786) );
  NAND2_X1 U877 ( .A1(n787), .A2(n786), .ZN(n991) );
  NAND2_X1 U878 ( .A1(G1996), .A2(n991), .ZN(n788) );
  NAND2_X1 U879 ( .A1(n789), .A2(n788), .ZN(n843) );
  NAND2_X1 U880 ( .A1(n843), .A2(n816), .ZN(n790) );
  XNOR2_X1 U881 ( .A(n790), .B(KEYINPUT95), .ZN(n809) );
  INV_X1 U882 ( .A(n809), .ZN(n791) );
  NAND2_X1 U883 ( .A1(n813), .A2(n791), .ZN(n792) );
  XOR2_X1 U884 ( .A(n792), .B(KEYINPUT96), .Z(n805) );
  AND2_X1 U885 ( .A1(n897), .A2(n805), .ZN(n793) );
  XNOR2_X1 U886 ( .A(G1986), .B(G290), .ZN(n901) );
  NAND2_X1 U887 ( .A1(n901), .A2(n816), .ZN(n822) );
  AND2_X1 U888 ( .A1(n793), .A2(n822), .ZN(n794) );
  NAND2_X1 U889 ( .A1(n795), .A2(n794), .ZN(n828) );
  NOR2_X1 U890 ( .A1(G2090), .A2(G303), .ZN(n796) );
  NAND2_X1 U891 ( .A1(G8), .A2(n796), .ZN(n797) );
  NAND2_X1 U892 ( .A1(n798), .A2(n797), .ZN(n800) );
  AND2_X1 U893 ( .A1(n803), .A2(n805), .ZN(n799) );
  AND2_X1 U894 ( .A1(n800), .A2(n799), .ZN(n821) );
  NOR2_X1 U895 ( .A1(G1981), .A2(G305), .ZN(n801) );
  XOR2_X1 U896 ( .A(n801), .B(KEYINPUT24), .Z(n802) );
  NOR2_X1 U897 ( .A1(n803), .A2(n802), .ZN(n804) );
  AND2_X1 U898 ( .A1(n805), .A2(n804), .ZN(n819) );
  NAND2_X1 U899 ( .A1(n1010), .A2(n806), .ZN(n865) );
  NOR2_X1 U900 ( .A1(G1996), .A2(n991), .ZN(n848) );
  NOR2_X1 U901 ( .A1(G1991), .A2(n992), .ZN(n844) );
  NOR2_X1 U902 ( .A1(G1986), .A2(G290), .ZN(n807) );
  NOR2_X1 U903 ( .A1(n844), .A2(n807), .ZN(n808) );
  NOR2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U905 ( .A1(n848), .A2(n810), .ZN(n811) );
  XNOR2_X1 U906 ( .A(KEYINPUT39), .B(n811), .ZN(n812) );
  XNOR2_X1 U907 ( .A(n812), .B(KEYINPUT108), .ZN(n814) );
  NAND2_X1 U908 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U909 ( .A1(n865), .A2(n815), .ZN(n817) );
  NAND2_X1 U910 ( .A1(n817), .A2(n816), .ZN(n824) );
  INV_X1 U911 ( .A(n824), .ZN(n818) );
  OR2_X1 U912 ( .A1(n819), .A2(n818), .ZN(n820) );
  NOR2_X1 U913 ( .A1(n821), .A2(n820), .ZN(n826) );
  INV_X1 U914 ( .A(n822), .ZN(n823) );
  AND2_X1 U915 ( .A1(n824), .A2(n823), .ZN(n825) );
  OR2_X1 U916 ( .A1(n826), .A2(n825), .ZN(n827) );
  NAND2_X1 U917 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U918 ( .A(n829), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U919 ( .A1(G2106), .A2(n830), .ZN(G217) );
  AND2_X1 U920 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U921 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U923 ( .A1(n833), .A2(n832), .ZN(G188) );
  XNOR2_X1 U924 ( .A(G96), .B(KEYINPUT109), .ZN(G221) );
  NAND2_X1 U926 ( .A1(n544), .A2(G112), .ZN(n840) );
  NAND2_X1 U927 ( .A1(G100), .A2(n1000), .ZN(n835) );
  NAND2_X1 U928 ( .A1(G136), .A2(n1001), .ZN(n834) );
  NAND2_X1 U929 ( .A1(n835), .A2(n834), .ZN(n838) );
  NAND2_X1 U930 ( .A1(n997), .A2(G124), .ZN(n836) );
  XOR2_X1 U931 ( .A(KEYINPUT44), .B(n836), .Z(n837) );
  NOR2_X1 U932 ( .A1(n838), .A2(n837), .ZN(n839) );
  NAND2_X1 U933 ( .A1(n840), .A2(n839), .ZN(n841) );
  XOR2_X1 U934 ( .A(KEYINPUT112), .B(n841), .Z(G162) );
  INV_X1 U935 ( .A(KEYINPUT55), .ZN(n893) );
  XNOR2_X1 U936 ( .A(KEYINPUT120), .B(KEYINPUT52), .ZN(n870) );
  XOR2_X1 U937 ( .A(G2084), .B(G160), .Z(n842) );
  NOR2_X1 U938 ( .A1(n984), .A2(n842), .ZN(n846) );
  NOR2_X1 U939 ( .A1(n844), .A2(n843), .ZN(n845) );
  NAND2_X1 U940 ( .A1(n846), .A2(n845), .ZN(n864) );
  XOR2_X1 U941 ( .A(G2090), .B(G162), .Z(n847) );
  NOR2_X1 U942 ( .A1(n848), .A2(n847), .ZN(n849) );
  XOR2_X1 U943 ( .A(KEYINPUT51), .B(n849), .Z(n862) );
  NAND2_X1 U944 ( .A1(G115), .A2(n544), .ZN(n851) );
  NAND2_X1 U945 ( .A1(G127), .A2(n997), .ZN(n850) );
  NAND2_X1 U946 ( .A1(n851), .A2(n850), .ZN(n852) );
  XNOR2_X1 U947 ( .A(n852), .B(KEYINPUT47), .ZN(n854) );
  NAND2_X1 U948 ( .A1(G103), .A2(n1000), .ZN(n853) );
  NAND2_X1 U949 ( .A1(n854), .A2(n853), .ZN(n857) );
  NAND2_X1 U950 ( .A1(n1001), .A2(G139), .ZN(n855) );
  XOR2_X1 U951 ( .A(KEYINPUT116), .B(n855), .Z(n856) );
  NOR2_X1 U952 ( .A1(n857), .A2(n856), .ZN(n985) );
  XOR2_X1 U953 ( .A(G2072), .B(n985), .Z(n859) );
  XOR2_X1 U954 ( .A(G164), .B(G2078), .Z(n858) );
  NOR2_X1 U955 ( .A1(n859), .A2(n858), .ZN(n860) );
  XNOR2_X1 U956 ( .A(KEYINPUT50), .B(n860), .ZN(n861) );
  NAND2_X1 U957 ( .A1(n862), .A2(n861), .ZN(n863) );
  NOR2_X1 U958 ( .A1(n864), .A2(n863), .ZN(n866) );
  NAND2_X1 U959 ( .A1(n866), .A2(n865), .ZN(n867) );
  NOR2_X1 U960 ( .A1(n868), .A2(n867), .ZN(n869) );
  XNOR2_X1 U961 ( .A(n870), .B(n869), .ZN(n871) );
  NAND2_X1 U962 ( .A1(n893), .A2(n871), .ZN(n872) );
  NAND2_X1 U963 ( .A1(n872), .A2(G29), .ZN(n948) );
  XNOR2_X1 U964 ( .A(G2090), .B(G35), .ZN(n888) );
  XNOR2_X1 U965 ( .A(G1996), .B(G32), .ZN(n875) );
  XNOR2_X1 U966 ( .A(n873), .B(G27), .ZN(n874) );
  NOR2_X1 U967 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U968 ( .A(KEYINPUT122), .B(n876), .ZN(n880) );
  XNOR2_X1 U969 ( .A(G2067), .B(G26), .ZN(n878) );
  XNOR2_X1 U970 ( .A(G33), .B(G2072), .ZN(n877) );
  NOR2_X1 U971 ( .A1(n878), .A2(n877), .ZN(n879) );
  NAND2_X1 U972 ( .A1(n880), .A2(n879), .ZN(n881) );
  XNOR2_X1 U973 ( .A(KEYINPUT123), .B(n881), .ZN(n882) );
  NAND2_X1 U974 ( .A1(n882), .A2(G28), .ZN(n885) );
  XOR2_X1 U975 ( .A(G25), .B(G1991), .Z(n883) );
  XNOR2_X1 U976 ( .A(KEYINPUT121), .B(n883), .ZN(n884) );
  NOR2_X1 U977 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U978 ( .A(KEYINPUT53), .B(n886), .ZN(n887) );
  NOR2_X1 U979 ( .A1(n888), .A2(n887), .ZN(n891) );
  XOR2_X1 U980 ( .A(G2084), .B(G34), .Z(n889) );
  XNOR2_X1 U981 ( .A(KEYINPUT54), .B(n889), .ZN(n890) );
  NAND2_X1 U982 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U983 ( .A(n893), .B(n892), .ZN(n895) );
  INV_X1 U984 ( .A(G29), .ZN(n894) );
  NAND2_X1 U985 ( .A1(n895), .A2(n894), .ZN(n896) );
  NAND2_X1 U986 ( .A1(G11), .A2(n896), .ZN(n946) );
  XNOR2_X1 U987 ( .A(G16), .B(KEYINPUT56), .ZN(n918) );
  XNOR2_X1 U988 ( .A(G1966), .B(G168), .ZN(n898) );
  NAND2_X1 U989 ( .A1(n898), .A2(n897), .ZN(n899) );
  XNOR2_X1 U990 ( .A(n899), .B(KEYINPUT57), .ZN(n912) );
  XNOR2_X1 U991 ( .A(G1956), .B(G299), .ZN(n900) );
  NOR2_X1 U992 ( .A1(n901), .A2(n900), .ZN(n903) );
  NAND2_X1 U993 ( .A1(G1971), .A2(G303), .ZN(n902) );
  NAND2_X1 U994 ( .A1(n903), .A2(n902), .ZN(n906) );
  XOR2_X1 U995 ( .A(G1348), .B(n978), .Z(n904) );
  XNOR2_X1 U996 ( .A(KEYINPUT124), .B(n904), .ZN(n905) );
  NOR2_X1 U997 ( .A1(n906), .A2(n905), .ZN(n908) );
  NAND2_X1 U998 ( .A1(n908), .A2(n907), .ZN(n910) );
  XNOR2_X1 U999 ( .A(G1961), .B(G301), .ZN(n909) );
  NOR2_X1 U1000 ( .A1(n910), .A2(n909), .ZN(n911) );
  NAND2_X1 U1001 ( .A1(n912), .A2(n911), .ZN(n914) );
  XNOR2_X1 U1002 ( .A(G1341), .B(n570), .ZN(n913) );
  NOR2_X1 U1003 ( .A1(n914), .A2(n913), .ZN(n915) );
  NAND2_X1 U1004 ( .A1(n916), .A2(n915), .ZN(n917) );
  NAND2_X1 U1005 ( .A1(n918), .A2(n917), .ZN(n944) );
  INV_X1 U1006 ( .A(G16), .ZN(n942) );
  XNOR2_X1 U1007 ( .A(G1348), .B(KEYINPUT59), .ZN(n919) );
  XNOR2_X1 U1008 ( .A(n919), .B(G4), .ZN(n923) );
  XNOR2_X1 U1009 ( .A(G1956), .B(G20), .ZN(n921) );
  XNOR2_X1 U1010 ( .A(G19), .B(G1341), .ZN(n920) );
  NOR2_X1 U1011 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1012 ( .A1(n923), .A2(n922), .ZN(n926) );
  XOR2_X1 U1013 ( .A(KEYINPUT125), .B(G1981), .Z(n924) );
  XNOR2_X1 U1014 ( .A(G6), .B(n924), .ZN(n925) );
  NOR2_X1 U1015 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1016 ( .A(KEYINPUT60), .B(n927), .ZN(n931) );
  XNOR2_X1 U1017 ( .A(G1966), .B(G21), .ZN(n929) );
  XNOR2_X1 U1018 ( .A(G5), .B(G1961), .ZN(n928) );
  NOR2_X1 U1019 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1020 ( .A1(n931), .A2(n930), .ZN(n939) );
  XNOR2_X1 U1021 ( .A(G1986), .B(G24), .ZN(n933) );
  XNOR2_X1 U1022 ( .A(G1971), .B(G22), .ZN(n932) );
  NOR2_X1 U1023 ( .A1(n933), .A2(n932), .ZN(n936) );
  XOR2_X1 U1024 ( .A(G1976), .B(KEYINPUT126), .Z(n934) );
  XNOR2_X1 U1025 ( .A(G23), .B(n934), .ZN(n935) );
  NAND2_X1 U1026 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1027 ( .A(KEYINPUT58), .B(n937), .ZN(n938) );
  NOR2_X1 U1028 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1029 ( .A(KEYINPUT61), .B(n940), .ZN(n941) );
  NAND2_X1 U1030 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1031 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1032 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1033 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1034 ( .A(KEYINPUT62), .B(n949), .Z(G311) );
  XNOR2_X1 U1035 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1036 ( .A(G108), .ZN(G238) );
  NOR2_X1 U1037 ( .A1(n951), .A2(n950), .ZN(G325) );
  INV_X1 U1038 ( .A(G325), .ZN(G261) );
  NAND2_X1 U1039 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1040 ( .A(n954), .B(KEYINPUT78), .ZN(n955) );
  XOR2_X1 U1041 ( .A(n956), .B(n955), .Z(G145) );
  INV_X1 U1042 ( .A(n957), .ZN(G319) );
  XOR2_X1 U1043 ( .A(G2096), .B(G2678), .Z(n959) );
  XNOR2_X1 U1044 ( .A(G2067), .B(G2072), .ZN(n958) );
  XNOR2_X1 U1045 ( .A(n959), .B(n958), .ZN(n960) );
  XOR2_X1 U1046 ( .A(n960), .B(KEYINPUT42), .Z(n962) );
  XNOR2_X1 U1047 ( .A(G2090), .B(KEYINPUT43), .ZN(n961) );
  XNOR2_X1 U1048 ( .A(n962), .B(n961), .ZN(n966) );
  XOR2_X1 U1049 ( .A(KEYINPUT110), .B(G2100), .Z(n964) );
  XNOR2_X1 U1050 ( .A(G2078), .B(G2084), .ZN(n963) );
  XNOR2_X1 U1051 ( .A(n964), .B(n963), .ZN(n965) );
  XNOR2_X1 U1052 ( .A(n966), .B(n965), .ZN(G227) );
  XOR2_X1 U1053 ( .A(G1981), .B(G1971), .Z(n968) );
  XNOR2_X1 U1054 ( .A(G1961), .B(G1956), .ZN(n967) );
  XNOR2_X1 U1055 ( .A(n968), .B(n967), .ZN(n972) );
  XOR2_X1 U1056 ( .A(KEYINPUT111), .B(G2474), .Z(n970) );
  XNOR2_X1 U1057 ( .A(G1996), .B(G1991), .ZN(n969) );
  XNOR2_X1 U1058 ( .A(n970), .B(n969), .ZN(n971) );
  XOR2_X1 U1059 ( .A(n972), .B(n971), .Z(n974) );
  XNOR2_X1 U1060 ( .A(G1976), .B(KEYINPUT41), .ZN(n973) );
  XNOR2_X1 U1061 ( .A(n974), .B(n973), .ZN(n976) );
  XOR2_X1 U1062 ( .A(G1986), .B(G1966), .Z(n975) );
  XNOR2_X1 U1063 ( .A(n976), .B(n975), .ZN(G229) );
  XOR2_X1 U1064 ( .A(KEYINPUT119), .B(n977), .Z(n980) );
  XNOR2_X1 U1065 ( .A(G171), .B(n978), .ZN(n979) );
  XNOR2_X1 U1066 ( .A(n980), .B(n979), .ZN(n982) );
  XNOR2_X1 U1067 ( .A(G286), .B(n570), .ZN(n981) );
  XNOR2_X1 U1068 ( .A(n982), .B(n981), .ZN(n983) );
  NOR2_X1 U1069 ( .A1(G37), .A2(n983), .ZN(G397) );
  XOR2_X1 U1070 ( .A(n985), .B(n984), .Z(n986) );
  XNOR2_X1 U1071 ( .A(G162), .B(n986), .ZN(n990) );
  XOR2_X1 U1072 ( .A(KEYINPUT115), .B(KEYINPUT46), .Z(n988) );
  XNOR2_X1 U1073 ( .A(KEYINPUT48), .B(KEYINPUT117), .ZN(n987) );
  XNOR2_X1 U1074 ( .A(n988), .B(n987), .ZN(n989) );
  XOR2_X1 U1075 ( .A(n990), .B(n989), .Z(n996) );
  XNOR2_X1 U1076 ( .A(G160), .B(n991), .ZN(n993) );
  XNOR2_X1 U1077 ( .A(n993), .B(n992), .ZN(n994) );
  XNOR2_X1 U1078 ( .A(G164), .B(n994), .ZN(n995) );
  XNOR2_X1 U1079 ( .A(n996), .B(n995), .ZN(n1012) );
  NAND2_X1 U1080 ( .A1(G118), .A2(n544), .ZN(n999) );
  NAND2_X1 U1081 ( .A1(G130), .A2(n997), .ZN(n998) );
  NAND2_X1 U1082 ( .A1(n999), .A2(n998), .ZN(n1008) );
  XNOR2_X1 U1083 ( .A(KEYINPUT45), .B(KEYINPUT114), .ZN(n1006) );
  NAND2_X1 U1084 ( .A1(n1000), .A2(G106), .ZN(n1004) );
  NAND2_X1 U1085 ( .A1(n1001), .A2(G142), .ZN(n1002) );
  XOR2_X1 U1086 ( .A(KEYINPUT113), .B(n1002), .Z(n1003) );
  NAND2_X1 U1087 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1088 ( .A(n1006), .B(n1005), .Z(n1007) );
  NOR2_X1 U1089 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1090 ( .A(n1010), .B(n1009), .Z(n1011) );
  XNOR2_X1 U1091 ( .A(n1012), .B(n1011), .ZN(n1013) );
  NOR2_X1 U1092 ( .A1(G37), .A2(n1013), .ZN(n1014) );
  XNOR2_X1 U1093 ( .A(KEYINPUT118), .B(n1014), .ZN(G395) );
  XOR2_X1 U1094 ( .A(G2446), .B(G2451), .Z(n1016) );
  XNOR2_X1 U1095 ( .A(G1341), .B(G2430), .ZN(n1015) );
  XNOR2_X1 U1096 ( .A(n1016), .B(n1015), .ZN(n1022) );
  XOR2_X1 U1097 ( .A(G2443), .B(G2438), .Z(n1018) );
  XNOR2_X1 U1098 ( .A(G2454), .B(G2435), .ZN(n1017) );
  XNOR2_X1 U1099 ( .A(n1018), .B(n1017), .ZN(n1020) );
  XOR2_X1 U1100 ( .A(G1348), .B(G2427), .Z(n1019) );
  XNOR2_X1 U1101 ( .A(n1020), .B(n1019), .ZN(n1021) );
  XOR2_X1 U1102 ( .A(n1022), .B(n1021), .Z(n1023) );
  NAND2_X1 U1103 ( .A1(G14), .A2(n1023), .ZN(n1029) );
  NAND2_X1 U1104 ( .A1(G319), .A2(n1029), .ZN(n1026) );
  NOR2_X1 U1105 ( .A1(G227), .A2(G229), .ZN(n1024) );
  XNOR2_X1 U1106 ( .A(KEYINPUT49), .B(n1024), .ZN(n1025) );
  NOR2_X1 U1107 ( .A1(n1026), .A2(n1025), .ZN(n1028) );
  NOR2_X1 U1108 ( .A1(G397), .A2(G395), .ZN(n1027) );
  NAND2_X1 U1109 ( .A1(n1028), .A2(n1027), .ZN(G225) );
  INV_X1 U1110 ( .A(G225), .ZN(G308) );
  INV_X1 U1111 ( .A(n1029), .ZN(G401) );
endmodule

