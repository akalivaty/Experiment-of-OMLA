//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 1 0 1 1 1 0 1 1 0 1 1 1 0 1 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 0 0 0 0 1 0 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:01 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n566,
    new_n568, new_n569, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1203, new_n1204, new_n1205;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT65), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  XNOR2_X1  g030(.A(G325), .B(KEYINPUT66), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT67), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(new_n453), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT68), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT69), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n462), .A2(new_n463), .A3(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  AOI21_X1  g040(.A(KEYINPUT69), .B1(new_n465), .B2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n465), .A2(G2104), .ZN(new_n467));
  OAI211_X1 g042(.A(G137), .B(new_n464), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G101), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n465), .A2(G2104), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n472), .A2(new_n473), .A3(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n471), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n470), .A2(new_n476), .ZN(G160));
  OAI21_X1  g052(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(KEYINPUT70), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(new_n464), .C1(new_n466), .C2(new_n467), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(new_n471), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n482), .A2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n484), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  NAND4_X1  g065(.A1(new_n472), .A2(new_n473), .A3(G138), .A4(new_n471), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n471), .A2(G102), .A3(G2104), .ZN(new_n494));
  AND3_X1   g069(.A1(new_n471), .A2(KEYINPUT4), .A3(G138), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n495), .B(new_n464), .C1(new_n466), .C2(new_n467), .ZN(new_n496));
  AND3_X1   g071(.A1(new_n493), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  OAI211_X1 g072(.A(G126), .B(new_n464), .C1(new_n466), .C2(new_n467), .ZN(new_n498));
  NAND2_X1  g073(.A1(G114), .A2(G2104), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  INV_X1    g078(.A(KEYINPUT73), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(G543), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n505), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n504), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(KEYINPUT6), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  OAI21_X1  g091(.A(KEYINPUT71), .B1(new_n516), .B2(G651), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT71), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n518), .A2(new_n513), .A3(KEYINPUT6), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n515), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n520), .A2(new_n511), .A3(G88), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n520), .A2(G50), .A3(G543), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n508), .A2(G543), .ZN(new_n524));
  AND3_X1   g099(.A1(new_n505), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n525));
  AOI21_X1  g100(.A(KEYINPUT72), .B1(new_n505), .B2(KEYINPUT5), .ZN(new_n526));
  OAI211_X1 g101(.A(G62), .B(new_n524), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(G75), .A2(G543), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n529), .A2(KEYINPUT73), .A3(G651), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n514), .A2(new_n523), .A3(new_n530), .ZN(G303));
  INV_X1    g106(.A(G303), .ZN(G166));
  NAND2_X1  g107(.A1(new_n520), .A2(new_n511), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G89), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n520), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G51), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT7), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n535), .A2(new_n538), .A3(new_n539), .A4(new_n541), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  INV_X1    g118(.A(KEYINPUT74), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n520), .A2(new_n511), .A3(G90), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n520), .A2(G52), .A3(G543), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI211_X1 g122(.A(G64), .B(new_n524), .C1(new_n525), .C2(new_n526), .ZN(new_n548));
  NAND2_X1  g123(.A1(G77), .A2(G543), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n513), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n544), .B1(new_n547), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NOR3_X1   g127(.A1(new_n547), .A2(new_n550), .A3(new_n544), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n552), .A2(new_n553), .ZN(G301));
  INV_X1    g129(.A(G301), .ZN(G171));
  INV_X1    g130(.A(G81), .ZN(new_n556));
  INV_X1    g131(.A(G43), .ZN(new_n557));
  OAI22_X1  g132(.A1(new_n556), .A2(new_n533), .B1(new_n536), .B2(new_n557), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT76), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n560));
  OR2_X1    g135(.A1(new_n560), .A2(KEYINPUT75), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(KEYINPUT75), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n561), .A2(G651), .A3(new_n562), .ZN(new_n563));
  AND2_X1   g138(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  AND3_X1   g140(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G36), .ZN(G176));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT8), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n566), .A2(new_n569), .ZN(G188));
  NAND3_X1  g145(.A1(new_n520), .A2(G53), .A3(G543), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT9), .ZN(new_n572));
  OAI211_X1 g147(.A(G65), .B(new_n524), .C1(new_n525), .C2(new_n526), .ZN(new_n573));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT77), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n573), .A2(KEYINPUT77), .A3(new_n574), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n577), .A2(G651), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n534), .A2(G91), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n572), .A2(new_n579), .A3(new_n580), .ZN(G299));
  INV_X1    g156(.A(KEYINPUT78), .ZN(new_n582));
  INV_X1    g157(.A(G87), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n533), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n520), .A2(G49), .A3(G543), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n520), .A2(new_n511), .A3(KEYINPUT78), .A4(G87), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n584), .A2(new_n585), .A3(new_n586), .A4(new_n587), .ZN(G288));
  NAND2_X1  g163(.A1(new_n511), .A2(G61), .ZN(new_n589));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n591), .A2(G651), .B1(new_n537), .B2(G48), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT79), .ZN(new_n593));
  INV_X1    g168(.A(G86), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n533), .B2(new_n594), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n520), .A2(new_n511), .A3(KEYINPUT79), .A4(G86), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n592), .A2(new_n597), .ZN(G305));
  INV_X1    g173(.A(G85), .ZN(new_n599));
  INV_X1    g174(.A(G47), .ZN(new_n600));
  OAI22_X1  g175(.A1(new_n599), .A2(new_n533), .B1(new_n536), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(new_n513), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  INV_X1    g181(.A(G92), .ZN(new_n607));
  OR3_X1    g182(.A1(new_n533), .A2(KEYINPUT10), .A3(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(KEYINPUT10), .B1(new_n533), .B2(new_n607), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g185(.A(KEYINPUT80), .B(G66), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n511), .A2(new_n611), .B1(G79), .B2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G54), .ZN(new_n613));
  OAI22_X1  g188(.A1(new_n612), .A2(new_n513), .B1(new_n613), .B2(new_n536), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n606), .B1(G868), .B2(new_n615), .ZN(G284));
  OAI21_X1  g191(.A(new_n606), .B1(G868), .B2(new_n615), .ZN(G321));
  NAND2_X1  g192(.A1(G286), .A2(G868), .ZN(new_n618));
  XOR2_X1   g193(.A(G299), .B(KEYINPUT81), .Z(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(G868), .ZN(G297));
  XNOR2_X1  g195(.A(G297), .B(KEYINPUT82), .ZN(G280));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n615), .B1(new_n622), .B2(G860), .ZN(G148));
  NAND2_X1  g198(.A1(new_n559), .A2(new_n563), .ZN(new_n624));
  INV_X1    g199(.A(G868), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(new_n615), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n627), .A2(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n626), .B1(new_n628), .B2(new_n625), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g205(.A1(new_n483), .A2(G123), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n485), .A2(G135), .ZN(new_n632));
  OAI21_X1  g207(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n633));
  INV_X1    g208(.A(KEYINPUT83), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n635), .B(new_n636), .C1(G111), .C2(new_n471), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n631), .A2(new_n632), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(G2096), .Z(new_n639));
  NAND3_X1  g214(.A1(new_n471), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT12), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT13), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(G2100), .Z(new_n643));
  NAND2_X1  g218(.A1(new_n639), .A2(new_n643), .ZN(G156));
  XOR2_X1   g219(.A(KEYINPUT15), .B(G2435), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2427), .B(G2430), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT84), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n646), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(KEYINPUT14), .ZN(new_n650));
  XOR2_X1   g225(.A(G2443), .B(G2446), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G1341), .B(G1348), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n652), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2451), .B(G2454), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(G14), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(G401));
  XNOR2_X1  g234(.A(G2084), .B(G2090), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT85), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2072), .B(G2078), .Z(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT86), .B(KEYINPUT18), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT88), .B(KEYINPUT17), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n664), .B(new_n668), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n669), .B1(new_n661), .B2(new_n662), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT87), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n662), .B1(new_n664), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n672), .B1(new_n671), .B2(new_n664), .ZN(new_n673));
  OAI211_X1 g248(.A(new_n670), .B(new_n663), .C1(new_n661), .C2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n667), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2096), .B(G2100), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(G227));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  NOR2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1971), .B(G1976), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT19), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n679), .A2(new_n680), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT20), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n685), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n682), .A2(new_n684), .A3(new_n686), .ZN(new_n690));
  OAI211_X1 g265(.A(new_n689), .B(new_n690), .C1(new_n688), .C2(new_n687), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1991), .B(G1996), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(G1981), .ZN(new_n695));
  INV_X1    g270(.A(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n693), .B(new_n697), .ZN(G229));
  INV_X1    g273(.A(KEYINPUT99), .ZN(new_n699));
  OAI21_X1  g274(.A(G16), .B1(new_n552), .B2(new_n553), .ZN(new_n700));
  NOR2_X1   g275(.A1(G5), .A2(G16), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n699), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n545), .A2(new_n546), .ZN(new_n705));
  INV_X1    g280(.A(new_n550), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n705), .A2(new_n706), .A3(KEYINPUT74), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n704), .B1(new_n707), .B2(new_n551), .ZN(new_n708));
  NOR3_X1   g283(.A1(new_n708), .A2(KEYINPUT99), .A3(new_n701), .ZN(new_n709));
  OAI21_X1  g284(.A(G1961), .B1(new_n703), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(KEYINPUT100), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT100), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n712), .B(G1961), .C1(new_n703), .C2(new_n709), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT28), .ZN(new_n715));
  INV_X1    g290(.A(G26), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(G29), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(G29), .ZN(new_n718));
  NAND4_X1  g293(.A1(new_n479), .A2(G140), .A3(new_n471), .A4(new_n481), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT93), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g296(.A1(new_n479), .A2(G128), .A3(G2105), .A4(new_n481), .ZN(new_n722));
  OR2_X1    g297(.A1(G104), .A2(G2105), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n723), .B(G2104), .C1(G116), .C2(new_n471), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n719), .A2(new_n720), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n721), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n718), .B1(new_n727), .B2(G29), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n717), .B1(new_n728), .B2(new_n715), .ZN(new_n729));
  INV_X1    g304(.A(G2067), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  OR2_X1    g306(.A1(G29), .A2(G32), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n483), .A2(G129), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n485), .A2(G141), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n471), .A2(G105), .A3(G2104), .ZN(new_n735));
  NAND3_X1  g310(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT26), .Z(new_n737));
  NAND4_X1  g312(.A1(new_n733), .A2(new_n734), .A3(new_n735), .A4(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G29), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n732), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT27), .B(G1996), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n489), .A2(G29), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n739), .A2(G35), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n745), .A2(KEYINPUT29), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n745), .A2(KEYINPUT29), .ZN(new_n747));
  OAI21_X1  g322(.A(G2090), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n714), .A2(new_n731), .A3(new_n742), .A4(new_n748), .ZN(new_n749));
  OR2_X1    g324(.A1(G16), .A2(G21), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G286), .B2(new_n704), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G1966), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n754), .A2(KEYINPUT97), .ZN(new_n755));
  NAND2_X1  g330(.A1(G299), .A2(G16), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n704), .A2(KEYINPUT23), .A3(G20), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT23), .ZN(new_n758));
  INV_X1    g333(.A(G20), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n759), .B2(G16), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n756), .A2(new_n757), .A3(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G1956), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(G27), .A2(G29), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G164), .B2(G29), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n765), .A2(G2078), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n754), .B2(KEYINPUT97), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n763), .B(new_n767), .C1(G1966), .C2(new_n752), .ZN(new_n768));
  NOR3_X1   g343(.A1(new_n703), .A2(new_n709), .A3(G1961), .ZN(new_n769));
  NOR4_X1   g344(.A1(new_n749), .A2(new_n755), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n704), .A2(G19), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n564), .B2(new_n704), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(G1341), .Z(new_n773));
  AND2_X1   g348(.A1(new_n704), .A2(G23), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G288), .B2(G16), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT33), .B(G1976), .Z(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  AOI211_X1 g353(.A(new_n776), .B(new_n774), .C1(G288), .C2(G16), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT90), .B(KEYINPUT91), .Z(new_n781));
  NAND3_X1  g356(.A1(new_n778), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  OR2_X1    g357(.A1(G16), .A2(G22), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G303), .B2(new_n704), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT92), .B(G1971), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(new_n781), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n775), .A2(new_n777), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(new_n779), .ZN(new_n789));
  AND3_X1   g364(.A1(new_n782), .A2(new_n786), .A3(new_n789), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT89), .B(G1981), .Z(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT32), .ZN(new_n793));
  NAND2_X1  g368(.A1(G305), .A2(G16), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n704), .A2(G6), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n793), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n704), .B1(new_n592), .B2(new_n597), .ZN(new_n797));
  INV_X1    g372(.A(new_n795), .ZN(new_n798));
  NOR3_X1   g373(.A1(new_n797), .A2(KEYINPUT32), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n792), .B1(new_n796), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n794), .A2(new_n793), .A3(new_n795), .ZN(new_n801));
  OAI21_X1  g376(.A(KEYINPUT32), .B1(new_n797), .B2(new_n798), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n801), .A2(new_n791), .A3(new_n802), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT34), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n790), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n782), .A2(new_n786), .A3(new_n789), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n800), .A2(new_n803), .ZN(new_n808));
  OAI21_X1  g383(.A(KEYINPUT34), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n704), .A2(G24), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n604), .B2(new_n704), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(new_n696), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n739), .A2(G25), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n483), .A2(G119), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n485), .A2(G131), .ZN(new_n815));
  OR2_X1    g390(.A1(G95), .A2(G2105), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n816), .B(G2104), .C1(G107), .C2(new_n471), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n814), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n813), .B1(new_n819), .B2(new_n739), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT35), .B(G1991), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n820), .B(new_n822), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n806), .A2(new_n809), .A3(new_n812), .A4(new_n823), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n824), .A2(KEYINPUT36), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n824), .A2(KEYINPUT36), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n770), .B(new_n773), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(G4), .A2(G16), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(new_n615), .B2(G16), .ZN(new_n829));
  INV_X1    g404(.A(G1348), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT30), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n739), .B1(new_n832), .B2(G28), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n833), .A2(KEYINPUT98), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(G28), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(KEYINPUT98), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n746), .A2(new_n747), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n831), .B(new_n837), .C1(new_n838), .C2(G2090), .ZN(new_n839));
  INV_X1    g414(.A(G11), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n765), .A2(G2078), .B1(KEYINPUT31), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(KEYINPUT31), .B2(new_n840), .ZN(new_n842));
  NOR3_X1   g417(.A1(new_n827), .A2(new_n839), .A3(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(KEYINPUT95), .A2(G2072), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n485), .A2(G139), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n472), .A2(new_n473), .A3(G127), .ZN(new_n846));
  INV_X1    g421(.A(G115), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n846), .B1(new_n847), .B2(new_n463), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(G2105), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT25), .Z(new_n851));
  NAND3_X1  g426(.A1(new_n845), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT94), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n853), .A2(new_n739), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n739), .A2(G33), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n844), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(KEYINPUT95), .A2(G2072), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  OR2_X1    g433(.A1(KEYINPUT24), .A2(G34), .ZN(new_n859));
  NAND2_X1  g434(.A1(KEYINPUT24), .A2(G34), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n859), .A2(new_n739), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(G160), .B2(new_n739), .ZN(new_n862));
  AOI22_X1  g437(.A1(new_n740), .A2(new_n741), .B1(G2084), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n858), .A2(new_n863), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(KEYINPUT96), .Z(new_n865));
  OR2_X1    g440(.A1(new_n862), .A2(G2084), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n638), .A2(new_n739), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NAND4_X1  g443(.A1(new_n843), .A2(new_n865), .A3(new_n866), .A4(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(G311));
  NAND2_X1  g445(.A1(new_n869), .A2(KEYINPUT101), .ZN(new_n871));
  NOR4_X1   g446(.A1(new_n827), .A2(new_n867), .A3(new_n839), .A4(new_n842), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT101), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n872), .A2(new_n873), .A3(new_n865), .A4(new_n866), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n871), .A2(new_n874), .ZN(G150));
  INV_X1    g450(.A(G93), .ZN(new_n876));
  INV_X1    g451(.A(G55), .ZN(new_n877));
  OAI22_X1  g452(.A1(new_n876), .A2(new_n533), .B1(new_n536), .B2(new_n877), .ZN(new_n878));
  AOI22_X1  g453(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n879), .A2(new_n513), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(G860), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n883), .B(KEYINPUT37), .Z(new_n884));
  XNOR2_X1  g459(.A(new_n624), .B(new_n881), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT39), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n615), .A2(G559), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT38), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n886), .B(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n884), .B1(new_n889), .B2(G860), .ZN(G145));
  NAND2_X1  g465(.A1(new_n483), .A2(G130), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n485), .A2(G142), .ZN(new_n892));
  OAI21_X1  g467(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n471), .A2(G118), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n891), .B(new_n892), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(new_n818), .ZN(new_n896));
  XOR2_X1   g471(.A(new_n896), .B(KEYINPUT102), .Z(new_n897));
  INV_X1    g472(.A(new_n641), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n896), .B(KEYINPUT102), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n641), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n738), .B(G164), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(new_n727), .ZN(new_n904));
  INV_X1    g479(.A(new_n852), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n904), .A2(new_n853), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n902), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n638), .B(G160), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(G162), .ZN(new_n911));
  INV_X1    g486(.A(new_n908), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n901), .B(new_n899), .C1(new_n912), .C2(new_n906), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n909), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n911), .B1(new_n909), .B2(new_n913), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(G37), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g494(.A(new_n885), .B(KEYINPUT103), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(new_n628), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n615), .B(G299), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(KEYINPUT41), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n922), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n921), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(KEYINPUT42), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n604), .B(G288), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT104), .ZN(new_n930));
  XNOR2_X1  g505(.A(G166), .B(G305), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n929), .B(KEYINPUT104), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n932), .B1(new_n934), .B2(new_n931), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n921), .A2(new_n924), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT42), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n936), .B(new_n937), .C1(new_n926), .C2(new_n921), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n928), .A2(new_n935), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n935), .B1(new_n928), .B2(new_n938), .ZN(new_n940));
  OAI21_X1  g515(.A(G868), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n882), .A2(new_n625), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(G295));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n942), .ZN(G331));
  XNOR2_X1  g519(.A(G301), .B(G286), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n885), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n885), .A2(new_n945), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT105), .B1(new_n948), .B2(new_n923), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n922), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT105), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n924), .A2(new_n951), .A3(new_n946), .A4(new_n947), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n949), .A2(new_n935), .A3(new_n950), .A4(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(new_n917), .ZN(new_n954));
  INV_X1    g529(.A(new_n935), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n949), .A2(new_n950), .A3(new_n952), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n958));
  INV_X1    g533(.A(new_n954), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n923), .A2(KEYINPUT106), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT41), .ZN(new_n961));
  NOR3_X1   g536(.A1(new_n922), .A2(KEYINPUT106), .A3(new_n961), .ZN(new_n962));
  OR2_X1    g537(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n950), .B1(new_n963), .B2(new_n948), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(new_n955), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n959), .A2(new_n965), .A3(KEYINPUT43), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT44), .B1(new_n958), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT43), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n959), .A2(new_n965), .A3(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n969), .B1(new_n957), .B2(new_n968), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n967), .A2(new_n972), .ZN(G397));
  INV_X1    g548(.A(G1384), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n493), .A2(new_n496), .A3(new_n494), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n471), .B1(new_n498), .B2(new_n499), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT45), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n476), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n468), .A2(new_n469), .ZN(new_n981));
  OAI211_X1 g556(.A(G40), .B(new_n980), .C1(new_n981), .C2(G2105), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n984), .A2(G1996), .ZN(new_n985));
  XOR2_X1   g560(.A(new_n985), .B(KEYINPUT46), .Z(new_n986));
  XNOR2_X1  g561(.A(new_n727), .B(G2067), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n983), .B1(new_n987), .B2(new_n738), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n989), .B(KEYINPUT127), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n990), .B(KEYINPUT47), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n738), .B(G1996), .ZN(new_n992));
  OR2_X1    g567(.A1(new_n992), .A2(new_n987), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n818), .A2(new_n821), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  OAI22_X1  g570(.A1(new_n993), .A2(new_n995), .B1(G2067), .B2(new_n727), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(new_n983), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n604), .A2(new_n696), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n984), .A2(new_n998), .ZN(new_n999));
  XOR2_X1   g574(.A(new_n999), .B(KEYINPUT48), .Z(new_n1000));
  NOR2_X1   g575(.A1(new_n819), .A2(new_n822), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n993), .A2(new_n1001), .A3(new_n994), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1000), .B1(new_n1002), .B2(new_n984), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n991), .A2(new_n997), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(G1384), .B1(new_n497), .B2(new_n501), .ZN(new_n1005));
  INV_X1    g580(.A(G40), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n470), .A2(new_n1006), .A3(new_n476), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1008), .A2(G2067), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n982), .B1(KEYINPUT50), .B2(new_n977), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT108), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT50), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1005), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1012), .B(new_n974), .C1(new_n975), .C2(new_n976), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT108), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1010), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1009), .B1(new_n1016), .B2(new_n830), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AOI211_X1 g594(.A(KEYINPUT118), .B(new_n1009), .C1(new_n1016), .C2(new_n830), .ZN(new_n1020));
  OAI21_X1  g595(.A(KEYINPUT60), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1021), .A2(KEYINPUT122), .A3(new_n627), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n1014), .B(new_n1011), .ZN(new_n1023));
  AOI21_X1  g598(.A(G1348), .B1(new_n1023), .B2(new_n1010), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT118), .B1(new_n1024), .B2(new_n1009), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  OR2_X1    g602(.A1(new_n1027), .A2(KEYINPUT60), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n627), .A2(KEYINPUT122), .ZN(new_n1029));
  OR2_X1    g604(.A1(new_n627), .A2(KEYINPUT122), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1027), .A2(KEYINPUT60), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1022), .A2(new_n1028), .A3(new_n1031), .ZN(new_n1032));
  OAI211_X1 g607(.A(KEYINPUT45), .B(new_n974), .C1(new_n975), .C2(new_n976), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n979), .A2(new_n1007), .A3(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g609(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n1035));
  XNOR2_X1  g610(.A(new_n1035), .B(G2072), .ZN(new_n1036));
  OR2_X1    g611(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n977), .A2(KEYINPUT50), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1038), .A2(new_n1007), .A3(new_n1014), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1039), .A2(new_n1040), .A3(new_n762), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1040), .B1(new_n1039), .B2(new_n762), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1037), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n573), .A2(KEYINPUT77), .A3(new_n574), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT77), .B1(new_n573), .B2(new_n574), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n1046), .A2(G651), .B1(G91), .B2(new_n534), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT57), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1047), .A2(KEYINPUT116), .A3(new_n1048), .A4(new_n572), .ZN(new_n1049));
  OR2_X1    g624(.A1(new_n1048), .A2(KEYINPUT116), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1048), .A2(KEYINPUT116), .ZN(new_n1051));
  NAND3_X1  g626(.A1(G299), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1043), .A2(new_n1053), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1055), .B(new_n1037), .C1(new_n1042), .C2(new_n1041), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n1057), .A2(KEYINPUT61), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1054), .A2(new_n1056), .A3(KEYINPUT61), .ZN(new_n1059));
  XOR2_X1   g634(.A(KEYINPUT58), .B(G1341), .Z(new_n1060));
  NAND2_X1  g635(.A1(new_n1008), .A2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g636(.A(KEYINPUT120), .B(G1996), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1061), .B1(new_n1034), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT121), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1063), .A2(new_n564), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT59), .ZN(new_n1066));
  OR2_X1    g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1068));
  AND3_X1   g643(.A1(new_n1059), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1032), .A2(new_n1058), .A3(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1043), .A2(new_n1053), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1025), .A2(new_n1026), .A3(new_n615), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1071), .B1(new_n1072), .B2(new_n1054), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n1073), .B(KEYINPUT119), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1070), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(G2084), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1010), .A2(new_n1013), .A3(new_n1076), .A4(new_n1015), .ZN(new_n1077));
  INV_X1    g652(.A(G1966), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1034), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(G8), .ZN(new_n1081));
  NAND2_X1  g656(.A1(G286), .A2(G8), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT123), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT51), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1081), .A2(new_n1082), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1080), .A2(G8), .A3(G286), .ZN(new_n1088));
  OAI211_X1 g663(.A(G8), .B(new_n1085), .C1(new_n1080), .C2(G286), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(KEYINPUT124), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT124), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1087), .A2(new_n1092), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT54), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT107), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1034), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(G2078), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n979), .A2(KEYINPUT107), .A3(new_n1007), .A4(new_n1033), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n1101));
  INV_X1    g676(.A(G1961), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1100), .A2(new_n1101), .B1(new_n1102), .B2(new_n1016), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n470), .A2(new_n1006), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1101), .A2(G2078), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n979), .A2(new_n1033), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n474), .A2(new_n475), .ZN(new_n1107));
  OAI21_X1  g682(.A(G2105), .B1(new_n1107), .B2(KEYINPUT125), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1108), .B1(KEYINPUT125), .B2(new_n1107), .ZN(new_n1109));
  OR2_X1    g684(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1110));
  AND3_X1   g685(.A1(new_n1103), .A2(G301), .A3(new_n1110), .ZN(new_n1111));
  OR2_X1    g686(.A1(new_n1106), .A2(new_n476), .ZN(new_n1112));
  AOI21_X1  g687(.A(G301), .B1(new_n1103), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1095), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1094), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(G1971), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1039), .A2(G2090), .ZN(new_n1117));
  OAI21_X1  g692(.A(G8), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT55), .ZN(new_n1119));
  INV_X1    g694(.A(G8), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1119), .B1(G166), .B2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT109), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT109), .ZN(new_n1124));
  NAND4_X1  g699(.A1(G303), .A2(new_n1124), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1123), .A2(KEYINPUT110), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT110), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1118), .A2(new_n1121), .A3(new_n1126), .A4(new_n1129), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n511), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1131));
  INV_X1    g706(.A(G48), .ZN(new_n1132));
  OAI22_X1  g707(.A1(new_n1131), .A2(new_n513), .B1(new_n1132), .B2(new_n536), .ZN(new_n1133));
  XOR2_X1   g708(.A(KEYINPUT113), .B(G86), .Z(new_n1134));
  NOR2_X1   g709(.A1(new_n533), .A2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(G1981), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1136), .B1(G305), .B2(G1981), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT49), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1120), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1136), .B(KEYINPUT49), .C1(G305), .C2(G1981), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT52), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n586), .A2(new_n585), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1144), .A2(G1976), .A3(new_n584), .A4(new_n587), .ZN(new_n1145));
  INV_X1    g720(.A(G1976), .ZN(new_n1146));
  NAND2_X1  g721(.A1(G288), .A2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1140), .A2(new_n1143), .A3(new_n1145), .A4(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1143), .B1(new_n1140), .B2(new_n1145), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1148), .B1(new_n1149), .B2(KEYINPUT112), .ZN(new_n1150));
  AND3_X1   g725(.A1(new_n1008), .A2(G8), .A3(new_n1145), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT112), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1151), .A2(new_n1152), .A3(new_n1143), .A4(new_n1147), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1142), .A2(new_n1150), .A3(new_n1153), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n1130), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1103), .A2(G301), .A3(new_n1112), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1016), .A2(new_n1102), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1157), .A2(new_n1158), .A3(new_n1110), .ZN(new_n1159));
  OAI211_X1 g734(.A(new_n1156), .B(KEYINPUT54), .C1(new_n1159), .C2(G301), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1129), .A2(new_n1121), .A3(new_n1126), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT111), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1129), .A2(KEYINPUT111), .A3(new_n1121), .A4(new_n1126), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1016), .A2(G2090), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1116), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1166), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1163), .A2(G8), .A3(new_n1164), .A4(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1155), .A2(new_n1160), .A3(new_n1168), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1115), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1075), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT114), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1081), .A2(G286), .ZN(new_n1173));
  OAI211_X1 g748(.A(new_n1154), .B(new_n1173), .C1(new_n1167), .C2(new_n1161), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(KEYINPUT63), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1142), .A2(new_n1146), .ZN(new_n1176));
  OAI22_X1  g751(.A1(new_n1176), .A2(G288), .B1(G1981), .B2(G305), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1177), .A2(new_n1140), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1175), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1154), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n1081), .A2(KEYINPUT63), .A3(G286), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1130), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1180), .B1(new_n1168), .B2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1172), .B1(new_n1179), .B2(new_n1183), .ZN(new_n1184));
  AOI22_X1  g759(.A1(new_n1174), .A2(KEYINPUT63), .B1(new_n1140), .B2(new_n1177), .ZN(new_n1185));
  AND2_X1   g760(.A1(new_n1164), .A2(G8), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1166), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1187));
  AOI22_X1  g762(.A1(new_n1186), .A2(new_n1187), .B1(new_n1130), .B2(new_n1181), .ZN(new_n1188));
  OAI211_X1 g763(.A(new_n1185), .B(KEYINPUT114), .C1(new_n1188), .C2(new_n1180), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1184), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n1191));
  AND3_X1   g766(.A1(new_n1171), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1191), .B1(new_n1171), .B2(new_n1190), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1155), .A2(new_n1168), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1113), .B1(new_n1094), .B2(KEYINPUT62), .ZN(new_n1195));
  AOI211_X1 g770(.A(new_n1194), .B(new_n1195), .C1(KEYINPUT62), .C2(new_n1094), .ZN(new_n1196));
  NOR3_X1   g771(.A1(new_n1192), .A2(new_n1193), .A3(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(new_n1002), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1198), .B1(G1986), .B2(G290), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n984), .B1(new_n1199), .B2(new_n998), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1004), .B1(new_n1197), .B2(new_n1200), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g776(.A(new_n677), .B1(new_n657), .B2(new_n658), .ZN(new_n1203));
  AOI21_X1  g777(.A(new_n1203), .B1(new_n916), .B2(new_n917), .ZN(new_n1204));
  INV_X1    g778(.A(G229), .ZN(new_n1205));
  NAND4_X1  g779(.A1(new_n1204), .A2(new_n970), .A3(G319), .A4(new_n1205), .ZN(G225));
  INV_X1    g780(.A(G225), .ZN(G308));
endmodule


