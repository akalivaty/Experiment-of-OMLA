

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735;

  NAND2_X1 U364 ( .A1(n372), .A2(n349), .ZN(n612) );
  XNOR2_X1 U365 ( .A(n500), .B(n499), .ZN(n720) );
  INV_X1 U366 ( .A(G953), .ZN(n722) );
  XNOR2_X2 U367 ( .A(n535), .B(n534), .ZN(n689) );
  XNOR2_X2 U368 ( .A(n507), .B(n365), .ZN(n672) );
  XNOR2_X1 U369 ( .A(n401), .B(G116), .ZN(n366) );
  INV_X1 U370 ( .A(n601), .ZN(n438) );
  NAND2_X2 U371 ( .A1(n541), .A2(n529), .ZN(n431) );
  INV_X2 U372 ( .A(G113), .ZN(n401) );
  OR2_X2 U373 ( .A1(n360), .A2(n494), .ZN(n426) );
  XNOR2_X1 U374 ( .A(n572), .B(n443), .ZN(n579) );
  INV_X1 U375 ( .A(n569), .ZN(n369) );
  OR2_X1 U376 ( .A1(n721), .A2(KEYINPUT2), .ZN(n693) );
  AND2_X1 U377 ( .A1(n357), .A2(n355), .ZN(n721) );
  XNOR2_X1 U378 ( .A(n376), .B(n375), .ZN(n735) );
  AND2_X1 U379 ( .A1(n382), .A2(n387), .ZN(n386) );
  NOR2_X1 U380 ( .A1(n583), .A2(n584), .ZN(n589) );
  NOR2_X1 U381 ( .A1(n579), .A2(n459), .ZN(n427) );
  NOR2_X1 U382 ( .A1(n531), .A2(n601), .ZN(n529) );
  XNOR2_X1 U383 ( .A(n368), .B(n367), .ZN(n674) );
  NAND2_X1 U384 ( .A1(n380), .A2(n656), .ZN(n572) );
  XNOR2_X1 U385 ( .A(n626), .B(n625), .ZN(n627) );
  XNOR2_X1 U386 ( .A(n366), .B(n444), .ZN(n361) );
  XNOR2_X1 U387 ( .A(KEYINPUT32), .B(KEYINPUT78), .ZN(n430) );
  XOR2_X1 U388 ( .A(G143), .B(G128), .Z(n464) );
  XNOR2_X2 U389 ( .A(n473), .B(G140), .ZN(n474) );
  NOR2_X1 U390 ( .A1(n668), .A2(n533), .ZN(n368) );
  NAND2_X1 U391 ( .A1(n558), .A2(n559), .ZN(n561) );
  NOR2_X2 U392 ( .A1(n374), .A2(n543), .ZN(n631) );
  INV_X1 U393 ( .A(G472), .ZN(n365) );
  NOR2_X1 U394 ( .A1(G902), .A2(n626), .ZN(n507) );
  INV_X1 U395 ( .A(G146), .ZN(n524) );
  INV_X1 U396 ( .A(G137), .ZN(n497) );
  XNOR2_X1 U397 ( .A(n402), .B(n432), .ZN(n527) );
  XNOR2_X1 U398 ( .A(n433), .B(G107), .ZN(n432) );
  XNOR2_X1 U399 ( .A(n434), .B(n445), .ZN(n402) );
  INV_X1 U400 ( .A(KEYINPUT72), .ZN(n433) );
  XNOR2_X1 U401 ( .A(n488), .B(n487), .ZN(n550) );
  XNOR2_X1 U402 ( .A(KEYINPUT13), .B(G475), .ZN(n487) );
  NAND2_X1 U403 ( .A1(n704), .A2(n350), .ZN(n397) );
  INV_X1 U404 ( .A(KEYINPUT47), .ZN(n415) );
  NOR2_X1 U405 ( .A1(n735), .A2(n733), .ZN(n595) );
  XNOR2_X1 U406 ( .A(n362), .B(KEYINPUT73), .ZN(n503) );
  NAND2_X1 U407 ( .A1(n722), .A2(n363), .ZN(n362) );
  INV_X1 U408 ( .A(G237), .ZN(n363) );
  XNOR2_X1 U409 ( .A(n540), .B(n539), .ZN(n559) );
  INV_X1 U410 ( .A(KEYINPUT44), .ZN(n539) );
  INV_X1 U411 ( .A(G134), .ZN(n465) );
  XNOR2_X1 U412 ( .A(n408), .B(n407), .ZN(n514) );
  INV_X1 U413 ( .A(KEYINPUT8), .ZN(n407) );
  NAND2_X1 U414 ( .A1(n722), .A2(G234), .ZN(n408) );
  XNOR2_X1 U415 ( .A(n498), .B(n346), .ZN(n371) );
  XNOR2_X1 U416 ( .A(KEYINPUT18), .B(KEYINPUT85), .ZN(n446) );
  XOR2_X1 U417 ( .A(KEYINPUT86), .B(KEYINPUT17), .Z(n447) );
  OR2_X1 U418 ( .A1(G237), .A2(G902), .ZN(n454) );
  XNOR2_X1 U419 ( .A(n522), .B(n521), .ZN(n668) );
  XNOR2_X1 U420 ( .A(G101), .B(KEYINPUT92), .ZN(n501) );
  XOR2_X1 U421 ( .A(KEYINPUT5), .B(KEYINPUT93), .Z(n502) );
  XNOR2_X1 U422 ( .A(KEYINPUT3), .B(G119), .ZN(n444) );
  XOR2_X1 U423 ( .A(KEYINPUT68), .B(KEYINPUT10), .Z(n475) );
  XNOR2_X1 U424 ( .A(G128), .B(G137), .ZN(n509) );
  XOR2_X1 U425 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n510) );
  XNOR2_X1 U426 ( .A(n720), .B(n441), .ZN(n700) );
  XNOR2_X1 U427 ( .A(n527), .B(n442), .ZN(n441) );
  XNOR2_X1 U428 ( .A(n526), .B(n525), .ZN(n442) );
  XNOR2_X1 U429 ( .A(n590), .B(KEYINPUT39), .ZN(n600) );
  XNOR2_X1 U430 ( .A(n422), .B(n421), .ZN(n420) );
  INV_X1 U431 ( .A(KEYINPUT28), .ZN(n421) );
  INV_X1 U432 ( .A(KEYINPUT107), .ZN(n388) );
  OR2_X1 U433 ( .A1(n343), .A2(n388), .ZN(n387) );
  XNOR2_X1 U434 ( .A(n427), .B(n460), .ZN(n360) );
  XOR2_X1 U435 ( .A(KEYINPUT102), .B(n552), .Z(n633) );
  INV_X1 U436 ( .A(KEYINPUT1), .ZN(n439) );
  NOR2_X1 U437 ( .A1(n396), .A2(n395), .ZN(n394) );
  NOR2_X1 U438 ( .A1(n429), .A2(G478), .ZN(n396) );
  XNOR2_X1 U439 ( .A(n354), .B(n470), .ZN(n702) );
  XNOR2_X1 U440 ( .A(n378), .B(n472), .ZN(n354) );
  XNOR2_X1 U441 ( .A(n351), .B(KEYINPUT101), .ZN(n469) );
  XNOR2_X1 U442 ( .A(n614), .B(KEYINPUT54), .ZN(n615) );
  NAND2_X1 U443 ( .A1(n643), .A2(n415), .ZN(n412) );
  NAND2_X1 U444 ( .A1(n591), .A2(n493), .ZN(n494) );
  NAND2_X1 U445 ( .A1(n597), .A2(n596), .ZN(n358) );
  XNOR2_X1 U446 ( .A(G104), .B(G101), .ZN(n434) );
  INV_X1 U447 ( .A(G110), .ZN(n445) );
  XNOR2_X1 U448 ( .A(G104), .B(G131), .ZN(n482) );
  XOR2_X1 U449 ( .A(KEYINPUT97), .B(KEYINPUT95), .Z(n479) );
  XNOR2_X1 U450 ( .A(G122), .B(G113), .ZN(n476) );
  XNOR2_X1 U451 ( .A(n524), .B(n523), .ZN(n525) );
  INV_X1 U452 ( .A(G140), .ZN(n523) );
  XNOR2_X1 U453 ( .A(KEYINPUT6), .B(KEYINPUT106), .ZN(n508) );
  INV_X1 U454 ( .A(KEYINPUT38), .ZN(n379) );
  INV_X1 U455 ( .A(n577), .ZN(n423) );
  NOR2_X1 U456 ( .A1(n356), .A2(n654), .ZN(n355) );
  XNOR2_X1 U457 ( .A(n358), .B(n598), .ZN(n357) );
  INV_X1 U458 ( .A(n653), .ZN(n356) );
  XNOR2_X1 U459 ( .A(KEYINPUT45), .B(KEYINPUT64), .ZN(n560) );
  NAND2_X1 U460 ( .A1(n468), .A2(n467), .ZN(n351) );
  XNOR2_X1 U461 ( .A(n471), .B(n341), .ZN(n378) );
  XNOR2_X1 U462 ( .A(n448), .B(n371), .ZN(n449) );
  NAND2_X1 U463 ( .A1(G234), .A2(G237), .ZN(n456) );
  XNOR2_X1 U464 ( .A(n603), .B(n364), .ZN(n571) );
  INV_X1 U465 ( .A(KEYINPUT111), .ZN(n364) );
  XNOR2_X1 U466 ( .A(n404), .B(KEYINPUT74), .ZN(n583) );
  XNOR2_X1 U467 ( .A(n353), .B(n352), .ZN(n551) );
  INV_X1 U468 ( .A(G478), .ZN(n352) );
  OR2_X1 U469 ( .A1(n702), .A2(G902), .ZN(n353) );
  INV_X1 U470 ( .A(KEYINPUT67), .ZN(n367) );
  INV_X1 U471 ( .A(G469), .ZN(n440) );
  NOR2_X1 U472 ( .A1(n700), .A2(G902), .ZN(n528) );
  BUF_X1 U473 ( .A(n668), .Z(n374) );
  NOR2_X2 U474 ( .A1(n530), .A2(n369), .ZN(n541) );
  XNOR2_X1 U475 ( .A(n720), .B(n424), .ZN(n626) );
  XNOR2_X1 U476 ( .A(n398), .B(n527), .ZN(n709) );
  XNOR2_X1 U477 ( .A(n361), .B(n399), .ZN(n398) );
  XNOR2_X1 U478 ( .A(n400), .B(KEYINPUT16), .ZN(n399) );
  INV_X1 U479 ( .A(G122), .ZN(n400) );
  XNOR2_X1 U480 ( .A(G110), .B(G119), .ZN(n512) );
  XNOR2_X1 U481 ( .A(n619), .B(n618), .ZN(n620) );
  INV_X1 U482 ( .A(KEYINPUT40), .ZN(n375) );
  XNOR2_X1 U483 ( .A(n389), .B(KEYINPUT35), .ZN(n730) );
  OR2_X1 U484 ( .A1(n593), .A2(n579), .ZN(n643) );
  NAND2_X1 U485 ( .A1(n385), .A2(n384), .ZN(n383) );
  AND2_X1 U486 ( .A1(n343), .A2(n388), .ZN(n384) );
  OR2_X1 U487 ( .A1(n550), .A2(n551), .ZN(n648) );
  NAND2_X1 U488 ( .A1(n393), .A2(n391), .ZN(n428) );
  NAND2_X1 U489 ( .A1(n392), .A2(n702), .ZN(n391) );
  AND2_X1 U490 ( .A1(n397), .A2(n394), .ZN(n393) );
  XNOR2_X1 U491 ( .A(n406), .B(n405), .ZN(n701) );
  XNOR2_X1 U492 ( .A(n700), .B(n699), .ZN(n405) );
  NAND2_X1 U493 ( .A1(n704), .A2(G469), .ZN(n406) );
  INV_X1 U494 ( .A(KEYINPUT56), .ZN(n435) );
  XOR2_X1 U495 ( .A(n463), .B(n462), .Z(n341) );
  XOR2_X1 U496 ( .A(n586), .B(KEYINPUT76), .Z(n342) );
  XNOR2_X1 U497 ( .A(n672), .B(n508), .ZN(n569) );
  AND2_X1 U498 ( .A1(n601), .A2(n532), .ZN(n343) );
  AND2_X1 U499 ( .A1(n692), .A2(n691), .ZN(n344) );
  AND2_X1 U500 ( .A1(n411), .A2(n412), .ZN(n345) );
  AND2_X1 U501 ( .A1(G224), .A2(n722), .ZN(n346) );
  AND2_X1 U502 ( .A1(n576), .A2(n403), .ZN(n347) );
  XNOR2_X1 U503 ( .A(KEYINPUT34), .B(KEYINPUT77), .ZN(n348) );
  XOR2_X1 U504 ( .A(n608), .B(KEYINPUT66), .Z(n349) );
  AND2_X1 U505 ( .A1(n429), .A2(G478), .ZN(n350) );
  XOR2_X1 U506 ( .A(G902), .B(KEYINPUT15), .Z(n489) );
  XOR2_X1 U507 ( .A(KEYINPUT84), .B(n617), .Z(n703) );
  INV_X1 U508 ( .A(n703), .ZN(n395) );
  XNOR2_X1 U509 ( .A(n351), .B(n497), .ZN(n500) );
  NAND2_X1 U510 ( .A1(n359), .A2(n652), .ZN(n410) );
  NAND2_X1 U511 ( .A1(n345), .A2(n409), .ZN(n359) );
  OR2_X1 U512 ( .A1(n360), .A2(n689), .ZN(n536) );
  OR2_X1 U513 ( .A1(n360), .A2(n581), .ZN(n548) );
  NOR2_X1 U514 ( .A1(n546), .A2(n360), .ZN(n547) );
  XNOR2_X1 U515 ( .A(n361), .B(n524), .ZN(n425) );
  NOR2_X1 U516 ( .A1(n410), .A2(n587), .ZN(n377) );
  NAND2_X1 U517 ( .A1(n570), .A2(n633), .ZN(n603) );
  XNOR2_X1 U518 ( .A(n506), .B(n425), .ZN(n424) );
  NAND2_X1 U519 ( .A1(n386), .A2(n383), .ZN(n732) );
  NAND2_X1 U520 ( .A1(n695), .A2(n418), .ZN(n417) );
  NAND2_X1 U521 ( .A1(n370), .A2(n369), .ZN(n535) );
  INV_X1 U522 ( .A(n544), .ZN(n370) );
  XNOR2_X1 U523 ( .A(n416), .B(KEYINPUT122), .ZN(n697) );
  NOR2_X1 U524 ( .A1(n732), .A2(n730), .ZN(n538) );
  XNOR2_X1 U525 ( .A(n516), .B(n517), .ZN(n706) );
  NAND2_X1 U526 ( .A1(n373), .A2(n489), .ZN(n372) );
  INV_X1 U527 ( .A(n610), .ZN(n373) );
  NAND2_X1 U528 ( .A1(n600), .A2(n633), .ZN(n376) );
  NAND2_X1 U529 ( .A1(n381), .A2(n721), .ZN(n610) );
  XNOR2_X1 U530 ( .A(n428), .B(KEYINPUT123), .ZN(G63) );
  XNOR2_X1 U531 ( .A(n377), .B(n588), .ZN(n597) );
  XNOR2_X1 U532 ( .A(n380), .B(n379), .ZN(n657) );
  NAND2_X1 U533 ( .A1(n589), .A2(n380), .ZN(n585) );
  NOR2_X1 U534 ( .A1(n606), .A2(n380), .ZN(n654) );
  XNOR2_X2 U535 ( .A(n453), .B(n452), .ZN(n380) );
  OR2_X1 U536 ( .A1(n381), .A2(KEYINPUT2), .ZN(n694) );
  NAND2_X1 U537 ( .A1(n381), .A2(n722), .ZN(n714) );
  XNOR2_X2 U538 ( .A(n561), .B(n560), .ZN(n381) );
  NAND2_X1 U539 ( .A1(n530), .A2(KEYINPUT107), .ZN(n382) );
  XNOR2_X1 U540 ( .A(n536), .B(n348), .ZN(n390) );
  INV_X1 U541 ( .A(n530), .ZN(n385) );
  NAND2_X1 U542 ( .A1(n390), .A2(n342), .ZN(n389) );
  INV_X1 U543 ( .A(n704), .ZN(n392) );
  AND2_X4 U544 ( .A1(n612), .A2(n611), .ZN(n704) );
  NAND2_X1 U545 ( .A1(n674), .A2(n576), .ZN(n581) );
  NAND2_X1 U546 ( .A1(n674), .A2(n347), .ZN(n404) );
  INV_X1 U547 ( .A(n582), .ZN(n403) );
  NAND2_X1 U548 ( .A1(n661), .A2(n415), .ZN(n411) );
  XOR2_X2 U549 ( .A(G125), .B(G146), .Z(n473) );
  XNOR2_X2 U550 ( .A(n475), .B(n474), .ZN(n719) );
  NAND2_X1 U551 ( .A1(n413), .A2(n414), .ZN(n409) );
  INV_X1 U552 ( .A(n643), .ZN(n413) );
  NOR2_X1 U553 ( .A1(n661), .A2(n415), .ZN(n414) );
  NAND2_X1 U554 ( .A1(n417), .A2(n344), .ZN(n416) );
  NOR2_X1 U555 ( .A1(n696), .A2(n419), .ZN(n418) );
  INV_X1 U556 ( .A(n694), .ZN(n419) );
  INV_X1 U557 ( .A(n672), .ZN(n578) );
  NAND2_X1 U558 ( .A1(n420), .A2(n576), .ZN(n593) );
  NAND2_X1 U559 ( .A1(n672), .A2(n423), .ZN(n422) );
  XNOR2_X2 U560 ( .A(n426), .B(n496), .ZN(n530) );
  INV_X1 U561 ( .A(n702), .ZN(n429) );
  NAND2_X1 U562 ( .A1(n538), .A2(n731), .ZN(n540) );
  XNOR2_X2 U563 ( .A(n431), .B(n430), .ZN(n731) );
  XNOR2_X1 U564 ( .A(n436), .B(n435), .ZN(G51) );
  NAND2_X1 U565 ( .A1(n437), .A2(n703), .ZN(n436) );
  XNOR2_X1 U566 ( .A(n616), .B(n615), .ZN(n437) );
  NAND2_X1 U567 ( .A1(n674), .A2(n438), .ZN(n544) );
  XNOR2_X2 U568 ( .A(n576), .B(n439), .ZN(n601) );
  XNOR2_X2 U569 ( .A(n528), .B(n440), .ZN(n576) );
  XNOR2_X1 U570 ( .A(KEYINPUT75), .B(KEYINPUT19), .ZN(n443) );
  XNOR2_X1 U571 ( .A(KEYINPUT81), .B(KEYINPUT48), .ZN(n598) );
  INV_X1 U572 ( .A(n533), .ZN(n493) );
  XNOR2_X1 U573 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U574 ( .A(n483), .B(n482), .ZN(n484) );
  INV_X1 U575 ( .A(KEYINPUT22), .ZN(n495) );
  XNOR2_X1 U576 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U577 ( .A(n495), .B(KEYINPUT71), .ZN(n496) );
  INV_X1 U578 ( .A(n374), .ZN(n531) );
  XNOR2_X1 U579 ( .A(KEYINPUT36), .B(KEYINPUT112), .ZN(n573) );
  XNOR2_X1 U580 ( .A(n621), .B(n620), .ZN(n622) );
  INV_X1 U581 ( .A(KEYINPUT60), .ZN(n623) );
  INV_X1 U582 ( .A(KEYINPUT0), .ZN(n460) );
  XNOR2_X1 U583 ( .A(n709), .B(n473), .ZN(n451) );
  XOR2_X1 U584 ( .A(KEYINPUT4), .B(KEYINPUT65), .Z(n498) );
  XNOR2_X1 U585 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U586 ( .A(n464), .B(n449), .Z(n450) );
  XNOR2_X1 U587 ( .A(n451), .B(n450), .ZN(n613) );
  NOR2_X1 U588 ( .A1(n613), .A2(n489), .ZN(n453) );
  NAND2_X1 U589 ( .A1(G210), .A2(n454), .ZN(n452) );
  NAND2_X1 U590 ( .A1(G214), .A2(n454), .ZN(n656) );
  XOR2_X1 U591 ( .A(KEYINPUT87), .B(G898), .Z(n711) );
  NOR2_X1 U592 ( .A1(n711), .A2(n722), .ZN(n708) );
  NAND2_X1 U593 ( .A1(n708), .A2(G902), .ZN(n455) );
  NAND2_X1 U594 ( .A1(G952), .A2(n722), .ZN(n562) );
  NAND2_X1 U595 ( .A1(n455), .A2(n562), .ZN(n458) );
  XOR2_X1 U596 ( .A(KEYINPUT14), .B(n456), .Z(n687) );
  INV_X1 U597 ( .A(n687), .ZN(n457) );
  NAND2_X1 U598 ( .A1(n458), .A2(n457), .ZN(n459) );
  XNOR2_X1 U599 ( .A(G107), .B(G122), .ZN(n461) );
  XNOR2_X1 U600 ( .A(n461), .B(KEYINPUT100), .ZN(n472) );
  XOR2_X1 U601 ( .A(KEYINPUT7), .B(KEYINPUT99), .Z(n463) );
  XNOR2_X1 U602 ( .A(G116), .B(KEYINPUT98), .ZN(n462) );
  NAND2_X1 U603 ( .A1(n465), .A2(n464), .ZN(n468) );
  XNOR2_X1 U604 ( .A(G143), .B(G128), .ZN(n466) );
  NAND2_X1 U605 ( .A1(G134), .A2(n466), .ZN(n467) );
  XNOR2_X1 U606 ( .A(n469), .B(KEYINPUT9), .ZN(n470) );
  NAND2_X1 U607 ( .A1(G217), .A2(n514), .ZN(n471) );
  INV_X1 U608 ( .A(n551), .ZN(n537) );
  XOR2_X1 U609 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n477) );
  XNOR2_X1 U610 ( .A(n477), .B(n476), .ZN(n481) );
  XNOR2_X1 U611 ( .A(G143), .B(KEYINPUT96), .ZN(n478) );
  XNOR2_X1 U612 ( .A(n479), .B(n478), .ZN(n480) );
  XOR2_X1 U613 ( .A(n481), .B(n480), .Z(n485) );
  NAND2_X1 U614 ( .A1(n503), .A2(G214), .ZN(n483) );
  XNOR2_X1 U615 ( .A(n719), .B(n486), .ZN(n619) );
  NOR2_X1 U616 ( .A1(G902), .A2(n619), .ZN(n488) );
  NOR2_X1 U617 ( .A1(n537), .A2(n550), .ZN(n591) );
  XOR2_X1 U618 ( .A(KEYINPUT89), .B(KEYINPUT21), .Z(n492) );
  INV_X1 U619 ( .A(n489), .ZN(n607) );
  NAND2_X1 U620 ( .A1(n607), .A2(G234), .ZN(n490) );
  XNOR2_X1 U621 ( .A(n490), .B(KEYINPUT20), .ZN(n518) );
  NAND2_X1 U622 ( .A1(n518), .A2(G221), .ZN(n491) );
  XNOR2_X1 U623 ( .A(n492), .B(n491), .ZN(n667) );
  XNOR2_X1 U624 ( .A(KEYINPUT90), .B(n667), .ZN(n533) );
  XNOR2_X1 U625 ( .A(n498), .B(G131), .ZN(n499) );
  XOR2_X1 U626 ( .A(n502), .B(n501), .Z(n505) );
  NAND2_X1 U627 ( .A1(n503), .A2(G210), .ZN(n504) );
  XNOR2_X1 U628 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U629 ( .A(n511), .B(KEYINPUT70), .Z(n513) );
  XNOR2_X1 U630 ( .A(n513), .B(n512), .ZN(n517) );
  NAND2_X1 U631 ( .A1(n514), .A2(G221), .ZN(n515) );
  XNOR2_X1 U632 ( .A(n515), .B(n719), .ZN(n516) );
  NOR2_X1 U633 ( .A1(G902), .A2(n706), .ZN(n522) );
  XOR2_X1 U634 ( .A(KEYINPUT88), .B(KEYINPUT25), .Z(n520) );
  NAND2_X1 U635 ( .A1(G217), .A2(n518), .ZN(n519) );
  XNOR2_X1 U636 ( .A(n520), .B(n519), .ZN(n521) );
  NAND2_X1 U637 ( .A1(G227), .A2(n722), .ZN(n526) );
  NOR2_X1 U638 ( .A1(n672), .A2(n531), .ZN(n532) );
  XOR2_X1 U639 ( .A(KEYINPUT108), .B(KEYINPUT33), .Z(n534) );
  NAND2_X1 U640 ( .A1(n537), .A2(n550), .ZN(n586) );
  XNOR2_X1 U641 ( .A(n541), .B(KEYINPUT82), .ZN(n542) );
  NAND2_X1 U642 ( .A1(n542), .A2(n601), .ZN(n543) );
  NOR2_X1 U643 ( .A1(n578), .A2(n544), .ZN(n545) );
  XNOR2_X1 U644 ( .A(KEYINPUT94), .B(n545), .ZN(n678) );
  INV_X1 U645 ( .A(n678), .ZN(n546) );
  XNOR2_X1 U646 ( .A(KEYINPUT31), .B(n547), .ZN(n647) );
  XNOR2_X1 U647 ( .A(n548), .B(KEYINPUT91), .ZN(n549) );
  NAND2_X1 U648 ( .A1(n549), .A2(n578), .ZN(n637) );
  NAND2_X1 U649 ( .A1(n647), .A2(n637), .ZN(n555) );
  XNOR2_X1 U650 ( .A(KEYINPUT103), .B(n648), .ZN(n599) );
  NAND2_X1 U651 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X1 U652 ( .A1(n599), .A2(n633), .ZN(n553) );
  XNOR2_X1 U653 ( .A(KEYINPUT104), .B(n553), .ZN(n661) );
  INV_X1 U654 ( .A(n661), .ZN(n554) );
  NAND2_X1 U655 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U656 ( .A(n556), .B(KEYINPUT105), .ZN(n557) );
  NOR2_X1 U657 ( .A1(n631), .A2(n557), .ZN(n558) );
  NOR2_X1 U658 ( .A1(n562), .A2(n687), .ZN(n567) );
  NAND2_X1 U659 ( .A1(G953), .A2(G902), .ZN(n563) );
  NOR2_X1 U660 ( .A1(n687), .A2(n563), .ZN(n564) );
  XNOR2_X1 U661 ( .A(n564), .B(KEYINPUT109), .ZN(n565) );
  NOR2_X1 U662 ( .A1(G900), .A2(n565), .ZN(n566) );
  NOR2_X1 U663 ( .A1(n567), .A2(n566), .ZN(n582) );
  NOR2_X1 U664 ( .A1(n582), .A2(n667), .ZN(n568) );
  NAND2_X1 U665 ( .A1(n568), .A2(n374), .ZN(n577) );
  NOR2_X1 U666 ( .A1(n569), .A2(n577), .ZN(n570) );
  NOR2_X1 U667 ( .A1(n572), .A2(n571), .ZN(n574) );
  XNOR2_X1 U668 ( .A(n574), .B(n573), .ZN(n575) );
  NAND2_X1 U669 ( .A1(n575), .A2(n438), .ZN(n652) );
  NAND2_X1 U670 ( .A1(n672), .A2(n656), .ZN(n580) );
  XNOR2_X1 U671 ( .A(KEYINPUT30), .B(n580), .ZN(n584) );
  NOR2_X1 U672 ( .A1(n586), .A2(n585), .ZN(n642) );
  XOR2_X1 U673 ( .A(KEYINPUT79), .B(n642), .Z(n587) );
  INV_X1 U674 ( .A(KEYINPUT69), .ZN(n588) );
  NAND2_X1 U675 ( .A1(n589), .A2(n657), .ZN(n590) );
  NAND2_X1 U676 ( .A1(n657), .A2(n656), .ZN(n662) );
  INV_X1 U677 ( .A(n591), .ZN(n658) );
  NOR2_X1 U678 ( .A1(n662), .A2(n658), .ZN(n592) );
  XNOR2_X1 U679 ( .A(KEYINPUT41), .B(n592), .ZN(n690) );
  NOR2_X1 U680 ( .A1(n593), .A2(n690), .ZN(n594) );
  XNOR2_X1 U681 ( .A(n594), .B(KEYINPUT42), .ZN(n733) );
  XNOR2_X1 U682 ( .A(KEYINPUT46), .B(n595), .ZN(n596) );
  NAND2_X1 U683 ( .A1(n600), .A2(n599), .ZN(n653) );
  NAND2_X1 U684 ( .A1(n601), .A2(n656), .ZN(n602) );
  NOR2_X1 U685 ( .A1(n603), .A2(n602), .ZN(n605) );
  XNOR2_X1 U686 ( .A(KEYINPUT43), .B(KEYINPUT110), .ZN(n604) );
  XNOR2_X1 U687 ( .A(n605), .B(n604), .ZN(n606) );
  INV_X1 U688 ( .A(KEYINPUT2), .ZN(n609) );
  NOR2_X1 U689 ( .A1(n607), .A2(n609), .ZN(n608) );
  NOR2_X2 U690 ( .A1(n610), .A2(n609), .ZN(n696) );
  INV_X1 U691 ( .A(n696), .ZN(n611) );
  NAND2_X1 U692 ( .A1(n704), .A2(G210), .ZN(n616) );
  XNOR2_X1 U693 ( .A(n613), .B(KEYINPUT55), .ZN(n614) );
  NOR2_X1 U694 ( .A1(G952), .A2(n722), .ZN(n617) );
  NAND2_X1 U695 ( .A1(n704), .A2(G475), .ZN(n621) );
  XOR2_X1 U696 ( .A(KEYINPUT59), .B(KEYINPUT83), .Z(n618) );
  NAND2_X1 U697 ( .A1(n622), .A2(n703), .ZN(n624) );
  XNOR2_X1 U698 ( .A(n624), .B(n623), .ZN(G60) );
  NAND2_X1 U699 ( .A1(n704), .A2(G472), .ZN(n628) );
  INV_X1 U700 ( .A(KEYINPUT62), .ZN(n625) );
  XNOR2_X1 U701 ( .A(n628), .B(n627), .ZN(n629) );
  NAND2_X1 U702 ( .A1(n629), .A2(n703), .ZN(n630) );
  XNOR2_X1 U703 ( .A(n630), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U704 ( .A(G101), .B(n631), .ZN(n632) );
  XNOR2_X1 U705 ( .A(n632), .B(KEYINPUT113), .ZN(G3) );
  INV_X1 U706 ( .A(n633), .ZN(n645) );
  NOR2_X1 U707 ( .A1(n645), .A2(n637), .ZN(n634) );
  XOR2_X1 U708 ( .A(G104), .B(n634), .Z(G6) );
  XOR2_X1 U709 ( .A(KEYINPUT114), .B(KEYINPUT26), .Z(n636) );
  XNOR2_X1 U710 ( .A(G107), .B(KEYINPUT27), .ZN(n635) );
  XNOR2_X1 U711 ( .A(n636), .B(n635), .ZN(n639) );
  NOR2_X1 U712 ( .A1(n648), .A2(n637), .ZN(n638) );
  XOR2_X1 U713 ( .A(n639), .B(n638), .Z(G9) );
  NOR2_X1 U714 ( .A1(n648), .A2(n643), .ZN(n641) );
  XNOR2_X1 U715 ( .A(G128), .B(KEYINPUT29), .ZN(n640) );
  XNOR2_X1 U716 ( .A(n641), .B(n640), .ZN(G30) );
  XOR2_X1 U717 ( .A(G143), .B(n642), .Z(G45) );
  NOR2_X1 U718 ( .A1(n645), .A2(n643), .ZN(n644) );
  XOR2_X1 U719 ( .A(G146), .B(n644), .Z(G48) );
  NOR2_X1 U720 ( .A1(n645), .A2(n647), .ZN(n646) );
  XOR2_X1 U721 ( .A(G113), .B(n646), .Z(G15) );
  NOR2_X1 U722 ( .A1(n648), .A2(n647), .ZN(n650) );
  XNOR2_X1 U723 ( .A(G116), .B(KEYINPUT115), .ZN(n649) );
  XNOR2_X1 U724 ( .A(n650), .B(n649), .ZN(G18) );
  XOR2_X1 U725 ( .A(G125), .B(KEYINPUT37), .Z(n651) );
  XNOR2_X1 U726 ( .A(n652), .B(n651), .ZN(G27) );
  XNOR2_X1 U727 ( .A(G134), .B(n653), .ZN(G36) );
  XOR2_X1 U728 ( .A(G140), .B(n654), .Z(n655) );
  XNOR2_X1 U729 ( .A(KEYINPUT116), .B(n655), .ZN(G42) );
  NOR2_X1 U730 ( .A1(n657), .A2(n656), .ZN(n659) );
  NOR2_X1 U731 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U732 ( .A(KEYINPUT119), .B(n660), .Z(n664) );
  NOR2_X1 U733 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U734 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U735 ( .A(n665), .B(KEYINPUT120), .ZN(n666) );
  NOR2_X1 U736 ( .A1(n689), .A2(n666), .ZN(n683) );
  NAND2_X1 U737 ( .A1(n374), .A2(n667), .ZN(n669) );
  XNOR2_X1 U738 ( .A(n669), .B(KEYINPUT49), .ZN(n670) );
  XOR2_X1 U739 ( .A(KEYINPUT117), .B(n670), .Z(n671) );
  NOR2_X1 U740 ( .A1(n672), .A2(n671), .ZN(n673) );
  XOR2_X1 U741 ( .A(KEYINPUT118), .B(n673), .Z(n677) );
  NOR2_X1 U742 ( .A1(n674), .A2(n438), .ZN(n675) );
  XNOR2_X1 U743 ( .A(KEYINPUT50), .B(n675), .ZN(n676) );
  NOR2_X1 U744 ( .A1(n677), .A2(n676), .ZN(n679) );
  NOR2_X1 U745 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U746 ( .A(KEYINPUT51), .B(n680), .Z(n681) );
  NOR2_X1 U747 ( .A1(n690), .A2(n681), .ZN(n682) );
  NOR2_X1 U748 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U749 ( .A(KEYINPUT121), .B(n684), .Z(n685) );
  XNOR2_X1 U750 ( .A(n685), .B(KEYINPUT52), .ZN(n686) );
  NOR2_X1 U751 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U752 ( .A1(G952), .A2(n688), .ZN(n692) );
  OR2_X1 U753 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U754 ( .A(n693), .B(KEYINPUT80), .ZN(n695) );
  NOR2_X1 U755 ( .A1(G953), .A2(n697), .ZN(n698) );
  XNOR2_X1 U756 ( .A(KEYINPUT53), .B(n698), .ZN(G75) );
  XOR2_X1 U757 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n699) );
  NOR2_X1 U758 ( .A1(n395), .A2(n701), .ZN(G54) );
  NAND2_X1 U759 ( .A1(G217), .A2(n704), .ZN(n705) );
  XNOR2_X1 U760 ( .A(n706), .B(n705), .ZN(n707) );
  NOR2_X1 U761 ( .A1(n395), .A2(n707), .ZN(G66) );
  NOR2_X1 U762 ( .A1(n709), .A2(n708), .ZN(n718) );
  NAND2_X1 U763 ( .A1(G953), .A2(G224), .ZN(n710) );
  XNOR2_X1 U764 ( .A(KEYINPUT61), .B(n710), .ZN(n712) );
  NAND2_X1 U765 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U766 ( .A(n713), .B(KEYINPUT124), .ZN(n715) );
  NAND2_X1 U767 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U768 ( .A(n716), .B(KEYINPUT125), .Z(n717) );
  XNOR2_X1 U769 ( .A(n718), .B(n717), .ZN(G69) );
  XNOR2_X1 U770 ( .A(n720), .B(n719), .ZN(n725) );
  XOR2_X1 U771 ( .A(n725), .B(n721), .Z(n723) );
  NAND2_X1 U772 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U773 ( .A(n724), .B(KEYINPUT126), .ZN(n729) );
  XNOR2_X1 U774 ( .A(G227), .B(n725), .ZN(n726) );
  NAND2_X1 U775 ( .A1(n726), .A2(G900), .ZN(n727) );
  NAND2_X1 U776 ( .A1(G953), .A2(n727), .ZN(n728) );
  NAND2_X1 U777 ( .A1(n729), .A2(n728), .ZN(G72) );
  XOR2_X1 U778 ( .A(n730), .B(G122), .Z(G24) );
  XNOR2_X1 U779 ( .A(n731), .B(G119), .ZN(G21) );
  XOR2_X1 U780 ( .A(G110), .B(n732), .Z(G12) );
  XNOR2_X1 U781 ( .A(G137), .B(KEYINPUT127), .ZN(n734) );
  XNOR2_X1 U782 ( .A(n734), .B(n733), .ZN(G39) );
  XOR2_X1 U783 ( .A(n735), .B(G131), .Z(G33) );
endmodule

