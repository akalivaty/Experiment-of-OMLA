//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 1 1 1 1 0 1 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 1 0 0 1 0 0 0 1 0 1 0 1 1 1 1 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n559, new_n561, new_n562, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n571, new_n572, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1167,
    new_n1168;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XOR2_X1   g016(.A(KEYINPUT65), .B(G108), .Z(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT66), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g020(.A(KEYINPUT67), .B(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT68), .Z(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n464), .A2(G137), .A3(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT70), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  AND3_X1   g045(.A1(new_n466), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n467), .B1(new_n466), .B2(new_n470), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n464), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n474), .B1(new_n475), .B2(new_n465), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  AND2_X1   g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(G125), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n477), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n482), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n476), .A2(new_n483), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n473), .A2(new_n484), .ZN(G160));
  NOR2_X1   g060(.A1(new_n480), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n480), .A2(new_n465), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n487), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  AND2_X1   g068(.A1(KEYINPUT71), .A2(G138), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n465), .B(new_n494), .C1(new_n478), .C2(new_n479), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n464), .A2(new_n497), .A3(new_n465), .A4(new_n494), .ZN(new_n498));
  AND2_X1   g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n469), .A2(G102), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n464), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(new_n465), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n499), .A2(new_n502), .ZN(G164));
  NAND2_X1  g078(.A1(G75), .A2(G543), .ZN(new_n504));
  AND3_X1   g079(.A1(KEYINPUT72), .A2(KEYINPUT5), .A3(G543), .ZN(new_n505));
  AOI21_X1  g080(.A(KEYINPUT5), .B1(KEYINPUT72), .B2(G543), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G62), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n504), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT6), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n509), .A2(G651), .B1(G50), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  OAI21_X1  g093(.A(KEYINPUT73), .B1(new_n507), .B2(new_n514), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT72), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT5), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(KEYINPUT72), .A2(KEYINPUT5), .A3(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT73), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT6), .B(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n519), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n517), .B1(new_n518), .B2(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  NAND3_X1  g105(.A1(new_n519), .A2(G89), .A3(new_n527), .ZN(new_n531));
  OAI211_X1 g106(.A(G63), .B(G651), .C1(new_n505), .C2(new_n506), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT74), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT74), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n524), .A2(new_n534), .A3(G63), .A4(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n516), .A2(G51), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AND3_X1   g115(.A1(new_n531), .A2(new_n536), .A3(new_n540), .ZN(G168));
  AND4_X1   g116(.A1(G52), .A2(new_n511), .A3(new_n513), .A4(G543), .ZN(new_n542));
  OAI21_X1  g117(.A(G64), .B1(new_n505), .B2(new_n506), .ZN(new_n543));
  NAND2_X1  g118(.A1(G77), .A2(G543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n542), .B1(new_n545), .B2(G651), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n519), .A2(G90), .A3(new_n527), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(G171));
  AND2_X1   g124(.A1(new_n519), .A2(new_n527), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G81), .ZN(new_n551));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G56), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n507), .B2(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n554), .A2(G651), .B1(G43), .B2(new_n516), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  AND3_X1   g133(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G36), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n562), .ZN(G188));
  AND3_X1   g138(.A1(new_n526), .A2(G53), .A3(G543), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n564), .B(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n519), .A2(G91), .A3(new_n527), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n524), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n568), .A2(new_n510), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(G299));
  AND3_X1   g145(.A1(new_n546), .A2(new_n547), .A3(KEYINPUT75), .ZN(new_n571));
  AOI21_X1  g146(.A(KEYINPUT75), .B1(new_n546), .B2(new_n547), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n571), .A2(new_n572), .ZN(G301));
  NAND3_X1  g148(.A1(new_n531), .A2(new_n536), .A3(new_n540), .ZN(G286));
  NAND3_X1  g149(.A1(new_n519), .A2(G87), .A3(new_n527), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT76), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n519), .A2(KEYINPUT76), .A3(new_n527), .A4(G87), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n577), .A2(new_n578), .B1(G49), .B2(new_n516), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT78), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT77), .ZN(new_n582));
  AND3_X1   g157(.A1(new_n579), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n580), .B1(new_n579), .B2(new_n582), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G288));
  NAND2_X1  g161(.A1(new_n550), .A2(G86), .ZN(new_n587));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n588), .B(KEYINPUT79), .ZN(new_n589));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n590), .B2(new_n507), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n591), .A2(G651), .B1(G48), .B2(new_n516), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n587), .A2(new_n592), .ZN(G305));
  NAND2_X1  g168(.A1(new_n516), .A2(G47), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G85), .ZN(new_n596));
  OAI221_X1 g171(.A(new_n594), .B1(new_n510), .B2(new_n595), .C1(new_n528), .C2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  XNOR2_X1  g174(.A(KEYINPUT80), .B(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n507), .B2(new_n600), .ZN(new_n601));
  AND2_X1   g176(.A1(new_n601), .A2(G651), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n550), .A2(KEYINPUT10), .A3(G92), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n528), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n602), .B1(new_n603), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n516), .A2(G54), .ZN(new_n608));
  AND2_X1   g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n598), .B1(new_n609), .B2(G868), .ZN(G284));
  OAI21_X1  g185(.A(new_n598), .B1(new_n609), .B2(G868), .ZN(G321));
  NAND2_X1  g186(.A1(G286), .A2(G868), .ZN(new_n612));
  INV_X1    g187(.A(G299), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(G868), .ZN(G297));
  OAI21_X1  g189(.A(new_n612), .B1(new_n613), .B2(G868), .ZN(G280));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n609), .B1(new_n616), .B2(G860), .ZN(G148));
  NAND2_X1  g192(.A1(new_n607), .A2(new_n608), .ZN(new_n618));
  OR3_X1    g193(.A1(new_n618), .A2(KEYINPUT81), .A3(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(KEYINPUT81), .B1(new_n618), .B2(G559), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G868), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n557), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n486), .A2(G135), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n488), .A2(G123), .ZN(new_n626));
  NOR2_X1   g201(.A1(G99), .A2(G2105), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(new_n465), .B2(G111), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n625), .B(new_n626), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT84), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2096), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n464), .A2(new_n469), .ZN(new_n632));
  XOR2_X1   g207(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT13), .ZN(new_n635));
  XOR2_X1   g210(.A(KEYINPUT83), .B(G2100), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n631), .A2(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2435), .ZN(new_n640));
  XOR2_X1   g215(.A(G2427), .B(G2438), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(KEYINPUT14), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT85), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n643), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n649), .B(new_n650), .Z(new_n651));
  AND2_X1   g226(.A1(new_n651), .A2(G14), .ZN(G401));
  XOR2_X1   g227(.A(G2067), .B(G2678), .Z(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AND2_X1   g231(.A1(new_n656), .A2(KEYINPUT17), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n654), .A2(new_n655), .ZN(new_n658));
  AOI21_X1  g233(.A(KEYINPUT18), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2072), .B(G2078), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT86), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(KEYINPUT18), .B2(new_n656), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n659), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2096), .B(G2100), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(G227));
  XNOR2_X1  g240(.A(G1971), .B(G1976), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  XOR2_X1   g242(.A(G1956), .B(G2474), .Z(new_n668));
  XOR2_X1   g243(.A(G1961), .B(G1966), .Z(new_n669));
  OR2_X1    g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT87), .Z(new_n672));
  NAND2_X1  g247(.A1(new_n668), .A2(new_n669), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT88), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(new_n667), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n667), .A2(new_n673), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT20), .Z(new_n678));
  NAND3_X1  g253(.A1(new_n672), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1991), .B(G1996), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1981), .B(G1986), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n683), .A2(new_n685), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(G229));
  MUX2_X1   g263(.A(G24), .B(G290), .S(G16), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G1986), .ZN(new_n690));
  INV_X1    g265(.A(G16), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n691), .A2(G23), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n577), .A2(new_n578), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n516), .A2(G49), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n693), .A2(new_n694), .A3(new_n582), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n692), .B1(new_n695), .B2(G16), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT33), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(G1976), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n696), .B(KEYINPUT33), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G1976), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n691), .A2(G6), .ZN(new_n703));
  INV_X1    g278(.A(G305), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n703), .B1(new_n704), .B2(new_n691), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT32), .B(G1981), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n691), .A2(G22), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G166), .B2(new_n691), .ZN(new_n709));
  INV_X1    g284(.A(G1971), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND4_X1  g286(.A1(new_n700), .A2(new_n702), .A3(new_n707), .A4(new_n711), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT91), .B(KEYINPUT34), .Z(new_n713));
  AOI21_X1  g288(.A(new_n690), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(G25), .A2(G29), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n486), .A2(G131), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n488), .A2(G119), .ZN(new_n717));
  NOR2_X1   g292(.A1(G95), .A2(G2105), .ZN(new_n718));
  OAI21_X1  g293(.A(G2104), .B1(new_n465), .B2(G107), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n716), .B(new_n717), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT89), .Z(new_n721));
  AOI21_X1  g296(.A(new_n715), .B1(new_n721), .B2(G29), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT35), .B(G1991), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT90), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n722), .B(new_n724), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n714), .B(new_n725), .C1(new_n713), .C2(new_n712), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT36), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n727), .A2(KEYINPUT92), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(G171), .A2(G16), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G5), .B2(G16), .ZN(new_n731));
  INV_X1    g306(.A(G1961), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT102), .Z(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT31), .B(G11), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n691), .A2(G21), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G168), .B2(new_n691), .ZN(new_n737));
  INV_X1    g312(.A(G1966), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n630), .A2(G29), .ZN(new_n740));
  INV_X1    g315(.A(G28), .ZN(new_n741));
  AOI21_X1  g316(.A(G29), .B1(new_n741), .B2(KEYINPUT30), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(KEYINPUT30), .B2(new_n741), .ZN(new_n743));
  AND3_X1   g318(.A1(new_n739), .A2(new_n740), .A3(new_n743), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n734), .A2(new_n735), .A3(new_n744), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n745), .A2(KEYINPUT103), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n691), .A2(G19), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n557), .B2(new_n691), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT94), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G1341), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n745), .A2(KEYINPUT103), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n691), .A2(G4), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n609), .B2(new_n691), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT93), .B(G1348), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n753), .B(new_n755), .ZN(new_n756));
  NAND4_X1  g331(.A1(new_n746), .A2(new_n750), .A3(new_n751), .A4(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(G29), .A2(G33), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n464), .A2(G127), .ZN(new_n759));
  AND2_X1   g334(.A1(G115), .A2(G2104), .ZN(new_n760));
  OAI21_X1  g335(.A(G2105), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT98), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n761), .A2(new_n762), .B1(G139), .B2(new_n486), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n469), .A2(G103), .ZN(new_n764));
  XOR2_X1   g339(.A(KEYINPUT97), .B(KEYINPUT25), .Z(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  OAI211_X1 g341(.A(KEYINPUT98), .B(G2105), .C1(new_n759), .C2(new_n760), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n763), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT99), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n763), .A2(KEYINPUT99), .A3(new_n766), .A4(new_n767), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(KEYINPUT100), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT100), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n770), .A2(new_n774), .A3(new_n771), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n758), .B1(new_n776), .B2(G29), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G2072), .ZN(new_n778));
  INV_X1    g353(.A(G29), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(G35), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G162), .B2(new_n779), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT106), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT29), .B(G2090), .Z(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(G160), .A2(new_n779), .ZN(new_n785));
  AND2_X1   g360(.A1(KEYINPUT24), .A2(G34), .ZN(new_n786));
  NOR2_X1   g361(.A1(KEYINPUT24), .A2(G34), .ZN(new_n787));
  NOR3_X1   g362(.A1(new_n786), .A2(new_n787), .A3(G29), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(G2084), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n779), .A2(G27), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G164), .B2(new_n779), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT105), .B(G2078), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NOR3_X1   g370(.A1(new_n784), .A2(new_n791), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n789), .A2(new_n790), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n731), .A2(new_n732), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n486), .A2(G141), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n488), .A2(G129), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n469), .A2(G105), .ZN(new_n801));
  NAND3_X1  g376(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT26), .Z(new_n803));
  NAND4_X1  g378(.A1(new_n799), .A2(new_n800), .A3(new_n801), .A4(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n805), .A2(G29), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G29), .B2(G32), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT27), .B(G1996), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n797), .B(new_n798), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT104), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n807), .A2(new_n808), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT101), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT107), .B(KEYINPUT23), .Z(new_n815));
  NAND2_X1  g390(.A1(new_n691), .A2(G20), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(new_n613), .B2(new_n691), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(G1956), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n814), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n796), .A2(new_n811), .A3(new_n812), .A4(new_n820), .ZN(new_n821));
  NOR3_X1   g396(.A1(new_n757), .A2(new_n778), .A3(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT28), .ZN(new_n823));
  AND2_X1   g398(.A1(new_n779), .A2(G26), .ZN(new_n824));
  OAI21_X1  g399(.A(G2104), .B1(new_n465), .B2(G116), .ZN(new_n825));
  INV_X1    g400(.A(G104), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n825), .B1(new_n826), .B2(new_n465), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT95), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n486), .A2(G140), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n488), .A2(G128), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  AOI211_X1 g406(.A(new_n823), .B(new_n824), .C1(new_n831), .C2(G29), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(new_n823), .B2(new_n824), .ZN(new_n833));
  XNOR2_X1  g408(.A(KEYINPUT96), .B(G2067), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n727), .A2(KEYINPUT92), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n726), .A2(new_n728), .A3(new_n836), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n729), .A2(new_n822), .A3(new_n835), .A4(new_n837), .ZN(G150));
  INV_X1    g413(.A(G150), .ZN(G311));
  NAND3_X1  g414(.A1(new_n519), .A2(G93), .A3(new_n527), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT109), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n516), .A2(G55), .ZN(new_n842));
  AND3_X1   g417(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n841), .B1(new_n840), .B2(new_n842), .ZN(new_n844));
  AOI22_X1  g419(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n845));
  OAI22_X1  g420(.A1(new_n843), .A2(new_n844), .B1(new_n510), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(G860), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT37), .Z(new_n848));
  NOR2_X1   g423(.A1(new_n618), .A2(new_n616), .ZN(new_n849));
  XOR2_X1   g424(.A(KEYINPUT108), .B(KEYINPUT38), .Z(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT39), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n849), .B(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n846), .B(new_n557), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n848), .B1(new_n854), .B2(G860), .ZN(G145));
  NAND2_X1  g430(.A1(new_n486), .A2(G142), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n488), .A2(G130), .ZN(new_n857));
  NOR2_X1   g432(.A1(G106), .A2(G2105), .ZN(new_n858));
  OAI21_X1  g433(.A(G2104), .B1(new_n465), .B2(G118), .ZN(new_n859));
  OAI211_X1 g434(.A(new_n856), .B(new_n857), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n720), .B(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n634), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n831), .A2(G164), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n831), .A2(G164), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n804), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n865), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n867), .A2(new_n805), .A3(new_n863), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n776), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n866), .A2(new_n868), .A3(new_n772), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n862), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(KEYINPUT110), .ZN(new_n873));
  XNOR2_X1  g448(.A(G160), .B(new_n492), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n630), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n870), .A2(new_n862), .A3(new_n871), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT110), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n873), .B(new_n875), .C1(new_n878), .C2(new_n872), .ZN(new_n879));
  INV_X1    g454(.A(G37), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n872), .A2(new_n875), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(new_n876), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT40), .ZN(G395));
  OR2_X1    g459(.A1(new_n846), .A2(G868), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n621), .A2(new_n853), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n618), .A2(new_n613), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n607), .A2(G299), .A3(new_n608), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n846), .B(new_n556), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n619), .A2(new_n620), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n887), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n893), .A2(KEYINPUT111), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(KEYINPUT111), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  XOR2_X1   g471(.A(G305), .B(KEYINPUT112), .Z(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(G166), .B(G290), .ZN(new_n899));
  INV_X1    g474(.A(new_n695), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n899), .A2(new_n900), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n898), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n903), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n905), .A2(new_n897), .A3(new_n901), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT42), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n907), .A2(new_n908), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT113), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n911), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT113), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n913), .A2(new_n909), .A3(new_n914), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n887), .A2(new_n892), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n888), .A2(KEYINPUT41), .A3(new_n889), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT41), .B1(new_n888), .B2(new_n889), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OR2_X1    g494(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n896), .A2(new_n912), .A3(new_n915), .A4(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n920), .A2(new_n895), .A3(new_n894), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n922), .A2(new_n914), .A3(new_n913), .A4(new_n909), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n886), .B1(new_n924), .B2(G868), .ZN(G295));
  AOI21_X1  g500(.A(new_n886), .B1(new_n924), .B2(G868), .ZN(G331));
  OAI21_X1  g501(.A(G168), .B1(new_n571), .B2(new_n572), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT114), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n928), .B1(G168), .B2(new_n548), .ZN(new_n929));
  NAND3_X1  g504(.A1(G171), .A2(G286), .A3(KEYINPUT114), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n927), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT115), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n927), .A2(new_n929), .A3(KEYINPUT115), .A4(new_n930), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n891), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n934), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n853), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n919), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n937), .A2(KEYINPUT116), .A3(new_n935), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT116), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n891), .A2(new_n933), .A3(new_n940), .A4(new_n934), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n938), .B1(new_n942), .B2(new_n890), .ZN(new_n943));
  AOI21_X1  g518(.A(G37), .B1(new_n943), .B2(new_n907), .ZN(new_n944));
  INV_X1    g519(.A(new_n907), .ZN(new_n945));
  INV_X1    g520(.A(new_n890), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n946), .B1(new_n939), .B2(new_n941), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n945), .B1(new_n947), .B2(new_n938), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT43), .B1(new_n944), .B2(new_n948), .ZN(new_n949));
  NOR3_X1   g524(.A1(new_n947), .A2(new_n945), .A3(new_n938), .ZN(new_n950));
  OR2_X1    g525(.A1(new_n917), .A2(new_n918), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n939), .A2(new_n951), .A3(new_n941), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n937), .A2(new_n890), .A3(new_n935), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n907), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT43), .ZN(new_n955));
  NOR4_X1   g530(.A1(new_n950), .A2(new_n954), .A3(new_n955), .A4(G37), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT44), .B1(new_n949), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n955), .B1(new_n944), .B2(new_n948), .ZN(new_n959));
  NOR4_X1   g534(.A1(new_n950), .A2(new_n954), .A3(KEYINPUT43), .A4(G37), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n957), .A2(new_n961), .ZN(G397));
  OR2_X1    g537(.A1(new_n831), .A2(G2067), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n831), .A2(G2067), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G1996), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n804), .B(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n723), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n721), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n963), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G1384), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n972), .B1(new_n499), .B2(new_n502), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT45), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n473), .A2(new_n484), .A3(G40), .ZN(new_n976));
  OR3_X1    g551(.A1(new_n975), .A2(new_n976), .A3(KEYINPUT117), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT117), .B1(new_n975), .B2(new_n976), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n971), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(G290), .A2(G1986), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  XOR2_X1   g557(.A(new_n982), .B(KEYINPUT48), .Z(new_n983));
  INV_X1    g558(.A(new_n968), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n720), .B(new_n969), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n983), .B1(new_n979), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n979), .A2(new_n966), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT46), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n989), .A2(KEYINPUT127), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n988), .B(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(KEYINPUT127), .ZN(new_n992));
  INV_X1    g567(.A(new_n965), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n979), .B1(new_n804), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n991), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  OR2_X1    g570(.A1(new_n995), .A2(KEYINPUT47), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(KEYINPUT47), .ZN(new_n997));
  AOI211_X1 g572(.A(new_n980), .B(new_n987), .C1(new_n996), .C2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G1981), .ZN(new_n999));
  XNOR2_X1  g574(.A(G305), .B(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT49), .ZN(new_n1001));
  OR2_X1    g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1003));
  NAND2_X1  g578(.A1(G114), .A2(G2104), .ZN(new_n1004));
  INV_X1    g579(.A(G126), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1004), .B1(new_n480), .B2(new_n1005), .ZN(new_n1006));
  AOI22_X1  g581(.A1(new_n1006), .A2(G2105), .B1(G102), .B2(new_n469), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n496), .A2(new_n498), .ZN(new_n1008));
  AOI21_X1  g583(.A(G1384), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1009), .A2(G40), .A3(new_n473), .A4(new_n484), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1010), .A2(KEYINPUT119), .A3(G8), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(G8), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT119), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  AOI22_X1  g589(.A1(new_n1002), .A2(new_n1003), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n900), .A2(G1976), .ZN(new_n1016));
  NAND2_X1  g591(.A1(KEYINPUT120), .A2(KEYINPUT52), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n1010), .A2(KEYINPUT119), .A3(G8), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT119), .B1(new_n1010), .B2(G8), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1016), .B(new_n1017), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT121), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n695), .A2(KEYINPUT78), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n579), .A2(new_n580), .A3(new_n582), .ZN(new_n1024));
  AOI21_X1  g599(.A(G1976), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1022), .B1(new_n1025), .B2(KEYINPUT52), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n699), .B1(new_n583), .B2(new_n584), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1027), .A2(KEYINPUT121), .A3(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1021), .A2(new_n1026), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1014), .A2(new_n1011), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n1016), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1032), .B1(KEYINPUT120), .B2(new_n1028), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1015), .B1(new_n1030), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(G303), .A2(G8), .ZN(new_n1035));
  XNOR2_X1  g610(.A(new_n1035), .B(KEYINPUT55), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n473), .A2(G40), .A3(new_n484), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n973), .A2(KEYINPUT50), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT50), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1009), .A2(new_n1039), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1037), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(G2090), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1009), .A2(KEYINPUT45), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1037), .A2(new_n975), .A3(new_n1043), .ZN(new_n1044));
  AOI22_X1  g619(.A1(new_n1041), .A2(new_n1042), .B1(new_n1044), .B2(new_n710), .ZN(new_n1045));
  INV_X1    g620(.A(G8), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1036), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT118), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1037), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1048), .B1(new_n1049), .B2(G2090), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1009), .B(KEYINPUT50), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1051), .A2(KEYINPUT118), .A3(new_n1042), .A4(new_n1037), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1044), .A2(new_n710), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1050), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(G8), .ZN(new_n1055));
  OR2_X1    g630(.A1(new_n1055), .A2(new_n1036), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1034), .A2(new_n1047), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n1058));
  INV_X1    g633(.A(G2078), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1037), .A2(new_n975), .A3(new_n1059), .A4(new_n1043), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g637(.A(new_n1009), .B(new_n974), .ZN(new_n1063));
  OAI211_X1 g638(.A(KEYINPUT53), .B(new_n1059), .C1(new_n475), .C2(new_n465), .ZN(new_n1064));
  NOR3_X1   g639(.A1(new_n1064), .A2(new_n471), .A3(new_n472), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1063), .A2(G40), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1049), .A2(new_n732), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1062), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1058), .B1(new_n1068), .B2(G171), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1063), .A2(KEYINPUT53), .A3(new_n1059), .A4(new_n1037), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1070), .A2(new_n1062), .A3(G301), .A4(new_n1067), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n1069), .A2(KEYINPUT126), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT126), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g649(.A(KEYINPUT124), .B(G1996), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1037), .A2(new_n975), .A3(new_n1043), .A4(new_n1075), .ZN(new_n1076));
  XOR2_X1   g651(.A(KEYINPUT58), .B(G1341), .Z(new_n1077));
  NAND2_X1  g652(.A1(new_n1010), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n556), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n1080));
  XNOR2_X1  g655(.A(new_n1079), .B(new_n1080), .ZN(new_n1081));
  OR2_X1    g656(.A1(KEYINPUT123), .A2(KEYINPUT57), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n566), .A2(new_n567), .A3(new_n569), .A4(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(KEYINPUT123), .A2(KEYINPUT57), .ZN(new_n1084));
  XNOR2_X1  g659(.A(new_n1083), .B(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(G1956), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1049), .A2(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g662(.A(KEYINPUT56), .B(G2072), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1037), .A2(new_n975), .A3(new_n1043), .A4(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT125), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(KEYINPUT61), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1085), .A2(new_n1087), .A3(new_n1089), .A4(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1049), .A2(new_n755), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1010), .A2(G2067), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT60), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1093), .A2(new_n1095), .A3(new_n1096), .A4(new_n609), .ZN(new_n1097));
  AND2_X1   g672(.A1(new_n1092), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n754), .B1(new_n1051), .B2(new_n1037), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n618), .B1(new_n1099), .B2(new_n1094), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1093), .A2(new_n1095), .A3(new_n609), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1100), .A2(KEYINPUT60), .A3(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1085), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1103), .A2(new_n1090), .A3(KEYINPUT61), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1081), .A2(new_n1098), .A3(new_n1102), .A4(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1085), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1103), .A2(new_n609), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1106), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1105), .A2(new_n1109), .ZN(new_n1110));
  AOI22_X1  g685(.A1(new_n1041), .A2(new_n790), .B1(new_n1044), .B2(new_n738), .ZN(new_n1111));
  NAND2_X1  g686(.A1(G286), .A2(G8), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT51), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1114), .B(new_n1112), .C1(new_n1111), .C2(new_n1046), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1044), .A2(new_n738), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1037), .A2(new_n1038), .A3(new_n790), .A4(new_n1040), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  OAI211_X1 g693(.A(KEYINPUT51), .B(G8), .C1(new_n1118), .C2(G286), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1113), .B1(new_n1115), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1070), .A2(new_n1062), .A3(new_n1067), .ZN(new_n1121));
  INV_X1    g696(.A(G301), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1062), .A2(new_n1066), .A3(new_n1067), .A4(G301), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT54), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1120), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1074), .A2(new_n1110), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1115), .A2(new_n1119), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1113), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT62), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1123), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1120), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1131), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1057), .B1(new_n1127), .B2(new_n1135), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1111), .A2(new_n1046), .A3(G286), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1030), .A2(new_n1033), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1015), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT63), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1140), .B1(new_n1055), .B2(new_n1036), .ZN(new_n1141));
  AND4_X1   g716(.A1(new_n1056), .A2(new_n1138), .A3(new_n1139), .A4(new_n1141), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1034), .A2(new_n1047), .A3(new_n1056), .A4(new_n1137), .ZN(new_n1143));
  AOI22_X1  g718(.A1(new_n1137), .A2(new_n1142), .B1(new_n1143), .B2(new_n1140), .ZN(new_n1144));
  NOR3_X1   g719(.A1(new_n1015), .A2(G1976), .A3(G288), .ZN(new_n1145));
  NOR2_X1   g720(.A1(G305), .A2(G1981), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1146), .B(KEYINPUT122), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1031), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1034), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1148), .B1(new_n1149), .B2(new_n1056), .ZN(new_n1150));
  NOR3_X1   g725(.A1(new_n1136), .A2(new_n1144), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(new_n979), .ZN(new_n1152));
  INV_X1    g727(.A(new_n986), .ZN(new_n1153));
  XOR2_X1   g728(.A(G290), .B(G1986), .Z(new_n1154));
  AOI21_X1  g729(.A(new_n1152), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n998), .B1(new_n1151), .B2(new_n1155), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g731(.A(G319), .B1(new_n686), .B2(new_n687), .ZN(new_n1158));
  AOI21_X1  g732(.A(G227), .B1(new_n651), .B2(G14), .ZN(new_n1159));
  NAND2_X1  g733(.A1(new_n883), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g734(.A1(new_n943), .A2(new_n907), .ZN(new_n1161));
  NAND3_X1  g735(.A1(new_n1161), .A2(new_n880), .A3(new_n948), .ZN(new_n1162));
  NAND2_X1  g736(.A1(new_n1162), .A2(KEYINPUT43), .ZN(new_n1163));
  INV_X1    g737(.A(new_n954), .ZN(new_n1164));
  NAND3_X1  g738(.A1(new_n944), .A2(new_n955), .A3(new_n1164), .ZN(new_n1165));
  AOI211_X1 g739(.A(new_n1158), .B(new_n1160), .C1(new_n1163), .C2(new_n1165), .ZN(G308));
  INV_X1    g740(.A(new_n1160), .ZN(new_n1167));
  INV_X1    g741(.A(new_n1158), .ZN(new_n1168));
  OAI211_X1 g742(.A(new_n1167), .B(new_n1168), .C1(new_n959), .C2(new_n960), .ZN(G225));
endmodule


