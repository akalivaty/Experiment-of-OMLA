//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 0 1 1 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1266, new_n1267,
    new_n1268, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1338, new_n1339, new_n1340;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n215));
  INV_X1    g0015(.A(G232), .ZN(new_n216));
  INV_X1    g0016(.A(G97), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n215), .B1(new_n202), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n211), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  OR2_X1    g0023(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n224));
  OAI21_X1  g0024(.A(G50), .B1(G58), .B2(G68), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT65), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(KEYINPUT64), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g0029(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n230));
  AND2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OR3_X1    g0031(.A1(new_n226), .A2(new_n209), .A3(new_n231), .ZN(new_n232));
  NAND3_X1  g0032(.A1(new_n214), .A2(new_n224), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G50), .B(G58), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT66), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  OAI21_X1  g0050(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  AND2_X1   g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  OAI21_X1  g0053(.A(KEYINPUT67), .B1(new_n253), .B2(new_n227), .ZN(new_n254));
  AND2_X1   g0054(.A1(G1), .A2(G13), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT67), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n252), .B1(new_n254), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G238), .ZN(new_n260));
  NOR3_X1   g0060(.A1(new_n253), .A2(KEYINPUT67), .A3(new_n227), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n256), .B1(new_n255), .B2(new_n257), .ZN(new_n262));
  OAI211_X1 g0062(.A(G274), .B(new_n252), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT3), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n270), .A2(G226), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G97), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n270), .A2(G1698), .ZN(new_n274));
  OAI211_X1 g0074(.A(new_n272), .B(new_n273), .C1(new_n274), .C2(new_n216), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n229), .A2(new_n230), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n257), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  AND3_X1   g0078(.A1(new_n275), .A2(KEYINPUT69), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(KEYINPUT69), .B1(new_n275), .B2(new_n278), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n265), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(KEYINPUT13), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT13), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n283), .B(new_n265), .C1(new_n279), .C2(new_n280), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT14), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(new_n286), .A3(G169), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT70), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n275), .A2(new_n278), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT69), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n275), .A2(KEYINPUT69), .A3(new_n278), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n264), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n288), .B1(new_n293), .B2(new_n283), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n281), .A2(KEYINPUT70), .A3(KEYINPUT13), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n294), .A2(G179), .A3(new_n284), .A4(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n287), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT72), .ZN(new_n298));
  INV_X1    g0098(.A(G169), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n299), .B1(new_n282), .B2(new_n284), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n298), .B1(new_n300), .B2(new_n286), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n285), .A2(G169), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n302), .A2(KEYINPUT72), .A3(KEYINPUT14), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n297), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G13), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n305), .A2(G1), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G20), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G68), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  XOR2_X1   g0110(.A(new_n310), .B(KEYINPUT12), .Z(new_n311));
  NOR2_X1   g0111(.A1(new_n267), .A2(G20), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G77), .ZN(new_n313));
  NOR2_X1   g0113(.A1(G20), .A2(G33), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  OAI221_X1 g0115(.A(new_n313), .B1(new_n209), .B2(G68), .C1(new_n201), .C2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n210), .A2(G33), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n231), .A2(new_n317), .ZN(new_n318));
  AND2_X1   g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n311), .B1(KEYINPUT11), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n320), .B1(KEYINPUT11), .B2(new_n319), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n318), .A2(new_n308), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n208), .A2(G20), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n322), .A2(G68), .A3(new_n323), .ZN(new_n324));
  XOR2_X1   g0124(.A(new_n324), .B(KEYINPUT71), .Z(new_n325));
  NOR2_X1   g0125(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n304), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n294), .A2(G190), .A3(new_n284), .A4(new_n295), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n285), .A2(G200), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n328), .A2(new_n326), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT68), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n274), .B(new_n333), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n334), .A2(G223), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n270), .A2(new_n271), .ZN(new_n336));
  INV_X1    g0136(.A(G222), .ZN(new_n337));
  INV_X1    g0137(.A(G77), .ZN(new_n338));
  OAI22_X1  g0138(.A1(new_n336), .A2(new_n337), .B1(new_n338), .B2(new_n270), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n278), .B1(new_n335), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G274), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n341), .B1(new_n254), .B2(new_n258), .ZN(new_n342));
  AOI22_X1  g0142(.A1(G226), .A2(new_n259), .B1(new_n342), .B2(new_n252), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G190), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n322), .A2(G50), .A3(new_n323), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n276), .B1(G33), .B2(new_n210), .ZN(new_n347));
  XNOR2_X1  g0147(.A(KEYINPUT8), .B(G58), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n349), .A2(new_n312), .B1(G150), .B2(new_n314), .ZN(new_n350));
  OAI21_X1  g0150(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI221_X1 g0152(.A(new_n346), .B1(G50), .B2(new_n307), .C1(new_n347), .C2(new_n352), .ZN(new_n353));
  XNOR2_X1  g0153(.A(new_n353), .B(KEYINPUT9), .ZN(new_n354));
  INV_X1    g0154(.A(G200), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n345), .B(new_n354), .C1(new_n355), .C2(new_n344), .ZN(new_n356));
  XNOR2_X1  g0156(.A(new_n356), .B(KEYINPUT10), .ZN(new_n357));
  INV_X1    g0157(.A(G179), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n344), .A2(new_n358), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n359), .B(new_n353), .C1(G169), .C2(new_n344), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n202), .A2(new_n309), .ZN(new_n363));
  NOR2_X1   g0163(.A1(G58), .A2(G68), .ZN(new_n364));
  OAI21_X1  g0164(.A(G20), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n314), .A2(G159), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  XNOR2_X1  g0168(.A(KEYINPUT73), .B(G33), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n209), .B(new_n268), .C1(new_n369), .C2(new_n266), .ZN(new_n370));
  OAI21_X1  g0170(.A(G68), .B1(new_n370), .B2(KEYINPUT7), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT7), .ZN(new_n372));
  NOR2_X1   g0172(.A1(KEYINPUT3), .A2(G33), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n267), .A2(KEYINPUT73), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT73), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G33), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n373), .B1(new_n377), .B2(KEYINPUT3), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n372), .B1(new_n378), .B2(new_n209), .ZN(new_n379));
  OAI211_X1 g0179(.A(KEYINPUT16), .B(new_n368), .C1(new_n371), .C2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT16), .ZN(new_n381));
  AOI21_X1  g0181(.A(G20), .B1(KEYINPUT3), .B2(G33), .ZN(new_n382));
  OAI211_X1 g0182(.A(KEYINPUT7), .B(new_n382), .C1(new_n377), .C2(KEYINPUT3), .ZN(new_n383));
  AOI21_X1  g0183(.A(KEYINPUT7), .B1(new_n268), .B2(new_n382), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n309), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n381), .B1(new_n386), .B2(new_n367), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n380), .A2(new_n318), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n348), .B1(new_n208), .B2(G20), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n322), .A2(new_n389), .B1(new_n308), .B2(new_n348), .ZN(new_n390));
  MUX2_X1   g0190(.A(G223), .B(G226), .S(G1698), .Z(new_n391));
  AOI21_X1  g0191(.A(new_n266), .B1(new_n374), .B2(new_n376), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n391), .B1(new_n392), .B2(new_n373), .ZN(new_n393));
  NAND2_X1  g0193(.A1(G33), .A2(G87), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n278), .ZN(new_n396));
  OAI211_X1 g0196(.A(G232), .B(new_n251), .C1(new_n261), .C2(new_n262), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n263), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(G190), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n396), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n277), .B1(new_n393), .B2(new_n394), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n263), .A2(new_n397), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n355), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  AND3_X1   g0203(.A1(new_n400), .A2(KEYINPUT74), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(KEYINPUT74), .B1(new_n400), .B2(new_n403), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n388), .B(new_n390), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n406), .B(KEYINPUT17), .ZN(new_n407));
  OAI21_X1  g0207(.A(G169), .B1(new_n401), .B2(new_n402), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n396), .A2(new_n398), .A3(G179), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n388), .A2(new_n390), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n410), .B(KEYINPUT18), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  XOR2_X1   g0213(.A(KEYINPUT15), .B(G87), .Z(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n312), .ZN(new_n415));
  OAI221_X1 g0215(.A(new_n415), .B1(new_n209), .B2(new_n338), .C1(new_n315), .C2(new_n348), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n416), .A2(new_n318), .B1(new_n338), .B2(new_n308), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n322), .A2(G77), .A3(new_n323), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n259), .A2(G244), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n263), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(G107), .ZN(new_n423));
  OAI22_X1  g0223(.A1(new_n336), .A2(new_n216), .B1(new_n423), .B2(new_n270), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n424), .B1(new_n334), .B2(G238), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n422), .B1(new_n425), .B2(new_n277), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n419), .B1(new_n426), .B2(new_n299), .ZN(new_n427));
  OR2_X1    g0227(.A1(new_n426), .A2(G179), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n426), .A2(G200), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n422), .B(G190), .C1(new_n425), .C2(new_n277), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n430), .A2(new_n431), .A3(new_n419), .ZN(new_n432));
  AND2_X1   g0232(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  AND4_X1   g0233(.A1(new_n332), .A2(new_n362), .A3(new_n413), .A4(new_n433), .ZN(new_n434));
  XNOR2_X1  g0234(.A(KEYINPUT5), .B(G41), .ZN(new_n435));
  INV_X1    g0235(.A(G45), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n436), .A2(G1), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n254), .A2(new_n258), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n435), .A2(new_n437), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n438), .A2(G270), .B1(new_n342), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT79), .ZN(new_n441));
  MUX2_X1   g0241(.A(G257), .B(G264), .S(G1698), .Z(new_n442));
  OAI21_X1  g0242(.A(new_n442), .B1(new_n392), .B2(new_n373), .ZN(new_n443));
  INV_X1    g0243(.A(new_n270), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(G303), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n441), .B1(new_n446), .B2(new_n278), .ZN(new_n447));
  AOI211_X1 g0247(.A(KEYINPUT79), .B(new_n277), .C1(new_n443), .C2(new_n445), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n440), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT80), .ZN(new_n450));
  AND2_X1   g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g0251(.A(KEYINPUT80), .B(new_n440), .C1(new_n447), .C2(new_n448), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(G190), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(G20), .B1(G33), .B2(G283), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n267), .A2(G97), .ZN(new_n456));
  INV_X1    g0256(.A(G116), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n455), .A2(new_n456), .B1(G20), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n318), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT20), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n318), .A2(KEYINPUT20), .A3(new_n458), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n461), .A2(new_n462), .B1(new_n457), .B2(new_n308), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n208), .A2(G33), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n231), .A2(new_n307), .A3(new_n317), .A4(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G116), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n449), .A2(new_n450), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n470), .A2(G200), .A3(new_n452), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n454), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT81), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT81), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n454), .A2(new_n474), .A3(new_n469), .A4(new_n471), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n299), .B1(new_n463), .B2(new_n467), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n470), .A2(new_n477), .A3(new_n452), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT21), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n449), .A2(new_n358), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n468), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n470), .A2(new_n477), .A3(KEYINPUT21), .A4(new_n452), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n268), .B1(new_n369), .B2(new_n266), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n484), .A2(KEYINPUT22), .A3(new_n209), .A4(G87), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n369), .A2(new_n457), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n209), .A2(G107), .ZN(new_n487));
  OR2_X1    g0287(.A1(new_n487), .A2(KEYINPUT23), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(KEYINPUT23), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n486), .A2(new_n209), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT22), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n209), .A2(G87), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n491), .B1(new_n444), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n485), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT24), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n485), .A2(new_n490), .A3(KEYINPUT24), .A4(new_n493), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n496), .A2(new_n318), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n466), .A2(G107), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT83), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n306), .A2(new_n487), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT82), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT25), .ZN(new_n503));
  OR2_X1    g0303(.A1(new_n502), .A2(KEYINPUT25), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n502), .A2(KEYINPUT25), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n504), .A2(new_n306), .A3(new_n505), .A4(new_n487), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n499), .A2(new_n500), .A3(new_n503), .A4(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n503), .B(new_n506), .C1(new_n465), .C2(new_n423), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT83), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n498), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(G250), .A2(G1698), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n512), .B1(new_n218), .B2(G1698), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n484), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(G294), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n514), .B1(new_n515), .B2(new_n369), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n516), .A2(new_n278), .B1(G264), .B2(new_n438), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n342), .A2(new_n439), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n299), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n517), .A2(new_n358), .A3(new_n518), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n511), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AND4_X1   g0322(.A1(new_n480), .A2(new_n482), .A3(new_n483), .A4(new_n522), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n438), .A2(G257), .B1(new_n342), .B2(new_n439), .ZN(new_n524));
  AND2_X1   g0324(.A1(KEYINPUT4), .A2(G244), .ZN(new_n525));
  AND2_X1   g0325(.A1(KEYINPUT3), .A2(G33), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n271), .B(new_n525), .C1(new_n526), .C2(new_n373), .ZN(new_n527));
  OAI211_X1 g0327(.A(G250), .B(G1698), .C1(new_n526), .C2(new_n373), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G33), .A2(G283), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  OAI211_X1 g0330(.A(G244), .B(new_n271), .C1(new_n392), .C2(new_n373), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT4), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n524), .B1(new_n533), .B2(new_n277), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G169), .ZN(new_n535));
  OAI211_X1 g0335(.A(G179), .B(new_n524), .C1(new_n533), .C2(new_n277), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT6), .ZN(new_n537));
  AND2_X1   g0337(.A1(G97), .A2(G107), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n537), .B1(new_n538), .B2(new_n205), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n423), .A2(KEYINPUT6), .A3(G97), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI22_X1  g0341(.A1(new_n541), .A2(new_n209), .B1(new_n338), .B2(new_n315), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n423), .B1(new_n383), .B2(new_n385), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n318), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n307), .A2(G97), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(new_n465), .B2(new_n217), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n535), .A2(new_n536), .B1(new_n544), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n534), .A2(G200), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT76), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n534), .A2(KEYINPUT76), .A3(G200), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n544), .A2(KEYINPUT75), .A3(new_n548), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT75), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n539), .A2(new_n540), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n557), .A2(G20), .B1(G77), .B2(new_n314), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n269), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n559), .B1(new_n369), .B2(new_n266), .ZN(new_n560));
  OAI21_X1  g0360(.A(G107), .B1(new_n560), .B2(new_n384), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n347), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n556), .B1(new_n562), .B2(new_n547), .ZN(new_n563));
  OAI211_X1 g0363(.A(G190), .B(new_n524), .C1(new_n533), .C2(new_n277), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n555), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n549), .B1(new_n554), .B2(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n484), .A2(KEYINPUT78), .A3(G244), .A4(G1698), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT77), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n271), .A2(G238), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n568), .B(new_n570), .C1(new_n392), .C2(new_n373), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n568), .B1(new_n484), .B2(new_n570), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n567), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(G244), .B(G1698), .C1(new_n392), .C2(new_n373), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT78), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n486), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n278), .B1(new_n574), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n437), .A2(G250), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(new_n341), .B2(new_n437), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n254), .A2(new_n258), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n580), .A2(new_n358), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n484), .A2(new_n209), .A3(G68), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT19), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n312), .A2(new_n587), .A3(G97), .ZN(new_n588));
  INV_X1    g0388(.A(G87), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n205), .A2(new_n589), .B1(new_n273), .B2(new_n209), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n588), .B1(new_n590), .B2(new_n587), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n586), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n318), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n466), .A2(new_n414), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n593), .B(new_n594), .C1(new_n307), .C2(new_n414), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n486), .B1(new_n575), .B2(new_n576), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n596), .B(new_n567), .C1(new_n573), .C2(new_n572), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n597), .A2(new_n278), .B1(new_n583), .B2(new_n582), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n585), .B(new_n595), .C1(new_n598), .C2(G169), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n580), .A2(G190), .A3(new_n584), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n593), .B1(new_n307), .B2(new_n414), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n465), .A2(new_n589), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n600), .B(new_n603), .C1(new_n598), .C2(new_n355), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n519), .A2(G200), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n517), .A2(G190), .A3(new_n518), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n605), .A2(new_n510), .A3(new_n498), .A4(new_n606), .ZN(new_n607));
  AND4_X1   g0407(.A1(new_n566), .A2(new_n599), .A3(new_n604), .A4(new_n607), .ZN(new_n608));
  AND4_X1   g0408(.A1(new_n434), .A2(new_n476), .A3(new_n523), .A4(new_n608), .ZN(G372));
  INV_X1    g0409(.A(new_n360), .ZN(new_n610));
  INV_X1    g0410(.A(new_n429), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n327), .B1(new_n330), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n407), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n411), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n610), .B1(new_n614), .B2(new_n357), .ZN(new_n615));
  INV_X1    g0415(.A(new_n599), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n480), .A2(new_n482), .A3(new_n483), .A4(new_n522), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n616), .B1(new_n608), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n535), .A2(new_n536), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n555), .A2(new_n563), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT84), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n619), .A2(new_n620), .A3(KEYINPUT84), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n623), .A2(new_n604), .A3(new_n599), .A4(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT26), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(KEYINPUT85), .A3(new_n626), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n604), .A2(new_n599), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n628), .A2(KEYINPUT26), .A3(new_n549), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(KEYINPUT85), .B1(new_n625), .B2(new_n626), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n618), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n434), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n615), .A2(new_n633), .ZN(G369));
  NAND3_X1  g0434(.A1(new_n480), .A2(new_n482), .A3(new_n483), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT86), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n306), .A2(new_n636), .A3(new_n209), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT86), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT27), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n637), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(G213), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n640), .B1(new_n637), .B2(new_n639), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(G343), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n468), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n635), .A2(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n476), .A2(new_n647), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n648), .B1(new_n649), .B2(new_n635), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(KEYINPUT87), .ZN(new_n651));
  XNOR2_X1  g0451(.A(KEYINPUT88), .B(G330), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT87), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n654), .B(new_n648), .C1(new_n649), .C2(new_n635), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n522), .A2(new_n646), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n511), .A2(new_n646), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n607), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n656), .B1(new_n658), .B2(new_n522), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n651), .A2(new_n653), .A3(new_n655), .A4(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n656), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n659), .A2(new_n635), .A3(new_n645), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(G399));
  INV_X1    g0463(.A(new_n212), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(G41), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(G1), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(new_n225), .B2(new_n666), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n669), .B(KEYINPUT28), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n625), .A2(new_n626), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT85), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n673), .A2(new_n629), .A3(new_n627), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n646), .B1(new_n674), .B2(new_n618), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(KEYINPUT29), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n623), .A2(new_n624), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT92), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n678), .A2(new_n628), .A3(new_n679), .A4(KEYINPUT26), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT92), .B1(new_n625), .B2(new_n626), .ZN(new_n681));
  AOI21_X1  g0481(.A(KEYINPUT26), .B1(new_n628), .B2(new_n549), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n599), .B(new_n680), .C1(new_n681), .C2(new_n682), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n566), .A2(new_n599), .A3(new_n604), .A4(new_n607), .ZN(new_n684));
  OAI21_X1  g0484(.A(KEYINPUT93), .B1(new_n523), .B2(new_n684), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n599), .A2(new_n604), .A3(new_n607), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT93), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n686), .A2(new_n617), .A3(new_n687), .A4(new_n566), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n645), .B1(new_n683), .B2(new_n689), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n690), .A2(KEYINPUT29), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n677), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n580), .A2(new_n517), .A3(new_n584), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT90), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n534), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n580), .A2(KEYINPUT90), .A3(new_n517), .A4(new_n584), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n695), .A2(new_n481), .A3(new_n696), .A4(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT30), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n696), .A2(KEYINPUT30), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n695), .A2(new_n481), .A3(new_n697), .A4(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(KEYINPUT91), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n519), .A2(new_n358), .A3(new_n534), .ZN(new_n705));
  INV_X1    g0505(.A(new_n598), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n451), .A2(new_n453), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n697), .A2(new_n481), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT91), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n710), .A2(new_n711), .A3(new_n695), .A4(new_n702), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n700), .A2(new_n704), .A3(new_n709), .A4(new_n712), .ZN(new_n713));
  XOR2_X1   g0513(.A(KEYINPUT89), .B(KEYINPUT31), .Z(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n713), .A2(new_n646), .A3(new_n715), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n476), .A2(new_n523), .A3(new_n608), .A4(new_n645), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n704), .A2(new_n712), .ZN(new_n718));
  AOI22_X1  g0518(.A1(new_n699), .A2(new_n698), .B1(new_n707), .B2(new_n708), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n645), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  OAI211_X1 g0520(.A(new_n716), .B(new_n717), .C1(new_n720), .C2(KEYINPUT31), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n653), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n692), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n670), .B1(new_n724), .B2(G1), .ZN(G364));
  NOR2_X1   g0525(.A1(new_n358), .A2(G200), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n726), .A2(G20), .A3(G190), .ZN(new_n727));
  INV_X1    g0527(.A(G322), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n209), .A2(G190), .ZN(new_n729));
  NOR2_X1   g0529(.A1(G179), .A2(G200), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(G329), .ZN(new_n732));
  OAI22_X1  g0532(.A1(new_n727), .A2(new_n728), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n729), .A2(new_n726), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  AOI211_X1 g0535(.A(new_n270), .B(new_n733), .C1(G311), .C2(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n399), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n738), .A2(KEYINPUT95), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(KEYINPUT95), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G326), .ZN(new_n743));
  NOR4_X1   g0543(.A1(new_n209), .A2(new_n399), .A3(new_n355), .A4(G179), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n209), .B1(new_n730), .B2(G190), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI22_X1  g0546(.A1(new_n744), .A2(G303), .B1(new_n746), .B2(G294), .ZN(new_n747));
  NOR4_X1   g0547(.A1(new_n209), .A2(new_n355), .A3(G179), .A4(G190), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n737), .A2(G190), .ZN(new_n749));
  XNOR2_X1  g0549(.A(KEYINPUT33), .B(G317), .ZN(new_n750));
  AOI22_X1  g0550(.A1(new_n748), .A2(G283), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n736), .A2(new_n743), .A3(new_n747), .A4(new_n751), .ZN(new_n752));
  XOR2_X1   g0552(.A(new_n745), .B(KEYINPUT97), .Z(new_n753));
  INV_X1    g0553(.A(new_n744), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n270), .B1(new_n754), .B2(new_n589), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT96), .ZN(new_n756));
  AOI22_X1  g0556(.A1(G97), .A2(new_n753), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  OAI221_X1 g0557(.A(new_n757), .B1(new_n756), .B2(new_n755), .C1(new_n201), .C2(new_n741), .ZN(new_n758));
  INV_X1    g0558(.A(new_n727), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n759), .A2(G58), .B1(new_n735), .B2(G77), .ZN(new_n760));
  INV_X1    g0560(.A(G159), .ZN(new_n761));
  OR3_X1    g0561(.A1(new_n731), .A2(KEYINPUT32), .A3(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(KEYINPUT32), .B1(new_n731), .B2(new_n761), .ZN(new_n763));
  AOI22_X1  g0563(.A1(new_n748), .A2(G107), .B1(new_n749), .B2(G68), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n760), .A2(new_n762), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n752), .B1(new_n758), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n231), .B1(G20), .B2(new_n299), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n305), .A2(G20), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n208), .B1(new_n769), .B2(G45), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n665), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n664), .A2(new_n444), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n774), .A2(G355), .B1(new_n457), .B2(new_n664), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n246), .A2(new_n436), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n664), .A2(new_n484), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(G45), .B2(new_n226), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n775), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n767), .ZN(new_n780));
  NOR3_X1   g0580(.A1(G13), .A2(G20), .A3(G33), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT94), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n773), .B1(new_n779), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n768), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n651), .A2(new_n655), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n787), .B1(new_n788), .B2(new_n781), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n651), .A2(new_n653), .A3(new_n655), .ZN(new_n790));
  AND2_X1   g0590(.A1(new_n790), .A2(new_n773), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n788), .A2(new_n652), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n789), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(G396));
  OAI21_X1  g0594(.A(new_n432), .B1(new_n419), .B2(new_n645), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(new_n429), .ZN(new_n796));
  INV_X1    g0596(.A(KEYINPUT99), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n427), .A2(new_n428), .A3(new_n645), .ZN(new_n798));
  AND3_X1   g0598(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n797), .B1(new_n796), .B2(new_n798), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n676), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n632), .A2(new_n645), .A3(new_n801), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT100), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n803), .B(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n772), .B1(new_n807), .B2(new_n722), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n808), .B1(new_n722), .B2(new_n807), .ZN(new_n809));
  NOR2_X1   g0609(.A1(G13), .A2(G33), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n767), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(G77), .ZN(new_n813));
  INV_X1    g0613(.A(new_n748), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(new_n309), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n815), .B1(G50), .B2(new_n744), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n202), .B2(new_n745), .ZN(new_n817));
  INV_X1    g0617(.A(new_n731), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n378), .B(new_n817), .C1(G132), .C2(new_n818), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n759), .A2(G143), .B1(new_n735), .B2(G159), .ZN(new_n820));
  INV_X1    g0620(.A(G150), .ZN(new_n821));
  INV_X1    g0621(.A(new_n749), .ZN(new_n822));
  INV_X1    g0622(.A(G137), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n820), .B1(new_n821), .B2(new_n822), .C1(new_n741), .C2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n819), .B1(KEYINPUT34), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT34), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n748), .A2(G87), .ZN(new_n829));
  INV_X1    g0629(.A(G311), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n829), .B1(new_n830), .B2(new_n731), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT98), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n444), .B1(new_n734), .B2(new_n457), .ZN(new_n833));
  INV_X1    g0633(.A(G283), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n754), .A2(new_n423), .B1(new_n834), .B2(new_n822), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n833), .B(new_n835), .C1(G294), .C2(new_n759), .ZN(new_n836));
  INV_X1    g0636(.A(new_n753), .ZN(new_n837));
  INV_X1    g0637(.A(G303), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n836), .B1(new_n217), .B2(new_n837), .C1(new_n838), .C2(new_n741), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n826), .A2(new_n828), .B1(new_n832), .B2(new_n839), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n773), .B(new_n813), .C1(new_n840), .C2(new_n767), .ZN(new_n841));
  INV_X1    g0641(.A(new_n810), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n841), .B1(new_n801), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n809), .A2(new_n843), .ZN(G384));
  NOR3_X1   g0644(.A1(new_n231), .A2(new_n209), .A3(new_n457), .ZN(new_n845));
  OR2_X1    g0645(.A1(new_n557), .A2(KEYINPUT35), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n557), .A2(KEYINPUT35), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  XOR2_X1   g0648(.A(new_n848), .B(KEYINPUT36), .Z(new_n849));
  OR3_X1    g0649(.A1(new_n363), .A2(new_n225), .A3(new_n338), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n201), .A2(G68), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n208), .B(G13), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(KEYINPUT102), .B1(new_n642), .B2(new_n643), .ZN(new_n854));
  INV_X1    g0654(.A(new_n643), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT102), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n855), .A2(new_n856), .A3(G213), .A4(new_n641), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  OR2_X1    g0659(.A1(new_n411), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n798), .B(KEYINPUT101), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n804), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n326), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT72), .B1(new_n302), .B2(KEYINPUT14), .ZN(new_n865));
  NOR3_X1   g0665(.A1(new_n300), .A2(new_n298), .A3(new_n286), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n287), .B(new_n296), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n864), .B(new_n646), .C1(new_n867), .C2(new_n331), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n864), .A2(new_n646), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n330), .B(new_n869), .C1(new_n304), .C2(new_n326), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n863), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT104), .ZN(new_n873));
  INV_X1    g0673(.A(new_n410), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT103), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n388), .A2(new_n390), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n875), .B1(new_n876), .B2(new_n859), .ZN(new_n877));
  AOI211_X1 g0677(.A(KEYINPUT103), .B(new_n858), .C1(new_n388), .C2(new_n390), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n406), .B(new_n874), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n873), .B1(new_n879), .B2(KEYINPUT37), .ZN(new_n880));
  INV_X1    g0680(.A(new_n877), .ZN(new_n881));
  INV_X1    g0681(.A(new_n878), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n405), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n400), .A2(new_n403), .A3(KEYINPUT74), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n876), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n410), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT37), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n883), .A2(new_n888), .A3(KEYINPUT104), .A4(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n880), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n368), .B1(new_n371), .B2(new_n379), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n892), .A2(new_n381), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n380), .A2(new_n318), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n390), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n409), .A2(new_n408), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n895), .A2(new_n644), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n406), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT37), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n891), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n898), .B1(new_n407), .B2(new_n411), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n901), .A2(KEYINPUT38), .A3(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT38), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n880), .A2(new_n890), .B1(KEYINPUT37), .B2(new_n899), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n905), .B1(new_n906), .B2(new_n902), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n860), .B1(new_n872), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n327), .A2(new_n645), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  XOR2_X1   g0712(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n913));
  AOI22_X1  g0713(.A1(new_n880), .A2(new_n890), .B1(KEYINPUT37), .B2(new_n879), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n883), .B1(new_n407), .B2(new_n411), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT39), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n904), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT106), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n908), .A2(KEYINPUT39), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT106), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n904), .A2(new_n916), .A3(new_n921), .A4(new_n917), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n919), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n910), .B1(new_n912), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n434), .B1(new_n677), .B2(new_n691), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n615), .ZN(new_n926));
  XOR2_X1   g0726(.A(new_n924), .B(new_n926), .Z(new_n927));
  NAND2_X1  g0727(.A1(new_n713), .A2(new_n646), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT108), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n713), .A2(KEYINPUT108), .A3(new_n646), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n930), .A2(new_n714), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n713), .A2(KEYINPUT31), .A3(new_n646), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n717), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n802), .B1(new_n870), .B2(new_n868), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n935), .A2(new_n936), .A3(new_n908), .ZN(new_n937));
  XOR2_X1   g0737(.A(KEYINPUT107), .B(KEYINPUT40), .Z(new_n938));
  NAND2_X1  g0738(.A1(new_n871), .A2(new_n801), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n932), .B2(new_n934), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT40), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n904), .B2(new_n916), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n937), .A2(new_n938), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n434), .A2(new_n935), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n943), .A2(new_n944), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n945), .A2(new_n653), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n927), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n208), .B2(new_n769), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n927), .A2(new_n947), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n853), .B1(new_n949), .B2(new_n950), .ZN(G367));
  NAND2_X1  g0751(.A1(new_n664), .A2(new_n414), .ZN(new_n952));
  INV_X1    g0752(.A(new_n777), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n952), .B1(new_n953), .B2(new_n241), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n772), .B1(new_n784), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n814), .A2(new_n217), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n378), .B1(new_n423), .B2(new_n745), .ZN(new_n957));
  AOI211_X1 g0757(.A(new_n956), .B(new_n957), .C1(G294), .C2(new_n749), .ZN(new_n958));
  INV_X1    g0758(.A(G317), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n727), .A2(new_n838), .B1(new_n731), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(KEYINPUT46), .B1(new_n744), .B2(G116), .ZN(new_n961));
  AOI211_X1 g0761(.A(new_n960), .B(new_n961), .C1(G283), .C2(new_n735), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n744), .A2(KEYINPUT46), .A3(G116), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n742), .A2(G311), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n958), .A2(new_n962), .A3(new_n963), .A4(new_n964), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n727), .A2(new_n821), .B1(new_n734), .B2(new_n201), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n754), .A2(new_n202), .B1(new_n761), .B2(new_n822), .ZN(new_n967));
  XNOR2_X1  g0767(.A(KEYINPUT112), .B(G137), .ZN(new_n968));
  AOI211_X1 g0768(.A(new_n966), .B(new_n967), .C1(new_n818), .C2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n753), .A2(G68), .ZN(new_n970));
  INV_X1    g0770(.A(G143), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n969), .B(new_n970), .C1(new_n971), .C2(new_n741), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n270), .B1(new_n814), .B2(new_n338), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT111), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n965), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT47), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n955), .B1(new_n976), .B2(new_n767), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n646), .B1(new_n601), .B2(new_n602), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n628), .A2(new_n978), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n599), .A2(new_n978), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n977), .B1(new_n981), .B2(new_n782), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n620), .A2(new_n646), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n566), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n619), .A2(new_n620), .A3(new_n646), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n662), .A2(new_n661), .A3(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT45), .Z(new_n988));
  NAND2_X1  g0788(.A1(new_n662), .A2(new_n661), .ZN(new_n989));
  INV_X1    g0789(.A(new_n986), .ZN(new_n990));
  XOR2_X1   g0790(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n991));
  NAND3_X1  g0791(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n986), .B1(new_n662), .B2(new_n661), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n993), .A2(new_n991), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n988), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n660), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n660), .A2(new_n988), .A3(new_n992), .A4(new_n994), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n635), .A2(new_n645), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n659), .B(new_n1000), .Z(new_n1001));
  XNOR2_X1  g0801(.A(new_n790), .B(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n724), .B1(new_n999), .B2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n665), .B(KEYINPUT41), .Z(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT110), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1003), .A2(KEYINPUT110), .A3(new_n1005), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n771), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n990), .A2(new_n522), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1011), .A2(new_n549), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n662), .A2(new_n990), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n1012), .A2(new_n645), .B1(new_n1013), .B2(KEYINPUT42), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(KEYINPUT42), .B2(new_n1013), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n981), .A2(KEYINPUT43), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n981), .A2(KEYINPUT43), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1017), .B(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n996), .A2(new_n986), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1019), .B(new_n1020), .Z(new_n1021));
  OAI21_X1  g0821(.A(new_n982), .B1(new_n1010), .B2(new_n1021), .ZN(G387));
  INV_X1    g0822(.A(new_n1002), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n771), .ZN(new_n1024));
  INV_X1    g0824(.A(G326), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n378), .B1(new_n1025), .B2(new_n731), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n744), .A2(G294), .B1(new_n746), .B2(G283), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n759), .A2(G317), .B1(new_n735), .B2(G303), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n830), .B2(new_n822), .C1(new_n741), .C2(new_n728), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT48), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1027), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT114), .Z(new_n1032));
  INV_X1    g0832(.A(new_n1029), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1032), .B1(KEYINPUT48), .B2(new_n1033), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT49), .Z(new_n1035));
  AOI211_X1 g0835(.A(new_n1026), .B(new_n1035), .C1(G116), .C2(new_n748), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n754), .A2(new_n338), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n956), .B(new_n1037), .C1(new_n349), .C2(new_n749), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n735), .A2(G68), .B1(new_n818), .B2(G150), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1038), .A2(new_n484), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n753), .A2(new_n414), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n201), .B2(new_n727), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT113), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1040), .B(new_n1043), .C1(G159), .C2(new_n742), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n767), .B1(new_n1036), .B2(new_n1044), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n659), .A2(new_n782), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n667), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n774), .A2(new_n1047), .B1(new_n423), .B2(new_n664), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n238), .A2(new_n436), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n349), .A2(new_n201), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT50), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n667), .B(new_n436), .C1(new_n309), .C2(new_n338), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n777), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1048), .B1(new_n1049), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n773), .B1(new_n1054), .B2(new_n785), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1045), .A2(new_n1046), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1002), .A2(new_n723), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(KEYINPUT115), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1002), .A2(new_n723), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1058), .A2(new_n1060), .A3(new_n665), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1057), .A2(KEYINPUT115), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1024), .B(new_n1056), .C1(new_n1061), .C2(new_n1062), .ZN(G393));
  AND2_X1   g0863(.A1(new_n997), .A2(new_n998), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n771), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n777), .A2(new_n249), .B1(G97), .B2(new_n664), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n773), .B1(new_n785), .B2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n837), .A2(new_n338), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n829), .B1(new_n201), .B2(new_n822), .C1(new_n754), .C2(new_n309), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n734), .A2(new_n348), .B1(new_n731), .B2(new_n971), .ZN(new_n1070));
  NOR4_X1   g0870(.A1(new_n1068), .A2(new_n1069), .A3(new_n378), .A4(new_n1070), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n741), .A2(new_n821), .B1(new_n761), .B2(new_n727), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT51), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n741), .A2(new_n959), .B1(new_n830), .B2(new_n727), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT52), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n754), .A2(new_n834), .B1(new_n457), .B2(new_n745), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n444), .B1(new_n731), .B2(new_n728), .C1(new_n515), .C2(new_n734), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n814), .A2(new_n423), .B1(new_n822), .B2(new_n838), .ZN(new_n1078));
  NOR3_X1   g0878(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1071), .A2(new_n1073), .B1(new_n1075), .B2(new_n1079), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1067), .B1(new_n780), .B2(new_n1080), .C1(new_n986), .C2(new_n782), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1065), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n666), .B1(new_n1059), .B2(new_n1064), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1060), .A2(new_n999), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1082), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(G390));
  OAI211_X1 g0886(.A(new_n645), .B(new_n801), .C1(new_n683), .C2(new_n689), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n798), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n871), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT116), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n912), .B1(new_n904), .B2(new_n916), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n868), .A2(new_n870), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n1087), .B2(new_n798), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n913), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n879), .A2(KEYINPUT37), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n891), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n915), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1095), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NOR3_X1   g0899(.A1(new_n906), .A2(new_n905), .A3(new_n902), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n911), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(KEYINPUT116), .B1(new_n1094), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1092), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n861), .B1(new_n675), .B2(new_n801), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n911), .B1(new_n1104), .B2(new_n1093), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1105), .A2(new_n919), .A3(new_n920), .A4(new_n922), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n721), .A2(new_n653), .A3(new_n801), .A4(new_n871), .ZN(new_n1107));
  AND3_X1   g0907(.A1(new_n1103), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(G330), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(new_n932), .B2(new_n934), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n936), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1093), .B1(new_n722), .B2(new_n802), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1104), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n871), .B1(new_n1110), .B2(new_n801), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1107), .A2(new_n798), .A3(new_n1087), .ZN(new_n1116));
  OAI21_X1  g0916(.A(KEYINPUT117), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n1107), .A2(new_n798), .A3(new_n1087), .ZN(new_n1118));
  AND3_X1   g0918(.A1(new_n713), .A2(KEYINPUT108), .A3(new_n646), .ZN(new_n1119));
  AOI21_X1  g0919(.A(KEYINPUT108), .B1(new_n713), .B2(new_n646), .ZN(new_n1120));
  NOR3_X1   g0920(.A1(new_n1119), .A2(new_n1120), .A3(new_n715), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n717), .A2(new_n933), .ZN(new_n1122));
  OAI211_X1 g0922(.A(G330), .B(new_n801), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n1093), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT117), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1118), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1114), .B1(new_n1117), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n434), .A2(new_n1110), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n925), .A2(new_n615), .A3(new_n1128), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n1108), .A2(new_n1112), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1114), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1125), .B1(new_n1118), .B2(new_n1124), .ZN(new_n1132));
  NOR3_X1   g0932(.A1(new_n1115), .A2(new_n1116), .A3(KEYINPUT117), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1131), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1090), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n1094), .A2(new_n1101), .A3(KEYINPUT116), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n912), .B1(new_n863), .B2(new_n871), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n1135), .A2(new_n1136), .B1(new_n923), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1111), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1103), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1129), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1134), .A2(new_n1140), .A3(new_n1141), .A4(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1130), .A2(new_n1143), .A3(new_n665), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1108), .A2(new_n1112), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n923), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n810), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n772), .B1(new_n812), .B2(new_n349), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1068), .B1(G283), .B2(new_n742), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n734), .A2(new_n217), .B1(new_n731), .B2(new_n515), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n270), .B(new_n1150), .C1(G116), .C2(new_n759), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n822), .A2(new_n423), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n1152), .B(new_n815), .C1(G87), .C2(new_n744), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1149), .A2(new_n1151), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n744), .A2(G150), .ZN(new_n1155));
  XOR2_X1   g0955(.A(new_n1155), .B(KEYINPUT53), .Z(new_n1156));
  INV_X1    g0956(.A(G132), .ZN(new_n1157));
  INV_X1    g0957(.A(G125), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n727), .A2(new_n1157), .B1(new_n731), .B2(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(KEYINPUT54), .B(G143), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n444), .B(new_n1159), .C1(new_n735), .C2(new_n1161), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n748), .A2(G50), .B1(new_n749), .B2(new_n968), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1156), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(G128), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n837), .A2(new_n761), .B1(new_n741), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1154), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1148), .B1(new_n1167), .B2(new_n767), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n1145), .A2(new_n771), .B1(new_n1147), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1144), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT118), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1144), .A2(new_n1169), .A3(KEYINPUT118), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(G378));
  INV_X1    g0975(.A(new_n924), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n937), .A2(new_n938), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n940), .A2(new_n942), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1177), .A2(new_n1178), .A3(G330), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n361), .A2(new_n353), .A3(new_n644), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n361), .B1(new_n353), .B2(new_n644), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  OR3_X1    g0983(.A1(new_n1180), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1183), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1179), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(new_n943), .B2(G330), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1176), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1179), .A2(new_n1186), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n943), .A2(G330), .A3(new_n1188), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1191), .A2(new_n1192), .A3(new_n924), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1190), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1186), .A2(new_n810), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n772), .B1(new_n812), .B2(G50), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n822), .A2(new_n217), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1197), .B(new_n1037), .C1(G58), .C2(new_n748), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n759), .A2(G107), .B1(new_n735), .B2(new_n414), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n834), .B2(new_n731), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n484), .A2(G41), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n742), .A2(G116), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1198), .A2(new_n1203), .A3(new_n970), .A4(new_n1204), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT58), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1202), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n822), .A2(new_n1157), .B1(new_n734), .B2(new_n823), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT119), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n759), .A2(G128), .B1(new_n744), .B2(new_n1161), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n837), .B2(new_n821), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1209), .B(new_n1211), .C1(G125), .C2(new_n742), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(KEYINPUT59), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n748), .A2(G159), .ZN(new_n1215));
  AOI211_X1 g1015(.A(G33), .B(G41), .C1(new_n818), .C2(G124), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1213), .A2(KEYINPUT59), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1206), .B(new_n1207), .C1(new_n1217), .C2(new_n1218), .ZN(new_n1219));
  OR2_X1    g1019(.A1(new_n1219), .A2(KEYINPUT120), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n780), .B1(new_n1219), .B2(KEYINPUT120), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1196), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1194), .A2(new_n771), .B1(new_n1195), .B2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1129), .B1(new_n1145), .B2(new_n1134), .ZN(new_n1224));
  AND3_X1   g1024(.A1(new_n1191), .A2(new_n1192), .A3(new_n924), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n924), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1226));
  OAI21_X1  g1026(.A(KEYINPUT57), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n665), .B1(new_n1224), .B2(new_n1227), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n1146), .A2(new_n1105), .B1(new_n1092), .B2(new_n1102), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1141), .B1(new_n1229), .B2(new_n1111), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1142), .B1(new_n1230), .B2(new_n1127), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT57), .B1(new_n1231), .B2(new_n1194), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1223), .B1(new_n1228), .B2(new_n1232), .ZN(G375));
  NAND2_X1  g1033(.A1(new_n1134), .A2(new_n1142), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1131), .B(new_n1129), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1234), .A2(new_n1005), .A3(new_n1235), .ZN(new_n1236));
  XOR2_X1   g1036(.A(new_n1236), .B(KEYINPUT121), .Z(new_n1237));
  NAND2_X1  g1037(.A1(new_n1093), .A2(new_n810), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n772), .B1(new_n812), .B2(G68), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n734), .A2(new_n423), .B1(new_n731), .B2(new_n838), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n270), .B(new_n1240), .C1(G283), .C2(new_n759), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n814), .A2(new_n338), .B1(new_n822), .B2(new_n457), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(G97), .B2(new_n744), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n742), .A2(G294), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1241), .A2(new_n1041), .A3(new_n1243), .A4(new_n1244), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n759), .A2(new_n968), .B1(new_n1161), .B2(new_n749), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n741), .B2(new_n1157), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(KEYINPUT122), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n753), .A2(G50), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n735), .A2(G150), .B1(new_n818), .B2(G128), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n744), .A2(G159), .B1(new_n748), .B2(G58), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1249), .A2(new_n484), .A3(new_n1250), .A4(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1245), .B1(new_n1248), .B2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1239), .B1(new_n1253), .B2(new_n767), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n1134), .A2(new_n771), .B1(new_n1238), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1237), .A2(new_n1255), .ZN(G381));
  INV_X1    g1056(.A(G384), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1085), .A2(new_n1257), .ZN(new_n1258));
  NOR4_X1   g1058(.A1(G387), .A2(G396), .A3(G393), .A4(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT123), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1170), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1144), .A2(new_n1169), .A3(KEYINPUT123), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1263), .A2(G375), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1259), .A2(new_n1264), .A3(new_n1255), .A4(new_n1237), .ZN(G407));
  INV_X1    g1065(.A(G213), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1266), .A2(G343), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1264), .A2(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(G407), .A2(G213), .A3(new_n1268), .ZN(G409));
  NAND3_X1  g1069(.A1(new_n1231), .A2(new_n1194), .A3(new_n1005), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1223), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1261), .A2(new_n1262), .A3(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n1174), .B2(G375), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT60), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1235), .A2(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1127), .A2(KEYINPUT60), .A3(new_n1129), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1275), .A2(new_n1234), .A3(new_n1276), .A4(new_n665), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1277), .A2(G384), .A3(new_n1255), .ZN(new_n1278));
  AOI21_X1  g1078(.A(G384), .B1(new_n1277), .B2(new_n1255), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n1280), .A2(KEYINPUT63), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1267), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1273), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT127), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1273), .A2(new_n1281), .A3(KEYINPUT127), .A4(new_n1282), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(G393), .B(G396), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n1003), .A2(KEYINPUT110), .A3(new_n1005), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT110), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n770), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(new_n1019), .B(new_n1020), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(G390), .B1(new_n1293), .B2(new_n982), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n982), .ZN(new_n1295));
  AOI211_X1 g1095(.A(new_n1295), .B(new_n1085), .C1(new_n1291), .C2(new_n1292), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1288), .B1(new_n1294), .B2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(G387), .A2(new_n1085), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(G393), .B(new_n793), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1293), .A2(new_n982), .A3(G390), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1298), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT61), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1297), .A2(new_n1301), .A3(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(G2897), .ZN(new_n1304));
  OAI22_X1  g1104(.A1(new_n1278), .A2(new_n1279), .B1(new_n1304), .B2(new_n1282), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1277), .A2(new_n1255), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1257), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1277), .A2(G384), .A3(new_n1255), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1282), .A2(new_n1304), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1307), .A2(new_n1308), .A3(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1305), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT126), .ZN(new_n1312));
  AOI22_X1  g1112(.A1(new_n1273), .A2(new_n1282), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1305), .A2(new_n1310), .A3(KEYINPUT126), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1303), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT125), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1231), .A2(new_n1194), .A3(KEYINPUT57), .ZN(new_n1318));
  AOI22_X1  g1118(.A1(new_n1143), .A2(new_n1142), .B1(new_n1190), .B2(new_n1193), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1318), .B(new_n665), .C1(new_n1319), .C2(KEYINPUT57), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1320), .A2(new_n1172), .A3(new_n1173), .A4(new_n1223), .ZN(new_n1321));
  AOI211_X1 g1121(.A(new_n1267), .B(new_n1317), .C1(new_n1321), .C2(new_n1272), .ZN(new_n1322));
  XNOR2_X1  g1122(.A(KEYINPUT124), .B(KEYINPUT63), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1316), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1273), .A2(new_n1282), .A3(new_n1280), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1323), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1325), .A2(KEYINPUT125), .A3(new_n1326), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1287), .A2(new_n1315), .A3(new_n1324), .A4(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1325), .A2(KEYINPUT62), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1273), .A2(new_n1282), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n1311), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT62), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1273), .A2(new_n1332), .A3(new_n1282), .A4(new_n1280), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1329), .A2(new_n1331), .A3(new_n1302), .A4(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1297), .A2(new_n1301), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1328), .A2(new_n1336), .ZN(G405));
  NAND3_X1  g1137(.A1(G375), .A2(new_n1261), .A3(new_n1262), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1338), .A2(new_n1321), .ZN(new_n1339));
  XNOR2_X1  g1139(.A(new_n1339), .B(new_n1280), .ZN(new_n1340));
  XNOR2_X1  g1140(.A(new_n1340), .B(new_n1335), .ZN(G402));
endmodule


