//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 1 0 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 0 1 0 0 1 0 1 1 0 0 0 0 1 0 0 0 1 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n822, new_n823, new_n825, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(G57gat), .B(G85gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(G127gat), .ZN(new_n206));
  INV_X1    g005(.A(G134gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G113gat), .ZN(new_n209));
  INV_X1    g008(.A(G120gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT1), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n212), .B1(G113gat), .B2(G120gat), .ZN(new_n213));
  XNOR2_X1  g012(.A(KEYINPUT67), .B(G127gat), .ZN(new_n214));
  OAI221_X1 g013(.A(new_n208), .B1(new_n211), .B2(new_n213), .C1(new_n214), .C2(new_n207), .ZN(new_n215));
  INV_X1    g014(.A(new_n213), .ZN(new_n216));
  XNOR2_X1  g015(.A(G127gat), .B(G134gat), .ZN(new_n217));
  XOR2_X1   g016(.A(KEYINPUT68), .B(G120gat), .Z(new_n218));
  OAI211_X1 g017(.A(new_n216), .B(new_n217), .C1(new_n218), .C2(new_n209), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT83), .ZN(new_n222));
  INV_X1    g021(.A(G141gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n223), .A2(G148gat), .ZN(new_n224));
  AND2_X1   g023(.A1(KEYINPUT81), .A2(G141gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(KEYINPUT81), .A2(G141gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n224), .B1(new_n227), .B2(G148gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT82), .ZN(new_n229));
  INV_X1    g028(.A(G155gat), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT2), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G162gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G155gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n230), .A2(G162gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n231), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n222), .B1(new_n228), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n235), .ZN(new_n237));
  INV_X1    g036(.A(new_n224), .ZN(new_n238));
  XNOR2_X1  g037(.A(KEYINPUT81), .B(G141gat), .ZN(new_n239));
  INV_X1    g038(.A(G148gat), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n237), .A2(new_n241), .A3(KEYINPUT83), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n236), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n233), .A2(new_n234), .ZN(new_n244));
  XNOR2_X1  g043(.A(G141gat), .B(G148gat), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n244), .B1(new_n245), .B2(KEYINPUT2), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n221), .B1(new_n247), .B2(KEYINPUT3), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n243), .A2(new_n249), .A3(new_n246), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(G225gat), .A2(G233gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n253), .A2(KEYINPUT5), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT85), .ZN(new_n255));
  AND2_X1   g054(.A1(new_n236), .A2(new_n242), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n215), .A2(new_n219), .A3(new_n246), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n243), .A2(new_n221), .A3(KEYINPUT85), .A4(new_n246), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(KEYINPUT4), .A3(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT86), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n256), .A2(new_n257), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT84), .B(KEYINPUT4), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n258), .A2(KEYINPUT86), .A3(new_n259), .A4(KEYINPUT4), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n262), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n254), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n247), .A2(new_n220), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n258), .A2(new_n269), .A3(new_n259), .ZN(new_n270));
  INV_X1    g069(.A(new_n252), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT4), .B1(new_n258), .B2(new_n259), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n263), .A2(new_n264), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI211_X1 g074(.A(KEYINPUT5), .B(new_n272), .C1(new_n275), .C2(new_n253), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n205), .B1(new_n268), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT87), .B(KEYINPUT6), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT96), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n277), .A2(KEYINPUT96), .A3(new_n279), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n277), .A2(new_n279), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n268), .A2(new_n205), .A3(new_n276), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  XOR2_X1   g087(.A(G211gat), .B(G218gat), .Z(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G197gat), .B(G204gat), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT22), .ZN(new_n292));
  INV_X1    g091(.A(G211gat), .ZN(new_n293));
  INV_X1    g092(.A(G218gat), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT29), .B1(new_n290), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n297), .B1(new_n290), .B2(new_n296), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT89), .ZN(new_n299));
  OR2_X1    g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n299), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(new_n249), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(new_n247), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT29), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n250), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n289), .A2(KEYINPUT74), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n306), .B(new_n296), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G228gat), .A2(G233gat), .ZN(new_n310));
  XOR2_X1   g109(.A(new_n310), .B(KEYINPUT88), .Z(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n249), .B1(new_n307), .B2(KEYINPUT29), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n310), .B1(new_n313), .B2(new_n247), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n308), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G22gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n316), .A2(G22gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT90), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n322), .B1(new_n317), .B2(new_n318), .ZN(new_n323));
  XNOR2_X1  g122(.A(G78gat), .B(G106gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(KEYINPUT31), .B(G50gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n324), .B(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n321), .B1(new_n323), .B2(new_n327), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n319), .A2(new_n322), .A3(new_n320), .A4(new_n326), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT35), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n288), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT73), .ZN(new_n333));
  INV_X1    g132(.A(G183gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT27), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT27), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(G183gat), .ZN(new_n337));
  INV_X1    g136(.A(G190gat), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n335), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT28), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT65), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT66), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n343), .B1(new_n339), .B2(new_n340), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT27), .B(G183gat), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n345), .A2(KEYINPUT66), .A3(KEYINPUT28), .A4(new_n338), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT65), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n339), .A2(new_n347), .A3(new_n340), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n342), .A2(new_n344), .A3(new_n346), .A4(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G169gat), .A2(G176gat), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(G169gat), .ZN(new_n352));
  INV_X1    g151(.A(G176gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n351), .B1(KEYINPUT26), .B2(new_n354), .ZN(new_n355));
  OR2_X1    g154(.A1(new_n354), .A2(KEYINPUT26), .ZN(new_n356));
  AOI22_X1  g155(.A1(new_n355), .A2(new_n356), .B1(G183gat), .B2(G190gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n349), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT64), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT24), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(G183gat), .A3(G190gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(G183gat), .B(G190gat), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n359), .B(new_n361), .C1(new_n362), .C2(new_n360), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT25), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n361), .B1(new_n362), .B2(new_n360), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n352), .A2(new_n353), .A3(KEYINPUT23), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT23), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n367), .B1(G169gat), .B2(G176gat), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n366), .A2(new_n368), .A3(new_n350), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n363), .B(new_n364), .C1(new_n365), .C2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n361), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n334), .A2(G190gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n338), .A2(G183gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n371), .B1(new_n374), .B2(KEYINPUT24), .ZN(new_n375));
  INV_X1    g174(.A(new_n369), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n375), .B(new_n376), .C1(new_n359), .C2(KEYINPUT25), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n370), .A2(new_n377), .ZN(new_n378));
  AND2_X1   g177(.A1(new_n358), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(new_n220), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n220), .B1(new_n358), .B2(new_n378), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(G227gat), .ZN(new_n383));
  INV_X1    g182(.A(G233gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n380), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT33), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT69), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT69), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n386), .A2(new_n390), .A3(new_n387), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  AND2_X1   g191(.A1(new_n386), .A2(KEYINPUT32), .ZN(new_n393));
  XNOR2_X1  g192(.A(G15gat), .B(G43gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(G71gat), .B(G99gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n392), .A2(new_n397), .ZN(new_n398));
  OR2_X1    g197(.A1(new_n396), .A2(new_n387), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n393), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n385), .A2(KEYINPUT34), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n358), .A2(new_n378), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n403), .A2(new_n221), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n402), .B1(new_n404), .B2(new_n381), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n380), .A2(KEYINPUT71), .A3(new_n382), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT71), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n407), .B1(new_n404), .B2(new_n381), .ZN(new_n408));
  INV_X1    g207(.A(new_n385), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n406), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT72), .ZN(new_n411));
  XOR2_X1   g210(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n412));
  NAND3_X1  g211(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n411), .B1(new_n410), .B2(new_n412), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n405), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n333), .B1(new_n401), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n416), .ZN(new_n418));
  AOI22_X1  g217(.A1(new_n392), .A2(new_n397), .B1(new_n393), .B2(new_n399), .ZN(new_n419));
  INV_X1    g218(.A(new_n415), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n413), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n419), .A2(new_n421), .A3(KEYINPUT73), .A4(new_n405), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n417), .A2(new_n418), .A3(new_n422), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n332), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT92), .ZN(new_n425));
  XOR2_X1   g224(.A(G8gat), .B(G36gat), .Z(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(KEYINPUT79), .ZN(new_n427));
  XNOR2_X1  g226(.A(G64gat), .B(G92gat), .ZN(new_n428));
  XOR2_X1   g227(.A(new_n427), .B(new_n428), .Z(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n307), .ZN(new_n431));
  NAND2_X1  g230(.A1(G226gat), .A2(G233gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(KEYINPUT75), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  OAI211_X1 g233(.A(KEYINPUT77), .B(new_n434), .C1(new_n379), .C2(KEYINPUT29), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT77), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT29), .B1(new_n358), .B2(new_n378), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n436), .B1(new_n437), .B2(new_n433), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT78), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT76), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n358), .A2(new_n441), .A3(new_n378), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n441), .B1(new_n358), .B2(new_n378), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n440), .B1(new_n444), .B2(new_n433), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n403), .A2(KEYINPUT76), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n358), .A2(new_n441), .A3(new_n378), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n446), .A2(new_n440), .A3(new_n433), .A4(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n431), .B(new_n439), .C1(new_n445), .C2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n403), .A2(new_n433), .ZN(new_n451));
  NOR3_X1   g250(.A1(new_n442), .A2(new_n443), .A3(KEYINPUT29), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n451), .B1(new_n452), .B2(new_n433), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n307), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n430), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n446), .A2(new_n304), .A3(new_n447), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n434), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n431), .B1(new_n458), .B2(new_n451), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n446), .A2(new_n433), .A3(new_n447), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT78), .ZN(new_n461));
  AOI22_X1  g260(.A1(new_n461), .A2(new_n448), .B1(new_n438), .B2(new_n435), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n459), .B1(new_n462), .B2(new_n431), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT80), .B1(new_n463), .B2(new_n430), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT30), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n456), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n450), .A2(new_n454), .A3(new_n430), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT80), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n467), .A2(new_n468), .A3(new_n465), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n425), .B1(new_n466), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n467), .A2(new_n468), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n455), .B1(new_n472), .B2(KEYINPUT30), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n473), .A2(KEYINPUT92), .A3(new_n469), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n424), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n473), .A2(new_n469), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n287), .A2(new_n280), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n419), .A2(new_n421), .A3(new_n405), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n418), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n478), .A2(new_n479), .A3(new_n481), .A4(new_n330), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT35), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n476), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT91), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n418), .A2(new_n480), .A3(KEYINPUT36), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT36), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n486), .B1(new_n487), .B2(new_n423), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n330), .B1(new_n478), .B2(new_n479), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n485), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n423), .A2(new_n487), .ZN(new_n491));
  INV_X1    g290(.A(new_n486), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n330), .ZN(new_n494));
  INV_X1    g293(.A(new_n479), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n494), .B1(new_n495), .B2(new_n477), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n493), .A2(new_n496), .A3(KEYINPUT91), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n490), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT37), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n430), .B1(new_n463), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n462), .A2(new_n307), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n499), .B1(new_n453), .B2(new_n431), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT38), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT95), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n500), .A2(KEYINPUT95), .A3(new_n503), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n282), .A2(new_n283), .B1(new_n286), .B2(new_n285), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n463), .A2(new_n499), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(new_n429), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n463), .A2(new_n499), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT38), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n510), .A2(new_n514), .A3(new_n467), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n330), .B1(new_n509), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT94), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT39), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT93), .ZN(new_n519));
  AOI211_X1 g318(.A(new_n519), .B(new_n252), .C1(new_n267), .C2(new_n251), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n260), .A2(new_n261), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n266), .A2(new_n265), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n251), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT93), .B1(new_n523), .B2(new_n271), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n518), .B1(new_n520), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n251), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n266), .A2(new_n265), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n526), .B1(new_n527), .B2(new_n262), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n519), .B1(new_n528), .B2(new_n252), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n523), .A2(KEYINPUT93), .A3(new_n271), .ZN(new_n530));
  INV_X1    g329(.A(new_n270), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n518), .B1(new_n531), .B2(new_n252), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n529), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n525), .A2(new_n205), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT40), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n277), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n525), .A2(new_n533), .A3(KEYINPUT40), .A4(new_n205), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n517), .B1(new_n475), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n541));
  NOR4_X1   g340(.A1(new_n470), .A2(new_n541), .A3(new_n425), .A4(new_n455), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT92), .B1(new_n473), .B2(new_n469), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n538), .A2(new_n537), .ZN(new_n545));
  INV_X1    g344(.A(new_n205), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n529), .A2(new_n530), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n546), .B1(new_n547), .B2(new_n518), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT40), .B1(new_n548), .B2(new_n533), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n544), .A2(new_n550), .A3(KEYINPUT94), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n516), .B1(new_n540), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n484), .B1(new_n498), .B2(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(G43gat), .B(G50gat), .Z(new_n554));
  INV_X1    g353(.A(KEYINPUT15), .ZN(new_n555));
  OAI21_X1  g354(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n556));
  OR3_X1    g355(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n557));
  AOI22_X1  g356(.A1(new_n554), .A2(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G43gat), .B(G50gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT15), .ZN(new_n560));
  NAND2_X1  g359(.A1(G29gat), .A2(G36gat), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n558), .A2(KEYINPUT99), .A3(new_n560), .A4(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT99), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n560), .A2(new_n561), .ZN(new_n564));
  INV_X1    g363(.A(new_n556), .ZN(new_n565));
  NOR3_X1   g364(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n566));
  OAI22_X1  g365(.A1(new_n559), .A2(KEYINPUT15), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n563), .B1(new_n564), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n562), .A2(new_n568), .ZN(new_n569));
  OR2_X1    g368(.A1(new_n556), .A2(KEYINPUT98), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n556), .A2(KEYINPUT98), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n570), .A2(new_n557), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n560), .B1(new_n572), .B2(new_n561), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G15gat), .B(G22gat), .ZN(new_n576));
  OR2_X1    g375(.A1(new_n576), .A2(G1gat), .ZN(new_n577));
  INV_X1    g376(.A(G8gat), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT16), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n576), .B1(new_n579), .B2(G1gat), .ZN(new_n580));
  AND3_X1   g379(.A1(new_n577), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n578), .B1(new_n577), .B2(new_n580), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n575), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G229gat), .A2(G233gat), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n573), .B1(new_n562), .B2(new_n568), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n583), .B1(new_n587), .B2(KEYINPUT17), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT17), .ZN(new_n589));
  AOI211_X1 g388(.A(new_n589), .B(new_n573), .C1(new_n568), .C2(new_n562), .ZN(new_n590));
  OAI211_X1 g389(.A(new_n585), .B(new_n586), .C1(new_n588), .C2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT100), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n592), .A2(KEYINPUT18), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n575), .A2(new_n589), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n587), .A2(KEYINPUT17), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n596), .A2(new_n583), .A3(new_n597), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n598), .A2(new_n585), .A3(new_n586), .A4(new_n593), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n586), .B(KEYINPUT13), .Z(new_n601));
  NOR2_X1   g400(.A1(new_n575), .A2(new_n584), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n587), .A2(new_n583), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT101), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI211_X1 g405(.A(KEYINPUT101), .B(new_n601), .C1(new_n602), .C2(new_n603), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G113gat), .B(G141gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(G197gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(KEYINPUT11), .B(G169gat), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n610), .B(new_n611), .Z(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT12), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n600), .A2(new_n608), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(KEYINPUT102), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT102), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n600), .A2(new_n608), .A3(new_n616), .A4(new_n613), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n600), .A2(new_n608), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n613), .B(KEYINPUT97), .Z(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  AND2_X1   g421(.A1(G232gat), .A2(G233gat), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n623), .A2(KEYINPUT41), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT7), .ZN(new_n626));
  INV_X1    g425(.A(G85gat), .ZN(new_n627));
  OAI21_X1  g426(.A(G92gat), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(G92gat), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n629), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n630));
  AOI22_X1  g429(.A1(new_n628), .A2(new_n630), .B1(new_n626), .B2(new_n627), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT8), .ZN(new_n632));
  NAND2_X1  g431(.A1(G99gat), .A2(G106gat), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n632), .B1(new_n633), .B2(KEYINPUT107), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n634), .B1(KEYINPUT107), .B2(new_n633), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(G99gat), .B(G106gat), .Z(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n637), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n631), .A2(new_n639), .A3(new_n635), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n596), .A2(new_n597), .A3(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n641), .ZN(new_n643));
  AOI22_X1  g442(.A1(new_n575), .A2(new_n643), .B1(KEYINPUT41), .B2(new_n623), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(G190gat), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n642), .A2(new_n338), .A3(new_n644), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(KEYINPUT106), .B1(new_n648), .B2(new_n294), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n646), .A2(G218gat), .A3(new_n647), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n625), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT106), .ZN(new_n652));
  INV_X1    g451(.A(new_n647), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n338), .B1(new_n642), .B2(new_n644), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n294), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  AND4_X1   g454(.A1(new_n652), .A2(new_n655), .A3(new_n625), .A4(new_n650), .ZN(new_n656));
  XOR2_X1   g455(.A(G134gat), .B(G162gat), .Z(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NOR3_X1   g457(.A1(new_n651), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n655), .A2(new_n652), .A3(new_n650), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(new_n624), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n649), .A2(new_n625), .A3(new_n650), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n657), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g463(.A(G57gat), .B(G64gat), .Z(new_n665));
  NAND2_X1  g464(.A1(G71gat), .A2(G78gat), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT9), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(G71gat), .ZN(new_n670));
  INV_X1    g469(.A(G78gat), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n672), .A2(KEYINPUT103), .A3(new_n666), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n666), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT103), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n669), .A2(new_n673), .A3(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n674), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n678), .A2(new_n665), .A3(KEYINPUT103), .A4(new_n668), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n680), .A2(KEYINPUT21), .ZN(new_n681));
  NAND2_X1  g480(.A1(G231gat), .A2(G233gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(new_n206), .ZN(new_n684));
  AND3_X1   g483(.A1(new_n677), .A2(KEYINPUT105), .A3(new_n679), .ZN(new_n685));
  AOI21_X1  g484(.A(KEYINPUT105), .B1(new_n677), .B2(new_n679), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT21), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n583), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n684), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT104), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(G155gat), .ZN(new_n693));
  XOR2_X1   g492(.A(G183gat), .B(G211gat), .Z(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n690), .B(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n664), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT108), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n638), .A2(KEYINPUT10), .A3(new_n640), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n699), .B1(new_n687), .B2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT10), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n641), .A2(new_n680), .ZN(new_n703));
  AOI22_X1  g502(.A1(new_n638), .A2(new_n640), .B1(new_n677), .B2(new_n679), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n700), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n706), .B(KEYINPUT108), .C1(new_n685), .C2(new_n686), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n701), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(G230gat), .A2(G233gat), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  OR3_X1    g509(.A1(new_n703), .A2(new_n709), .A3(new_n704), .ZN(new_n711));
  XOR2_X1   g510(.A(G120gat), .B(G148gat), .Z(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT109), .ZN(new_n713));
  XNOR2_X1  g512(.A(G176gat), .B(G204gat), .ZN(new_n714));
  XOR2_X1   g513(.A(new_n713), .B(new_n714), .Z(new_n715));
  NAND3_X1  g514(.A1(new_n710), .A2(new_n711), .A3(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT110), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n710), .A2(KEYINPUT110), .A3(new_n711), .A4(new_n715), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n710), .A2(new_n711), .ZN(new_n721));
  INV_X1    g520(.A(new_n715), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n698), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n553), .A2(new_n622), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(KEYINPUT111), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT111), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n553), .A2(new_n728), .A3(new_n622), .A4(new_n725), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n495), .ZN(new_n731));
  XNOR2_X1  g530(.A(KEYINPUT112), .B(G1gat), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n731), .B(new_n732), .ZN(G1324gat));
  XNOR2_X1  g532(.A(KEYINPUT16), .B(G8gat), .ZN(new_n734));
  AOI211_X1 g533(.A(new_n475), .B(new_n734), .C1(new_n727), .C2(new_n729), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n735), .A2(KEYINPUT42), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n578), .B1(new_n730), .B2(new_n544), .ZN(new_n737));
  OAI21_X1  g536(.A(KEYINPUT42), .B1(new_n737), .B2(new_n735), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(G1325gat));
  NOR2_X1   g538(.A1(new_n423), .A2(G15gat), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n730), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(G15gat), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n493), .B1(new_n727), .B2(new_n729), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT113), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT113), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n741), .B(new_n746), .C1(new_n742), .C2(new_n743), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(G1326gat));
  NAND2_X1  g547(.A1(new_n730), .A2(new_n494), .ZN(new_n749));
  XNOR2_X1  g548(.A(KEYINPUT43), .B(G22gat), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n749), .B(new_n750), .ZN(G1327gat));
  NAND2_X1  g550(.A1(new_n553), .A2(new_n622), .ZN(new_n752));
  INV_X1    g551(.A(new_n724), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n696), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n664), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  NOR4_X1   g555(.A1(new_n752), .A2(G29gat), .A3(new_n479), .A4(new_n756), .ZN(new_n757));
  OR2_X1    g556(.A1(new_n757), .A2(KEYINPUT45), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(KEYINPUT45), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n488), .A2(new_n489), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n484), .B1(new_n552), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n658), .B1(new_n651), .B2(new_n656), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n661), .A2(new_n662), .A3(new_n657), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT44), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n664), .A2(new_n767), .ZN(new_n768));
  AOI22_X1  g567(.A1(new_n766), .A2(new_n767), .B1(new_n553), .B2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n622), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n754), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(KEYINPUT114), .B1(new_n772), .B2(new_n479), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(G29gat), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n772), .A2(KEYINPUT114), .A3(new_n479), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n758), .B(new_n759), .C1(new_n774), .C2(new_n775), .ZN(G1328gat));
  NOR4_X1   g575(.A1(new_n752), .A2(G36gat), .A3(new_n475), .A4(new_n756), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(KEYINPUT46), .ZN(new_n778));
  OAI21_X1  g577(.A(G36gat), .B1(new_n772), .B2(new_n475), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(G1329gat));
  AOI22_X1  g579(.A1(new_n424), .A2(new_n475), .B1(KEYINPUT35), .B2(new_n482), .ZN(new_n781));
  INV_X1    g580(.A(new_n515), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n494), .B1(new_n782), .B2(new_n508), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n475), .A2(new_n517), .A3(new_n539), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT94), .B1(new_n544), .B2(new_n550), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n783), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n781), .B1(new_n786), .B2(new_n760), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n767), .B1(new_n787), .B2(new_n664), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n553), .A2(new_n768), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n788), .A2(new_n488), .A3(new_n789), .A4(new_n771), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(G43gat), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n423), .A2(G43gat), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n752), .A2(new_n756), .A3(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n791), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT47), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n794), .B1(new_n790), .B2(G43gat), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT47), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n799), .A2(KEYINPUT115), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n798), .A2(new_n801), .ZN(G1330gat));
  NAND4_X1  g601(.A1(new_n788), .A2(new_n494), .A3(new_n789), .A4(new_n771), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(G50gat), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n330), .A2(G50gat), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n553), .A2(new_n622), .A3(new_n755), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT48), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n807), .B(new_n808), .ZN(G1331gat));
  NOR3_X1   g608(.A1(new_n698), .A2(new_n622), .A3(new_n753), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n762), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n495), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g613(.A1(new_n811), .A2(new_n475), .ZN(new_n815));
  NOR2_X1   g614(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n816));
  AND2_X1   g615(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n818), .B1(new_n815), .B2(new_n816), .ZN(G1333gat));
  OAI21_X1  g618(.A(G71gat), .B1(new_n811), .B2(new_n493), .ZN(new_n820));
  INV_X1    g619(.A(new_n423), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n670), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n820), .B1(new_n811), .B2(new_n822), .ZN(new_n823));
  XOR2_X1   g622(.A(new_n823), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g623(.A1(new_n811), .A2(new_n330), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(new_n671), .ZN(G1335gat));
  NOR2_X1   g625(.A1(new_n697), .A2(new_n622), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n724), .ZN(new_n828));
  XOR2_X1   g627(.A(new_n828), .B(KEYINPUT116), .Z(new_n829));
  NAND2_X1  g628(.A1(new_n769), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(G85gat), .B1(new_n830), .B2(new_n479), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n787), .A2(new_n664), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT117), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n832), .A2(new_n833), .A3(KEYINPUT51), .A4(new_n827), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n762), .A2(new_n765), .A3(new_n827), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT51), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT117), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n836), .ZN(new_n838));
  AND3_X1   g637(.A1(new_n834), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n495), .A2(new_n627), .A3(new_n724), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n831), .B1(new_n839), .B2(new_n840), .ZN(G1336gat));
  NAND4_X1  g640(.A1(new_n788), .A2(new_n544), .A3(new_n789), .A4(new_n829), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT52), .B1(new_n842), .B2(G92gat), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n475), .A2(G92gat), .A3(new_n753), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n843), .B1(new_n839), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT118), .ZN(new_n847));
  AND3_X1   g646(.A1(new_n835), .A2(new_n847), .A3(KEYINPUT51), .ZN(new_n848));
  AOI21_X1  g647(.A(KEYINPUT51), .B1(new_n835), .B2(new_n847), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI22_X1  g649(.A1(new_n850), .A2(new_n844), .B1(G92gat), .B2(new_n842), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT52), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n846), .B1(new_n851), .B2(new_n852), .ZN(G1337gat));
  NOR2_X1   g652(.A1(new_n830), .A2(new_n493), .ZN(new_n854));
  XNOR2_X1  g653(.A(KEYINPUT119), .B(G99gat), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n821), .A2(new_n724), .A3(new_n855), .ZN(new_n856));
  OAI22_X1  g655(.A1(new_n854), .A2(new_n855), .B1(new_n839), .B2(new_n856), .ZN(G1338gat));
  NOR3_X1   g656(.A1(new_n330), .A2(G106gat), .A3(new_n753), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n848), .A2(new_n849), .A3(new_n859), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n788), .A2(new_n494), .A3(new_n789), .A4(new_n829), .ZN(new_n861));
  XNOR2_X1  g660(.A(KEYINPUT120), .B(G106gat), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT53), .B1(new_n860), .B2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n866), .B1(new_n839), .B2(new_n859), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n861), .A2(KEYINPUT121), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n769), .A2(new_n869), .A3(new_n494), .A4(new_n829), .ZN(new_n870));
  AND3_X1   g669(.A1(new_n868), .A2(new_n870), .A3(new_n863), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n865), .B1(new_n867), .B2(new_n871), .ZN(G1339gat));
  INV_X1    g671(.A(KEYINPUT55), .ZN(new_n873));
  INV_X1    g672(.A(new_n709), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n701), .A2(new_n705), .A3(new_n707), .A4(new_n874), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n710), .A2(KEYINPUT54), .A3(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n708), .A2(new_n877), .A3(new_n709), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n722), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n873), .B1(new_n876), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n710), .A2(KEYINPUT54), .A3(new_n875), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n881), .A2(KEYINPUT55), .A3(new_n722), .A4(new_n878), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n880), .A2(new_n720), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n586), .B1(new_n598), .B2(new_n585), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n602), .A2(new_n603), .A3(new_n601), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI22_X1  g685(.A1(new_n615), .A2(new_n617), .B1(new_n612), .B2(new_n886), .ZN(new_n887));
  AOI22_X1  g686(.A1(new_n622), .A2(new_n883), .B1(new_n887), .B2(new_n724), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n888), .A2(new_n765), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n883), .A2(new_n887), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n890), .B1(new_n764), .B2(new_n763), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n696), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n698), .A2(new_n622), .A3(new_n724), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n895), .A2(new_n479), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n481), .A2(new_n330), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n544), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(G113gat), .B1(new_n900), .B2(new_n622), .ZN(new_n901));
  INV_X1    g700(.A(new_n894), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n892), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n330), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n475), .A2(new_n495), .A3(new_n821), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n770), .A2(new_n209), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n901), .B1(new_n906), .B2(new_n907), .ZN(G1340gat));
  NAND3_X1  g707(.A1(new_n900), .A2(new_n218), .A3(new_n724), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n904), .A2(new_n753), .A3(new_n905), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n910), .B2(new_n210), .ZN(new_n911));
  XOR2_X1   g710(.A(new_n911), .B(KEYINPUT122), .Z(G1341gat));
  NAND3_X1  g711(.A1(new_n900), .A2(new_n214), .A3(new_n697), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n904), .A2(new_n696), .A3(new_n905), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n913), .B1(new_n914), .B2(new_n214), .ZN(G1342gat));
  AOI21_X1  g714(.A(new_n207), .B1(new_n906), .B2(new_n765), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n900), .A2(new_n207), .A3(new_n765), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n916), .B1(new_n917), .B2(KEYINPUT56), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n918), .B1(KEYINPUT56), .B2(new_n917), .ZN(G1343gat));
  INV_X1    g718(.A(KEYINPUT123), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n920), .B1(new_n895), .B2(new_n479), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n493), .A2(new_n494), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n922), .A2(new_n544), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n924), .B1(KEYINPUT123), .B2(new_n896), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n925), .A2(new_n223), .A3(new_n622), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n493), .A2(new_n495), .A3(new_n475), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT57), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n928), .B1(new_n895), .B2(new_n330), .ZN(new_n929));
  OAI211_X1 g728(.A(KEYINPUT57), .B(new_n494), .C1(new_n893), .C2(new_n894), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n927), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n931), .A2(new_n622), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n926), .B1(new_n227), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(KEYINPUT58), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT58), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n926), .B(new_n935), .C1(new_n227), .C2(new_n932), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(G1344gat));
  NAND3_X1  g736(.A1(new_n925), .A2(new_n240), .A3(new_n724), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT59), .ZN(new_n939));
  OAI21_X1  g738(.A(KEYINPUT124), .B1(new_n889), .B2(new_n891), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n887), .B(new_n883), .C1(new_n659), .C2(new_n663), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT124), .ZN(new_n942));
  OAI211_X1 g741(.A(new_n941), .B(new_n942), .C1(new_n765), .C2(new_n888), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n940), .A2(new_n696), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(new_n902), .ZN(new_n945));
  AOI21_X1  g744(.A(KEYINPUT57), .B1(new_n945), .B2(new_n494), .ZN(new_n946));
  INV_X1    g745(.A(new_n930), .ZN(new_n947));
  OR2_X1    g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n927), .A2(new_n753), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n939), .B1(new_n950), .B2(G148gat), .ZN(new_n951));
  AOI211_X1 g750(.A(KEYINPUT59), .B(new_n240), .C1(new_n931), .C2(new_n724), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n938), .B1(new_n951), .B2(new_n952), .ZN(G1345gat));
  XOR2_X1   g752(.A(KEYINPUT82), .B(G155gat), .Z(new_n954));
  NAND3_X1  g753(.A1(new_n925), .A2(new_n697), .A3(new_n954), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n931), .A2(new_n697), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n955), .B1(new_n956), .B2(new_n954), .ZN(G1346gat));
  AOI21_X1  g756(.A(G162gat), .B1(new_n925), .B2(new_n765), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n664), .A2(new_n232), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n958), .B1(new_n931), .B2(new_n959), .ZN(G1347gat));
  NOR4_X1   g759(.A1(new_n895), .A2(new_n495), .A3(new_n897), .A4(new_n475), .ZN(new_n961));
  AOI21_X1  g760(.A(G169gat), .B1(new_n961), .B2(new_n622), .ZN(new_n962));
  NOR4_X1   g761(.A1(new_n904), .A2(new_n495), .A3(new_n475), .A4(new_n423), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n770), .A2(new_n352), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(G1348gat));
  NAND3_X1  g764(.A1(new_n961), .A2(new_n353), .A3(new_n724), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n963), .A2(new_n724), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n966), .B1(new_n967), .B2(new_n353), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n968), .B(KEYINPUT125), .ZN(G1349gat));
  NAND3_X1  g768(.A1(new_n961), .A2(new_n345), .A3(new_n697), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n963), .A2(new_n697), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n970), .B1(new_n971), .B2(new_n334), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g772(.A1(new_n961), .A2(new_n338), .A3(new_n765), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n963), .A2(new_n765), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(G190gat), .ZN(new_n976));
  AND2_X1   g775(.A1(new_n976), .A2(KEYINPUT61), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n976), .A2(KEYINPUT61), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n974), .B1(new_n977), .B2(new_n978), .ZN(G1351gat));
  OR3_X1    g778(.A1(new_n922), .A2(KEYINPUT126), .A3(new_n475), .ZN(new_n980));
  OAI21_X1  g779(.A(KEYINPUT126), .B1(new_n922), .B2(new_n475), .ZN(new_n981));
  AND4_X1   g780(.A1(new_n479), .A2(new_n980), .A3(new_n903), .A4(new_n981), .ZN(new_n982));
  AOI21_X1  g781(.A(G197gat), .B1(new_n982), .B2(new_n622), .ZN(new_n983));
  NOR3_X1   g782(.A1(new_n488), .A2(new_n475), .A3(new_n495), .ZN(new_n984));
  AND2_X1   g783(.A1(new_n948), .A2(new_n984), .ZN(new_n985));
  AND2_X1   g784(.A1(new_n622), .A2(G197gat), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n983), .B1(new_n985), .B2(new_n986), .ZN(G1352gat));
  INV_X1    g786(.A(G204gat), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n988), .B1(new_n985), .B2(new_n724), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n982), .A2(new_n988), .A3(new_n724), .ZN(new_n990));
  XNOR2_X1  g789(.A(new_n990), .B(KEYINPUT62), .ZN(new_n991));
  OR2_X1    g790(.A1(new_n989), .A2(new_n991), .ZN(G1353gat));
  NAND3_X1  g791(.A1(new_n982), .A2(new_n293), .A3(new_n697), .ZN(new_n993));
  OAI211_X1 g792(.A(new_n697), .B(new_n984), .C1(new_n946), .C2(new_n947), .ZN(new_n994));
  AND3_X1   g793(.A1(new_n994), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n995));
  AOI21_X1  g794(.A(KEYINPUT63), .B1(new_n994), .B2(G211gat), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n993), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT127), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI211_X1 g798(.A(KEYINPUT127), .B(new_n993), .C1(new_n995), .C2(new_n996), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n999), .A2(new_n1000), .ZN(G1354gat));
  NAND3_X1  g800(.A1(new_n982), .A2(new_n294), .A3(new_n765), .ZN(new_n1002));
  AND2_X1   g801(.A1(new_n985), .A2(new_n765), .ZN(new_n1003));
  OAI21_X1  g802(.A(new_n1002), .B1(new_n1003), .B2(new_n294), .ZN(G1355gat));
endmodule


