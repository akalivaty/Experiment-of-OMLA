

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XNOR2_X1 U321 ( .A(n289), .B(n332), .ZN(n375) );
  NOR2_X2 U322 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X2 U323 ( .A1(n478), .A2(n477), .ZN(n571) );
  NOR2_X1 U324 ( .A1(n463), .A2(n462), .ZN(n486) );
  XOR2_X1 U325 ( .A(n344), .B(n343), .Z(n578) );
  INV_X1 U326 ( .A(KEYINPUT124), .ZN(n439) );
  XNOR2_X1 U327 ( .A(KEYINPUT119), .B(KEYINPUT55), .ZN(n475) );
  XNOR2_X1 U328 ( .A(n309), .B(n308), .ZN(n546) );
  XOR2_X1 U329 ( .A(KEYINPUT69), .B(KEYINPUT13), .Z(n289) );
  AND2_X1 U330 ( .A1(G226GAT), .A2(G233GAT), .ZN(n290) );
  XOR2_X1 U331 ( .A(KEYINPUT110), .B(n377), .Z(n291) );
  XOR2_X1 U332 ( .A(G218GAT), .B(G162GAT), .Z(n292) );
  XNOR2_X1 U333 ( .A(n349), .B(n292), .ZN(n350) );
  XNOR2_X1 U334 ( .A(n351), .B(n350), .ZN(n355) );
  XNOR2_X1 U335 ( .A(n390), .B(n290), .ZN(n391) );
  XNOR2_X1 U336 ( .A(KEYINPUT36), .B(KEYINPUT98), .ZN(n359) );
  XNOR2_X1 U337 ( .A(KEYINPUT37), .B(KEYINPUT100), .ZN(n466) );
  XNOR2_X1 U338 ( .A(n392), .B(n391), .ZN(n394) );
  XNOR2_X1 U339 ( .A(n380), .B(n359), .ZN(n582) );
  XNOR2_X1 U340 ( .A(n476), .B(n475), .ZN(n478) );
  XNOR2_X1 U341 ( .A(n467), .B(n466), .ZN(n515) );
  XNOR2_X1 U342 ( .A(n403), .B(n402), .ZN(n518) );
  XNOR2_X1 U343 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U344 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U345 ( .A(n447), .B(n446), .ZN(G1352GAT) );
  XNOR2_X1 U346 ( .A(n472), .B(n471), .ZN(G1330GAT) );
  XOR2_X1 U347 ( .A(KEYINPUT126), .B(KEYINPUT125), .Z(n443) );
  XOR2_X1 U348 ( .A(G57GAT), .B(G85GAT), .Z(n294) );
  XNOR2_X1 U349 ( .A(G29GAT), .B(G148GAT), .ZN(n293) );
  XNOR2_X1 U350 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U351 ( .A(KEYINPUT6), .B(KEYINPUT85), .Z(n296) );
  XNOR2_X1 U352 ( .A(KEYINPUT4), .B(KEYINPUT5), .ZN(n295) );
  XNOR2_X1 U353 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U354 ( .A(n298), .B(n297), .ZN(n309) );
  XOR2_X1 U355 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n300) );
  XNOR2_X1 U356 ( .A(G141GAT), .B(G162GAT), .ZN(n299) );
  XNOR2_X1 U357 ( .A(n300), .B(n299), .ZN(n410) );
  XOR2_X1 U358 ( .A(G127GAT), .B(G155GAT), .Z(n336) );
  XOR2_X1 U359 ( .A(n410), .B(n336), .Z(n302) );
  NAND2_X1 U360 ( .A1(G225GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U361 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U362 ( .A(n303), .B(KEYINPUT1), .Z(n307) );
  XOR2_X1 U363 ( .A(G120GAT), .B(KEYINPUT0), .Z(n305) );
  XNOR2_X1 U364 ( .A(G113GAT), .B(G134GAT), .ZN(n304) );
  XNOR2_X1 U365 ( .A(n305), .B(n304), .ZN(n421) );
  XNOR2_X1 U366 ( .A(G1GAT), .B(n421), .ZN(n306) );
  XNOR2_X1 U367 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U368 ( .A(KEYINPUT54), .B(KEYINPUT118), .Z(n406) );
  INV_X1 U369 ( .A(KEYINPUT111), .ZN(n379) );
  XOR2_X1 U370 ( .A(G169GAT), .B(G8GAT), .Z(n399) );
  XNOR2_X1 U371 ( .A(G15GAT), .B(G22GAT), .ZN(n310) );
  XNOR2_X1 U372 ( .A(n310), .B(G1GAT), .ZN(n333) );
  XOR2_X1 U373 ( .A(n399), .B(n333), .Z(n312) );
  NAND2_X1 U374 ( .A1(G229GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U375 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U376 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n314) );
  XNOR2_X1 U377 ( .A(KEYINPUT67), .B(KEYINPUT64), .ZN(n313) );
  XNOR2_X1 U378 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U379 ( .A(n316), .B(n315), .Z(n326) );
  XOR2_X1 U380 ( .A(G43GAT), .B(G29GAT), .Z(n318) );
  XNOR2_X1 U381 ( .A(G50GAT), .B(KEYINPUT8), .ZN(n317) );
  XNOR2_X1 U382 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U383 ( .A(n319), .B(KEYINPUT65), .Z(n321) );
  XNOR2_X1 U384 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n320) );
  XNOR2_X1 U385 ( .A(n321), .B(n320), .ZN(n356) );
  XOR2_X1 U386 ( .A(KEYINPUT66), .B(G197GAT), .Z(n323) );
  XNOR2_X1 U387 ( .A(G113GAT), .B(G141GAT), .ZN(n322) );
  XNOR2_X1 U388 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U389 ( .A(n356), .B(n324), .ZN(n325) );
  XOR2_X1 U390 ( .A(n326), .B(n325), .Z(n547) );
  XOR2_X1 U391 ( .A(n547), .B(KEYINPUT68), .Z(n561) );
  XOR2_X1 U392 ( .A(KEYINPUT78), .B(KEYINPUT15), .Z(n328) );
  XNOR2_X1 U393 ( .A(KEYINPUT79), .B(KEYINPUT75), .ZN(n327) );
  XNOR2_X1 U394 ( .A(n328), .B(n327), .ZN(n344) );
  XOR2_X1 U395 ( .A(KEYINPUT76), .B(KEYINPUT14), .Z(n330) );
  NAND2_X1 U396 ( .A1(G231GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U397 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U398 ( .A(n331), .B(KEYINPUT12), .Z(n335) );
  XNOR2_X1 U399 ( .A(G71GAT), .B(G57GAT), .ZN(n332) );
  XNOR2_X1 U400 ( .A(n333), .B(n375), .ZN(n334) );
  XNOR2_X1 U401 ( .A(n335), .B(n334), .ZN(n340) );
  XOR2_X1 U402 ( .A(G183GAT), .B(G211GAT), .Z(n390) );
  XOR2_X1 U403 ( .A(G64GAT), .B(n390), .Z(n338) );
  XNOR2_X1 U404 ( .A(G78GAT), .B(n336), .ZN(n337) );
  XNOR2_X1 U405 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U406 ( .A(n340), .B(n339), .Z(n342) );
  XNOR2_X1 U407 ( .A(G8GAT), .B(KEYINPUT77), .ZN(n341) );
  XNOR2_X1 U408 ( .A(n342), .B(n341), .ZN(n343) );
  INV_X1 U409 ( .A(n578), .ZN(n554) );
  XOR2_X1 U410 ( .A(KEYINPUT72), .B(KEYINPUT71), .Z(n346) );
  XOR2_X1 U411 ( .A(G99GAT), .B(G85GAT), .Z(n371) );
  XOR2_X1 U412 ( .A(G190GAT), .B(KEYINPUT74), .Z(n395) );
  XNOR2_X1 U413 ( .A(n371), .B(n395), .ZN(n345) );
  XNOR2_X1 U414 ( .A(n346), .B(n345), .ZN(n351) );
  XOR2_X1 U415 ( .A(G92GAT), .B(KEYINPUT11), .Z(n348) );
  XNOR2_X1 U416 ( .A(G134GAT), .B(G106GAT), .ZN(n347) );
  XNOR2_X1 U417 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U418 ( .A(KEYINPUT10), .B(KEYINPUT73), .Z(n353) );
  NAND2_X1 U419 ( .A1(G232GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U420 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U421 ( .A(n355), .B(n354), .ZN(n358) );
  XNOR2_X1 U422 ( .A(n356), .B(KEYINPUT9), .ZN(n357) );
  XNOR2_X1 U423 ( .A(n358), .B(n357), .ZN(n380) );
  NOR2_X1 U424 ( .A1(n554), .A2(n582), .ZN(n361) );
  XNOR2_X1 U425 ( .A(KEYINPUT45), .B(KEYINPUT109), .ZN(n360) );
  XNOR2_X1 U426 ( .A(n361), .B(n360), .ZN(n376) );
  XOR2_X1 U427 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n363) );
  NAND2_X1 U428 ( .A1(G230GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U429 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U430 ( .A(n364), .B(KEYINPUT70), .Z(n369) );
  XOR2_X1 U431 ( .A(G78GAT), .B(G148GAT), .Z(n366) );
  XNOR2_X1 U432 ( .A(G106GAT), .B(G204GAT), .ZN(n365) );
  XNOR2_X1 U433 ( .A(n366), .B(n365), .ZN(n412) );
  XNOR2_X1 U434 ( .A(G176GAT), .B(G92GAT), .ZN(n367) );
  XNOR2_X1 U435 ( .A(n367), .B(G64GAT), .ZN(n396) );
  XNOR2_X1 U436 ( .A(n412), .B(n396), .ZN(n368) );
  XNOR2_X1 U437 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U438 ( .A(n370), .B(KEYINPUT33), .Z(n373) );
  XNOR2_X1 U439 ( .A(G120GAT), .B(n371), .ZN(n372) );
  XNOR2_X1 U440 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U441 ( .A(n375), .B(n374), .ZN(n448) );
  INV_X1 U442 ( .A(n448), .ZN(n574) );
  NOR2_X1 U443 ( .A1(n376), .A2(n574), .ZN(n377) );
  NOR2_X1 U444 ( .A1(n561), .A2(n291), .ZN(n378) );
  XNOR2_X1 U445 ( .A(n379), .B(n378), .ZN(n386) );
  INV_X1 U446 ( .A(n380), .ZN(n570) );
  INV_X1 U447 ( .A(n547), .ZN(n441) );
  XOR2_X1 U448 ( .A(KEYINPUT41), .B(n574), .Z(n549) );
  NAND2_X1 U449 ( .A1(n441), .A2(n549), .ZN(n381) );
  XNOR2_X1 U450 ( .A(KEYINPUT46), .B(n381), .ZN(n382) );
  XOR2_X1 U451 ( .A(KEYINPUT108), .B(n578), .Z(n565) );
  NAND2_X1 U452 ( .A1(n382), .A2(n565), .ZN(n383) );
  NOR2_X1 U453 ( .A1(n570), .A2(n383), .ZN(n384) );
  XOR2_X1 U454 ( .A(KEYINPUT47), .B(n384), .Z(n385) );
  NOR2_X1 U455 ( .A1(n386), .A2(n385), .ZN(n387) );
  XNOR2_X1 U456 ( .A(n387), .B(KEYINPUT48), .ZN(n527) );
  XOR2_X1 U457 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n389) );
  XNOR2_X1 U458 ( .A(KEYINPUT83), .B(KEYINPUT17), .ZN(n388) );
  XNOR2_X1 U459 ( .A(n389), .B(n388), .ZN(n426) );
  XOR2_X1 U460 ( .A(n426), .B(KEYINPUT86), .Z(n392) );
  XNOR2_X1 U461 ( .A(G36GAT), .B(G204GAT), .ZN(n393) );
  XNOR2_X1 U462 ( .A(n394), .B(n393), .ZN(n403) );
  XOR2_X1 U463 ( .A(n396), .B(n395), .Z(n401) );
  XOR2_X1 U464 ( .A(KEYINPUT84), .B(KEYINPUT21), .Z(n398) );
  XNOR2_X1 U465 ( .A(G197GAT), .B(G218GAT), .ZN(n397) );
  XNOR2_X1 U466 ( .A(n398), .B(n397), .ZN(n413) );
  XNOR2_X1 U467 ( .A(n399), .B(n413), .ZN(n400) );
  XOR2_X1 U468 ( .A(n401), .B(n400), .Z(n402) );
  INV_X1 U469 ( .A(n518), .ZN(n404) );
  NOR2_X1 U470 ( .A1(n527), .A2(n404), .ZN(n405) );
  XNOR2_X1 U471 ( .A(n406), .B(n405), .ZN(n407) );
  NOR2_X1 U472 ( .A1(n546), .A2(n407), .ZN(n474) );
  XOR2_X1 U473 ( .A(G155GAT), .B(KEYINPUT23), .Z(n409) );
  XNOR2_X1 U474 ( .A(G50GAT), .B(G22GAT), .ZN(n408) );
  XNOR2_X1 U475 ( .A(n409), .B(n408), .ZN(n411) );
  XOR2_X1 U476 ( .A(n411), .B(n410), .Z(n415) );
  XNOR2_X1 U477 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U478 ( .A(n415), .B(n414), .ZN(n420) );
  XOR2_X1 U479 ( .A(KEYINPUT22), .B(G211GAT), .Z(n417) );
  NAND2_X1 U480 ( .A1(G228GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U481 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U482 ( .A(KEYINPUT24), .B(n418), .Z(n419) );
  XNOR2_X1 U483 ( .A(n420), .B(n419), .ZN(n473) );
  XOR2_X1 U484 ( .A(n421), .B(G127GAT), .Z(n423) );
  NAND2_X1 U485 ( .A1(G227GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U486 ( .A(n423), .B(n422), .ZN(n437) );
  XOR2_X1 U487 ( .A(G190GAT), .B(G99GAT), .Z(n425) );
  XNOR2_X1 U488 ( .A(G43GAT), .B(KEYINPUT81), .ZN(n424) );
  XNOR2_X1 U489 ( .A(n425), .B(n424), .ZN(n427) );
  XOR2_X1 U490 ( .A(n427), .B(n426), .Z(n435) );
  XOR2_X1 U491 ( .A(G176GAT), .B(KEYINPUT20), .Z(n429) );
  XNOR2_X1 U492 ( .A(KEYINPUT80), .B(KEYINPUT82), .ZN(n428) );
  XNOR2_X1 U493 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U494 ( .A(G183GAT), .B(G71GAT), .Z(n431) );
  XNOR2_X1 U495 ( .A(G169GAT), .B(G15GAT), .ZN(n430) );
  XNOR2_X1 U496 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U497 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U498 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U499 ( .A(n437), .B(n436), .ZN(n530) );
  NOR2_X1 U500 ( .A1(n473), .A2(n530), .ZN(n438) );
  XNOR2_X1 U501 ( .A(n438), .B(KEYINPUT26), .ZN(n450) );
  NAND2_X1 U502 ( .A1(n474), .A2(n450), .ZN(n440) );
  XNOR2_X2 U503 ( .A(n440), .B(n439), .ZN(n580) );
  NAND2_X1 U504 ( .A1(n580), .A2(n441), .ZN(n442) );
  XNOR2_X1 U505 ( .A(n443), .B(n442), .ZN(n447) );
  XNOR2_X1 U506 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n445) );
  INV_X1 U507 ( .A(KEYINPUT59), .ZN(n444) );
  NAND2_X1 U508 ( .A1(n561), .A2(n448), .ZN(n488) );
  XNOR2_X1 U509 ( .A(KEYINPUT27), .B(KEYINPUT87), .ZN(n449) );
  XOR2_X1 U510 ( .A(n449), .B(n518), .Z(n458) );
  NAND2_X1 U511 ( .A1(n450), .A2(n458), .ZN(n543) );
  XNOR2_X1 U512 ( .A(n543), .B(KEYINPUT89), .ZN(n455) );
  NAND2_X1 U513 ( .A1(n530), .A2(n518), .ZN(n451) );
  NAND2_X1 U514 ( .A1(n451), .A2(n473), .ZN(n452) );
  XNOR2_X1 U515 ( .A(n452), .B(KEYINPUT90), .ZN(n453) );
  XNOR2_X1 U516 ( .A(KEYINPUT25), .B(n453), .ZN(n454) );
  NOR2_X1 U517 ( .A1(n455), .A2(n454), .ZN(n456) );
  NOR2_X1 U518 ( .A1(n546), .A2(n456), .ZN(n457) );
  XOR2_X1 U519 ( .A(KEYINPUT91), .B(n457), .Z(n463) );
  INV_X1 U520 ( .A(n458), .ZN(n459) );
  XOR2_X1 U521 ( .A(KEYINPUT28), .B(n473), .Z(n524) );
  NOR2_X1 U522 ( .A1(n459), .A2(n524), .ZN(n460) );
  NAND2_X1 U523 ( .A1(n546), .A2(n460), .ZN(n528) );
  NOR2_X1 U524 ( .A1(n530), .A2(n528), .ZN(n461) );
  XNOR2_X1 U525 ( .A(KEYINPUT88), .B(n461), .ZN(n462) );
  NOR2_X1 U526 ( .A1(n578), .A2(n486), .ZN(n464) );
  XNOR2_X1 U527 ( .A(n464), .B(KEYINPUT99), .ZN(n465) );
  NOR2_X1 U528 ( .A1(n582), .A2(n465), .ZN(n467) );
  NOR2_X1 U529 ( .A1(n488), .A2(n515), .ZN(n468) );
  XNOR2_X1 U530 ( .A(n468), .B(KEYINPUT38), .ZN(n504) );
  NAND2_X1 U531 ( .A1(n504), .A2(n530), .ZN(n472) );
  XOR2_X1 U532 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n470) );
  XNOR2_X1 U533 ( .A(G43GAT), .B(KEYINPUT104), .ZN(n469) );
  NAND2_X1 U534 ( .A1(n474), .A2(n473), .ZN(n476) );
  INV_X1 U535 ( .A(n530), .ZN(n477) );
  NAND2_X1 U536 ( .A1(n571), .A2(n549), .ZN(n481) );
  XOR2_X1 U537 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n479) );
  XNOR2_X1 U538 ( .A(n479), .B(G176GAT), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n481), .B(n480), .ZN(G1349GAT) );
  XNOR2_X1 U540 ( .A(G1GAT), .B(KEYINPUT94), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n482), .B(KEYINPUT34), .ZN(n483) );
  XOR2_X1 U542 ( .A(KEYINPUT93), .B(n483), .Z(n490) );
  NOR2_X1 U543 ( .A1(n570), .A2(n554), .ZN(n484) );
  XOR2_X1 U544 ( .A(KEYINPUT16), .B(n484), .Z(n485) );
  NOR2_X1 U545 ( .A1(n486), .A2(n485), .ZN(n487) );
  XOR2_X1 U546 ( .A(KEYINPUT92), .B(n487), .Z(n506) );
  NOR2_X1 U547 ( .A1(n506), .A2(n488), .ZN(n496) );
  NAND2_X1 U548 ( .A1(n496), .A2(n546), .ZN(n489) );
  XNOR2_X1 U549 ( .A(n490), .B(n489), .ZN(G1324GAT) );
  XOR2_X1 U550 ( .A(G8GAT), .B(KEYINPUT95), .Z(n492) );
  NAND2_X1 U551 ( .A1(n496), .A2(n518), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n492), .B(n491), .ZN(G1325GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT96), .B(KEYINPUT35), .Z(n494) );
  NAND2_X1 U554 ( .A1(n496), .A2(n530), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U556 ( .A(G15GAT), .B(n495), .ZN(G1326GAT) );
  XOR2_X1 U557 ( .A(G22GAT), .B(KEYINPUT97), .Z(n498) );
  NAND2_X1 U558 ( .A1(n496), .A2(n524), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n498), .B(n497), .ZN(G1327GAT) );
  NAND2_X1 U560 ( .A1(n504), .A2(n546), .ZN(n501) );
  XNOR2_X1 U561 ( .A(G29GAT), .B(KEYINPUT101), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n499), .B(KEYINPUT39), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n501), .B(n500), .ZN(G1328GAT) );
  NAND2_X1 U564 ( .A1(n504), .A2(n518), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n502), .B(KEYINPUT102), .ZN(n503) );
  XNOR2_X1 U566 ( .A(G36GAT), .B(n503), .ZN(G1329GAT) );
  NAND2_X1 U567 ( .A1(n504), .A2(n524), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n505), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n508) );
  NAND2_X1 U570 ( .A1(n549), .A2(n547), .ZN(n514) );
  NOR2_X1 U571 ( .A1(n506), .A2(n514), .ZN(n511) );
  NAND2_X1 U572 ( .A1(n546), .A2(n511), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n508), .B(n507), .ZN(G1332GAT) );
  NAND2_X1 U574 ( .A1(n511), .A2(n518), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n509), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U576 ( .A1(n530), .A2(n511), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n510), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U578 ( .A(G78GAT), .B(KEYINPUT43), .Z(n513) );
  NAND2_X1 U579 ( .A1(n511), .A2(n524), .ZN(n512) );
  XNOR2_X1 U580 ( .A(n513), .B(n512), .ZN(G1335GAT) );
  XOR2_X1 U581 ( .A(G85GAT), .B(KEYINPUT105), .Z(n517) );
  NOR2_X1 U582 ( .A1(n515), .A2(n514), .ZN(n523) );
  NAND2_X1 U583 ( .A1(n523), .A2(n546), .ZN(n516) );
  XNOR2_X1 U584 ( .A(n517), .B(n516), .ZN(G1336GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n520) );
  NAND2_X1 U586 ( .A1(n523), .A2(n518), .ZN(n519) );
  XNOR2_X1 U587 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U588 ( .A(G92GAT), .B(n521), .ZN(G1337GAT) );
  NAND2_X1 U589 ( .A1(n530), .A2(n523), .ZN(n522) );
  XNOR2_X1 U590 ( .A(n522), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U591 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n525), .B(KEYINPUT44), .ZN(n526) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(n526), .ZN(G1339GAT) );
  BUF_X1 U594 ( .A(n527), .Z(n544) );
  NOR2_X1 U595 ( .A1(n544), .A2(n528), .ZN(n529) );
  NAND2_X1 U596 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U597 ( .A(KEYINPUT112), .B(n531), .ZN(n536) );
  INV_X1 U598 ( .A(n536), .ZN(n539) );
  NAND2_X1 U599 ( .A1(n539), .A2(n561), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n532), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT113), .B(KEYINPUT49), .Z(n534) );
  NAND2_X1 U602 ( .A1(n549), .A2(n539), .ZN(n533) );
  XNOR2_X1 U603 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U604 ( .A(G120GAT), .B(n535), .Z(G1341GAT) );
  NOR2_X1 U605 ( .A1(n565), .A2(n536), .ZN(n537) );
  XOR2_X1 U606 ( .A(KEYINPUT50), .B(n537), .Z(n538) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n541) );
  NAND2_X1 U609 ( .A1(n570), .A2(n539), .ZN(n540) );
  XNOR2_X1 U610 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U611 ( .A(G134GAT), .B(n542), .ZN(G1343GAT) );
  NOR2_X1 U612 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U613 ( .A1(n546), .A2(n545), .ZN(n558) );
  NOR2_X1 U614 ( .A1(n547), .A2(n558), .ZN(n548) );
  XOR2_X1 U615 ( .A(G141GAT), .B(n548), .Z(G1344GAT) );
  INV_X1 U616 ( .A(n549), .ZN(n550) );
  NOR2_X1 U617 ( .A1(n550), .A2(n558), .ZN(n552) );
  XNOR2_X1 U618 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(n553), .ZN(G1345GAT) );
  NOR2_X1 U621 ( .A1(n554), .A2(n558), .ZN(n556) );
  XNOR2_X1 U622 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U624 ( .A(G155GAT), .B(n557), .ZN(G1346GAT) );
  NOR2_X1 U625 ( .A1(n380), .A2(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G162GAT), .B(KEYINPUT117), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1347GAT) );
  NAND2_X1 U628 ( .A1(n571), .A2(n561), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(KEYINPUT120), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(G169GAT), .ZN(G1348GAT) );
  INV_X1 U631 ( .A(n571), .ZN(n564) );
  NOR2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U633 ( .A(G183GAT), .B(n566), .Z(G1350GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n568) );
  XNOR2_X1 U635 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n567) );
  XNOR2_X1 U636 ( .A(n568), .B(n567), .ZN(n569) );
  XOR2_X1 U637 ( .A(KEYINPUT121), .B(n569), .Z(n573) );
  NAND2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1351GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n576) );
  NAND2_X1 U641 ( .A1(n574), .A2(n580), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XOR2_X1 U643 ( .A(G204GAT), .B(n577), .Z(G1353GAT) );
  NAND2_X1 U644 ( .A1(n578), .A2(n580), .ZN(n579) );
  XNOR2_X1 U645 ( .A(G211GAT), .B(n579), .ZN(G1354GAT) );
  INV_X1 U646 ( .A(n580), .ZN(n581) );
  XOR2_X1 U647 ( .A(KEYINPUT62), .B(n583), .Z(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

