//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 1 0 0 1 0 1 0 0 1 1 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n777, new_n778,
    new_n779, new_n781, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n989, new_n990;
  XOR2_X1   g000(.A(KEYINPUT31), .B(G50gat), .Z(new_n202));
  XNOR2_X1  g001(.A(G155gat), .B(G162gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  OR2_X1    g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206));
  AND2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT2), .ZN(new_n209));
  NAND4_X1  g008(.A1(new_n204), .A2(new_n207), .A3(KEYINPUT76), .A4(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT76), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n203), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G155gat), .ZN(new_n213));
  INV_X1    g012(.A(G162gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n215), .A2(KEYINPUT76), .A3(new_n208), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n209), .A2(new_n205), .A3(new_n206), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n212), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n210), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT3), .ZN(new_n220));
  AOI21_X1  g019(.A(KEYINPUT29), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  XOR2_X1   g020(.A(G197gat), .B(G204gat), .Z(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G211gat), .B(G218gat), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT72), .B(G211gat), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n225), .A2(G218gat), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n223), .B(new_n224), .C1(new_n226), .C2(KEYINPUT22), .ZN(new_n227));
  INV_X1    g026(.A(new_n224), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT22), .B1(new_n225), .B2(G218gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n228), .B1(new_n229), .B2(new_n222), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n221), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT29), .B1(new_n227), .B2(new_n230), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n210), .B(new_n218), .C1(new_n234), .C2(KEYINPUT3), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT81), .ZN(new_n236));
  NAND2_X1  g035(.A1(G228gat), .A2(G233gat), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n233), .A2(new_n235), .A3(new_n236), .A4(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT29), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n231), .A2(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n219), .B1(new_n241), .B2(new_n220), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n238), .B1(new_n221), .B2(new_n231), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT81), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n239), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT80), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n232), .B1(new_n235), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n242), .A2(KEYINPUT80), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n238), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n202), .B1(new_n245), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n202), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n239), .A2(new_n244), .ZN(new_n252));
  AND2_X1   g051(.A1(new_n247), .A2(new_n248), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n251), .B(new_n252), .C1(new_n253), .C2(new_n238), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(G78gat), .B(G106gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(G22gat), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n250), .A2(new_n254), .A3(new_n257), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  XOR2_X1   g060(.A(G183gat), .B(G190gat), .Z(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT24), .ZN(new_n263));
  NOR2_X1   g062(.A1(G169gat), .A2(G176gat), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT23), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(G183gat), .A2(G190gat), .ZN(new_n267));
  INV_X1    g066(.A(G169gat), .ZN(new_n268));
  INV_X1    g067(.A(G176gat), .ZN(new_n269));
  OAI22_X1  g068(.A1(new_n267), .A2(KEYINPUT24), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n263), .A2(new_n266), .A3(KEYINPUT25), .A4(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT64), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n263), .A2(new_n266), .A3(new_n271), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT25), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n270), .B1(new_n262), .B2(KEYINPUT24), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n278), .A2(KEYINPUT64), .A3(KEYINPUT25), .A4(new_n266), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n274), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n268), .A2(new_n269), .ZN(new_n281));
  NOR3_X1   g080(.A1(new_n281), .A2(KEYINPUT26), .A3(new_n264), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n264), .A2(KEYINPUT26), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(new_n267), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  XOR2_X1   g084(.A(KEYINPUT27), .B(G183gat), .Z(new_n286));
  INV_X1    g085(.A(KEYINPUT65), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(G183gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT27), .ZN(new_n290));
  AOI21_X1  g089(.A(G190gat), .B1(new_n290), .B2(KEYINPUT65), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT28), .B1(new_n288), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT28), .ZN(new_n293));
  NOR3_X1   g092(.A1(new_n286), .A2(new_n293), .A3(G190gat), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n285), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT67), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G113gat), .ZN(new_n299));
  INV_X1    g098(.A(G120gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT1), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n302), .B1(G113gat), .B2(G120gat), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT66), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G127gat), .B(G134gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n305), .B(KEYINPUT66), .C1(new_n301), .C2(new_n303), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n280), .A2(KEYINPUT67), .A3(new_n295), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n298), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n309), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n280), .A2(KEYINPUT67), .A3(new_n312), .A4(new_n295), .ZN(new_n313));
  AND2_X1   g112(.A1(G227gat), .A2(G233gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n311), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT32), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT33), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  XOR2_X1   g117(.A(KEYINPUT68), .B(G71gat), .Z(new_n319));
  XNOR2_X1  g118(.A(new_n319), .B(G99gat), .ZN(new_n320));
  XOR2_X1   g119(.A(G15gat), .B(G43gat), .Z(new_n321));
  XOR2_X1   g120(.A(new_n320), .B(new_n321), .Z(new_n322));
  NAND3_X1  g121(.A1(new_n316), .A2(new_n318), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n322), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n315), .B(KEYINPUT32), .C1(new_n317), .C2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT69), .ZN(new_n327));
  AND2_X1   g126(.A1(new_n311), .A2(new_n313), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n327), .B(KEYINPUT34), .C1(new_n328), .C2(new_n314), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT34), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n314), .B1(new_n311), .B2(new_n313), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n330), .B1(new_n331), .B2(KEYINPUT69), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n326), .A2(new_n333), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n261), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n296), .A2(new_n240), .ZN(new_n336));
  NAND2_X1  g135(.A1(G226gat), .A2(G233gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n337), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT73), .B1(new_n296), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT73), .ZN(new_n341));
  AOI211_X1 g140(.A(new_n341), .B(new_n337), .C1(new_n280), .C2(new_n295), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n338), .B(new_n231), .C1(new_n340), .C2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n296), .A2(new_n339), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT29), .B1(new_n280), .B2(new_n295), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n344), .B1(new_n339), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n231), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT74), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT74), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n343), .A2(new_n351), .A3(new_n348), .ZN(new_n352));
  XNOR2_X1  g151(.A(G8gat), .B(G36gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n353), .B(KEYINPUT75), .ZN(new_n354));
  XNOR2_X1  g153(.A(G64gat), .B(G92gat), .ZN(new_n355));
  XOR2_X1   g154(.A(new_n354), .B(new_n355), .Z(new_n356));
  NAND3_X1  g155(.A1(new_n350), .A2(new_n352), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n356), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n343), .A2(new_n348), .A3(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT30), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OR2_X1    g160(.A1(new_n359), .A2(new_n360), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n357), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n219), .A2(new_n220), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n210), .A2(new_n218), .A3(KEYINPUT3), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n364), .A2(new_n312), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(G225gat), .A2(G233gat), .ZN(new_n367));
  AND2_X1   g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  XOR2_X1   g167(.A(KEYINPUT77), .B(KEYINPUT5), .Z(new_n369));
  NAND2_X1  g168(.A1(new_n219), .A2(new_n309), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT78), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n370), .A2(new_n371), .A3(KEYINPUT4), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(KEYINPUT4), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT4), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n219), .A2(new_n374), .A3(new_n309), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(KEYINPUT78), .A3(new_n375), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n368), .A2(new_n369), .A3(new_n372), .A4(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G1gat), .B(G29gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n378), .B(KEYINPUT0), .ZN(new_n379));
  XNOR2_X1  g178(.A(G57gat), .B(G85gat), .ZN(new_n380));
  XOR2_X1   g179(.A(new_n379), .B(new_n380), .Z(new_n381));
  NAND4_X1  g180(.A1(new_n210), .A2(new_n218), .A3(new_n308), .A4(new_n307), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n370), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n367), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n369), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n373), .A2(new_n375), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n366), .A2(new_n367), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n377), .A2(new_n381), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT79), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n377), .A2(new_n388), .ZN(new_n392));
  INV_X1    g191(.A(new_n381), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT6), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n377), .A2(new_n388), .A3(KEYINPUT79), .A4(new_n381), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n391), .A2(new_n394), .A3(new_n395), .A4(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n381), .B1(new_n377), .B2(new_n388), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT6), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n363), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n326), .A2(new_n333), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT70), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT70), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n326), .A2(new_n333), .A3(new_n405), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n335), .A2(new_n402), .A3(new_n404), .A4(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT35), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n323), .A2(new_n329), .A3(new_n332), .A4(new_n325), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n403), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n410), .A2(new_n261), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT35), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n411), .A2(new_n412), .A3(new_n402), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n408), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n397), .A2(new_n399), .A3(new_n359), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT37), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n416), .B1(new_n346), .B2(new_n231), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n338), .B(new_n347), .C1(new_n340), .C2(new_n342), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT38), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n343), .A2(new_n416), .A3(new_n348), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n419), .A2(new_n356), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT85), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n419), .A2(KEYINPUT85), .A3(new_n356), .A4(new_n420), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n415), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n350), .A2(KEYINPUT37), .A3(new_n352), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n420), .A2(new_n356), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT38), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n261), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n376), .A2(new_n366), .A3(new_n372), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n384), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT39), .ZN(new_n432));
  INV_X1    g231(.A(new_n383), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n432), .B1(new_n433), .B2(new_n367), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n430), .A2(new_n432), .A3(new_n384), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n436), .A2(KEYINPUT83), .A3(new_n381), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT83), .B1(new_n436), .B2(new_n381), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n435), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT40), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n394), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n436), .A2(new_n381), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT83), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI22_X1  g244(.A1(new_n445), .A2(new_n437), .B1(new_n431), .B2(new_n434), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n446), .A2(KEYINPUT40), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n442), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT84), .B1(new_n448), .B2(new_n363), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n398), .B1(new_n446), .B2(KEYINPUT40), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n440), .A2(new_n441), .ZN(new_n451));
  AND4_X1   g250(.A1(KEYINPUT84), .A2(new_n363), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n429), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  AND3_X1   g252(.A1(new_n250), .A2(new_n254), .A3(new_n257), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n257), .B1(new_n250), .B2(new_n254), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n357), .A2(new_n361), .A3(new_n362), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n456), .B1(new_n457), .B2(new_n400), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n409), .A2(KEYINPUT36), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n459), .A2(new_n404), .A3(new_n406), .ZN(new_n460));
  XOR2_X1   g259(.A(KEYINPUT71), .B(KEYINPUT36), .Z(new_n461));
  NAND2_X1  g260(.A1(new_n410), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n458), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT82), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n453), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n326), .A2(new_n405), .A3(new_n333), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n405), .B1(new_n326), .B2(new_n333), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI22_X1  g267(.A1(new_n468), .A2(new_n459), .B1(new_n410), .B2(new_n461), .ZN(new_n469));
  NOR3_X1   g268(.A1(new_n469), .A2(KEYINPUT82), .A3(new_n458), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n414), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  XOR2_X1   g270(.A(KEYINPUT93), .B(KEYINPUT18), .Z(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(G22gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(G15gat), .ZN(new_n475));
  INV_X1    g274(.A(G15gat), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(G22gat), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT91), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n475), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(G8gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(G15gat), .B(G22gat), .ZN(new_n481));
  INV_X1    g280(.A(G8gat), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n481), .A2(new_n478), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT16), .ZN(new_n485));
  AOI21_X1  g284(.A(G1gat), .B1(new_n481), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n486), .A2(new_n480), .A3(new_n483), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AND2_X1   g289(.A1(G43gat), .A2(G50gat), .ZN(new_n491));
  OR2_X1    g290(.A1(KEYINPUT88), .A2(KEYINPUT15), .ZN(new_n492));
  NAND2_X1  g291(.A1(KEYINPUT88), .A2(KEYINPUT15), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(G43gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT89), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT89), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(G43gat), .ZN(new_n498));
  INV_X1    g297(.A(G50gat), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n496), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(G29gat), .A2(G36gat), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G43gat), .B(G50gat), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n503), .B1(new_n504), .B2(KEYINPUT15), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT14), .ZN(new_n507));
  INV_X1    g306(.A(G29gat), .ZN(new_n508));
  INV_X1    g307(.A(G36gat), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT90), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT90), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n512), .A2(new_n507), .A3(new_n508), .A4(new_n509), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n511), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n510), .A2(new_n514), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n502), .ZN(new_n517));
  NOR2_X1   g316(.A1(G43gat), .A2(G50gat), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT15), .B1(new_n491), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n517), .A2(KEYINPUT87), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT87), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n503), .B1(new_n510), .B2(new_n514), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n522), .B1(new_n523), .B2(new_n519), .ZN(new_n524));
  AOI22_X1  g323(.A1(new_n506), .A2(new_n515), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n490), .B1(new_n525), .B2(KEYINPUT17), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n515), .A2(new_n501), .A3(new_n505), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT87), .B1(new_n517), .B2(new_n520), .ZN(new_n528));
  NOR3_X1   g327(.A1(new_n523), .A2(new_n522), .A3(new_n519), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n527), .B(KEYINPUT17), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT92), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n521), .A2(new_n524), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n533), .A2(KEYINPUT92), .A3(KEYINPUT17), .A4(new_n527), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n526), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(G229gat), .A2(G233gat), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n536), .B1(new_n525), .B2(new_n490), .ZN(new_n537));
  OAI211_X1 g336(.A(KEYINPUT94), .B(new_n473), .C1(new_n535), .C2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT94), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n532), .A2(new_n534), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n486), .A2(new_n480), .A3(new_n483), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n481), .A2(new_n485), .ZN(new_n542));
  INV_X1    g341(.A(G1gat), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n480), .A2(new_n483), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n537), .B1(new_n540), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n539), .B1(new_n549), .B2(new_n472), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n545), .A2(new_n547), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n533), .B(new_n527), .C1(new_n541), .C2(new_n544), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n551), .A2(new_n552), .A3(KEYINPUT95), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT95), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n525), .A2(new_n554), .A3(new_n490), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  XOR2_X1   g355(.A(new_n536), .B(KEYINPUT13), .Z(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n549), .A2(KEYINPUT18), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n538), .A2(new_n550), .A3(new_n558), .A4(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(G113gat), .B(G141gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G169gat), .B(G197gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT12), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n560), .A2(new_n567), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n557), .A2(new_n556), .B1(new_n549), .B2(KEYINPUT18), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT96), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n570), .B(new_n473), .C1(new_n535), .C2(new_n537), .ZN(new_n571));
  OAI21_X1  g370(.A(KEYINPUT96), .B1(new_n549), .B2(new_n472), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n569), .A2(new_n566), .A3(new_n571), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n471), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(G71gat), .ZN(new_n576));
  INV_X1    g375(.A(G78gat), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(G71gat), .A2(G78gat), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT9), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G57gat), .B(G64gat), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT97), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(G57gat), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n586), .A2(G64gat), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n586), .A2(G64gat), .ZN(new_n588));
  NOR3_X1   g387(.A1(new_n587), .A2(new_n588), .A3(KEYINPUT97), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n580), .B1(new_n585), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT99), .ZN(new_n591));
  NAND2_X1  g390(.A1(KEYINPUT98), .A2(G64gat), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(KEYINPUT98), .A2(G64gat), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n591), .B(G57gat), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n579), .B1(new_n578), .B2(new_n581), .ZN(new_n596));
  INV_X1    g395(.A(new_n594), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n586), .B1(new_n597), .B2(new_n592), .ZN(new_n598));
  INV_X1    g397(.A(G64gat), .ZN(new_n599));
  OAI21_X1  g398(.A(KEYINPUT99), .B1(new_n599), .B2(G57gat), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n595), .B(new_n596), .C1(new_n598), .C2(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(KEYINPUT21), .B1(new_n590), .B2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT100), .ZN(new_n603));
  XNOR2_X1  g402(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT101), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n603), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G183gat), .B(G211gat), .ZN(new_n607));
  OR2_X1    g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n590), .A2(new_n601), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT21), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n490), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G127gat), .B(G155gat), .ZN(new_n614));
  NAND2_X1  g413(.A1(G231gat), .A2(G233gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n613), .B(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n610), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n608), .A2(new_n617), .A3(new_n609), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AND2_X1   g420(.A1(G232gat), .A2(G233gat), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n622), .A2(KEYINPUT41), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT102), .ZN(new_n624));
  XNOR2_X1  g423(.A(G134gat), .B(G162gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(G85gat), .A2(G92gat), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(KEYINPUT7), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT7), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n630), .A2(G85gat), .A3(G92gat), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(G99gat), .A2(G106gat), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(G99gat), .A2(G106gat), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(G85gat), .ZN(new_n637));
  INV_X1    g436(.A(G92gat), .ZN(new_n638));
  AOI22_X1  g437(.A1(KEYINPUT8), .A2(new_n633), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AND3_X1   g438(.A1(new_n632), .A2(new_n636), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n636), .B1(new_n632), .B2(new_n639), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  OAI211_X1 g441(.A(new_n540), .B(new_n642), .C1(KEYINPUT17), .C2(new_n525), .ZN(new_n643));
  XOR2_X1   g442(.A(G190gat), .B(G218gat), .Z(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n632), .A2(new_n639), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n646), .B1(new_n634), .B2(new_n635), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n632), .A2(new_n636), .A3(new_n639), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI22_X1  g448(.A1(new_n547), .A2(new_n649), .B1(KEYINPUT41), .B2(new_n622), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n643), .A2(new_n645), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n645), .B1(new_n643), .B2(new_n650), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n627), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n653), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n655), .A2(new_n626), .A3(new_n651), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT105), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n646), .A2(KEYINPUT103), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n590), .A2(new_n601), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(new_n649), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n642), .A2(new_n601), .A3(new_n590), .A4(new_n659), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT10), .ZN(new_n664));
  OAI21_X1  g463(.A(KEYINPUT10), .B1(new_n640), .B2(new_n641), .ZN(new_n665));
  OAI21_X1  g464(.A(KEYINPUT104), .B1(new_n611), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n664), .B1(new_n647), .B2(new_n648), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT104), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n667), .A2(new_n668), .A3(new_n601), .A4(new_n590), .ZN(new_n669));
  AOI22_X1  g468(.A1(new_n663), .A2(new_n664), .B1(new_n666), .B2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(G230gat), .ZN(new_n671));
  INV_X1    g470(.A(G233gat), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n658), .B1(new_n670), .B2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n673), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n669), .A2(new_n666), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(KEYINPUT10), .B1(new_n661), .B2(new_n662), .ZN(new_n678));
  OAI211_X1 g477(.A(KEYINPUT105), .B(new_n675), .C1(new_n677), .C2(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n663), .A2(new_n675), .ZN(new_n680));
  XNOR2_X1  g479(.A(G120gat), .B(G148gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(G176gat), .B(G204gat), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n681), .B(new_n682), .Z(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n674), .A2(new_n679), .A3(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n678), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n673), .B1(new_n687), .B2(new_n676), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n684), .B1(new_n688), .B2(new_n680), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n621), .A2(new_n657), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n575), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n400), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(new_n543), .ZN(G1324gat));
  XOR2_X1   g493(.A(KEYINPUT16), .B(G8gat), .Z(new_n695));
  NAND4_X1  g494(.A1(new_n575), .A2(new_n363), .A3(new_n691), .A4(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT42), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(G8gat), .B1(new_n692), .B2(new_n457), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n699), .A2(new_n696), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n698), .B1(new_n700), .B2(new_n697), .ZN(G1325gat));
  NAND2_X1  g500(.A1(new_n460), .A2(new_n462), .ZN(new_n702));
  OAI21_X1  g501(.A(G15gat), .B1(new_n692), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n410), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(new_n476), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n703), .B1(new_n692), .B2(new_n705), .ZN(G1326gat));
  NOR2_X1   g505(.A1(new_n692), .A2(new_n456), .ZN(new_n707));
  XOR2_X1   g506(.A(KEYINPUT43), .B(G22gat), .Z(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(G1327gat));
  INV_X1    g508(.A(new_n690), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n621), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n657), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n575), .A2(new_n713), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n714), .A2(G29gat), .A3(new_n400), .ZN(new_n715));
  OR2_X1    g514(.A1(new_n715), .A2(KEYINPUT45), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(KEYINPUT45), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n453), .A2(new_n463), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n414), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n657), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n712), .A2(new_n718), .ZN(new_n722));
  AOI22_X1  g521(.A1(new_n718), .A2(new_n721), .B1(new_n471), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n574), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n711), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(G29gat), .B1(new_n726), .B2(new_n400), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n716), .A2(new_n717), .A3(new_n727), .ZN(G1328gat));
  NOR3_X1   g527(.A1(new_n714), .A2(G36gat), .A3(new_n457), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT46), .ZN(new_n730));
  OR2_X1    g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(G36gat), .B1(new_n726), .B2(new_n457), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n729), .A2(new_n730), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(G1329gat));
  INV_X1    g533(.A(KEYINPUT106), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT47), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n575), .A2(new_n704), .A3(new_n713), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n496), .A2(new_n498), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n735), .A2(new_n736), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n702), .A2(new_n739), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n723), .A2(new_n725), .A3(new_n742), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n740), .A2(new_n741), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n741), .B1(new_n740), .B2(new_n743), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n744), .A2(new_n745), .ZN(G1330gat));
  NOR2_X1   g545(.A1(new_n456), .A2(G50gat), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n575), .A2(new_n713), .A3(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT107), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT48), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n471), .A2(new_n722), .ZN(new_n752));
  AOI22_X1  g551(.A1(new_n463), .A2(new_n453), .B1(new_n408), .B2(new_n413), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n718), .B1(new_n753), .B2(new_n712), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n752), .A2(new_n261), .A3(new_n754), .A4(new_n725), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n499), .A2(KEYINPUT48), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n751), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n723), .A2(KEYINPUT108), .A3(new_n261), .A4(new_n725), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT108), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n755), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n758), .A2(new_n760), .A3(G50gat), .ZN(new_n761));
  OR2_X1    g560(.A1(new_n748), .A2(KEYINPUT107), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n757), .B1(new_n763), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g563(.A1(new_n621), .A2(new_n657), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n765), .A2(new_n724), .A3(new_n690), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT109), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n720), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n768), .A2(new_n400), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(new_n586), .ZN(G1332gat));
  INV_X1    g569(.A(new_n768), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n457), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(KEYINPUT110), .ZN(new_n774));
  OR2_X1    g573(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n774), .B(new_n775), .ZN(G1333gat));
  OAI21_X1  g575(.A(G71gat), .B1(new_n768), .B2(new_n702), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n704), .A2(new_n576), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n768), .B2(new_n778), .ZN(new_n779));
  XOR2_X1   g578(.A(new_n779), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g579(.A1(new_n768), .A2(new_n456), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(new_n577), .ZN(G1335gat));
  INV_X1    g581(.A(new_n621), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n783), .A2(new_n574), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n690), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(KEYINPUT111), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n723), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(G85gat), .B1(new_n787), .B2(new_n400), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n712), .B1(new_n719), .B2(new_n414), .ZN(new_n789));
  AND3_X1   g588(.A1(new_n789), .A2(KEYINPUT51), .A3(new_n784), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT51), .B1(new_n789), .B2(new_n784), .ZN(new_n791));
  OR2_X1    g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n401), .A2(new_n637), .A3(new_n690), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n788), .B1(new_n793), .B2(new_n794), .ZN(G1336gat));
  NAND4_X1  g594(.A1(new_n752), .A2(new_n363), .A3(new_n754), .A4(new_n786), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(G92gat), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n457), .A2(G92gat), .A3(new_n710), .ZN(new_n798));
  XOR2_X1   g597(.A(new_n798), .B(KEYINPUT112), .Z(new_n799));
  OAI21_X1  g598(.A(new_n799), .B1(new_n790), .B2(new_n791), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n797), .A2(KEYINPUT52), .A3(new_n800), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n723), .A2(KEYINPUT113), .A3(new_n363), .A4(new_n786), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n796), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n802), .A2(new_n804), .A3(G92gat), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n792), .A2(new_n798), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n801), .B1(new_n807), .B2(new_n808), .ZN(G1337gat));
  NOR2_X1   g608(.A1(new_n787), .A2(new_n702), .ZN(new_n810));
  XNOR2_X1  g609(.A(KEYINPUT114), .B(G99gat), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n704), .A2(new_n690), .A3(new_n811), .ZN(new_n812));
  OAI22_X1  g611(.A1(new_n810), .A2(new_n811), .B1(new_n793), .B2(new_n812), .ZN(G1338gat));
  NAND3_X1  g612(.A1(new_n723), .A2(new_n261), .A3(new_n786), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(G106gat), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n456), .A2(G106gat), .A3(new_n710), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n792), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT53), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n815), .A2(new_n817), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(G1339gat));
  NAND3_X1  g621(.A1(new_n765), .A2(new_n724), .A3(new_n710), .ZN(new_n823));
  INV_X1    g622(.A(new_n686), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n825), .B1(new_n670), .B2(new_n673), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n674), .A2(new_n826), .A3(new_n679), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n683), .B1(new_n688), .B2(new_n825), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n824), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n827), .A2(KEYINPUT55), .A3(new_n828), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n540), .A2(new_n548), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n536), .B1(new_n834), .B2(new_n551), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n557), .B1(new_n553), .B2(new_n555), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n565), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT115), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n839), .B(new_n565), .C1(new_n835), .C2(new_n836), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n657), .A2(new_n841), .A3(new_n573), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n833), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n574), .A2(new_n831), .A3(new_n832), .ZN(new_n844));
  INV_X1    g643(.A(new_n840), .ZN(new_n845));
  INV_X1    g644(.A(new_n551), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n846), .B1(new_n540), .B2(new_n548), .ZN(new_n847));
  OAI22_X1  g646(.A1(new_n556), .A2(new_n557), .B1(new_n847), .B2(new_n536), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n839), .B1(new_n848), .B2(new_n565), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n845), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n573), .A2(new_n690), .ZN(new_n851));
  OAI21_X1  g650(.A(KEYINPUT116), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT116), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n841), .A2(new_n853), .A3(new_n573), .A4(new_n690), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n844), .A2(new_n852), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n843), .B1(new_n855), .B2(new_n712), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n823), .B1(new_n856), .B2(new_n783), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n857), .A2(new_n411), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n363), .A2(new_n400), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(G113gat), .B1(new_n860), .B2(new_n724), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n468), .A2(new_n335), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n857), .A2(new_n401), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n457), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n574), .A2(new_n299), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n861), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  XOR2_X1   g665(.A(new_n866), .B(KEYINPUT117), .Z(G1340gat));
  NOR3_X1   g666(.A1(new_n860), .A2(new_n300), .A3(new_n710), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n863), .A2(new_n457), .A3(new_n690), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n868), .B1(new_n869), .B2(new_n300), .ZN(G1341gat));
  OAI21_X1  g669(.A(G127gat), .B1(new_n860), .B2(new_n621), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n621), .A2(G127gat), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n871), .B1(new_n864), .B2(new_n872), .ZN(G1342gat));
  OAI21_X1  g672(.A(G134gat), .B1(new_n860), .B2(new_n712), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(KEYINPUT119), .ZN(new_n875));
  INV_X1    g674(.A(G134gat), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n457), .A2(new_n657), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT118), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n863), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  XOR2_X1   g679(.A(new_n880), .B(KEYINPUT56), .Z(new_n881));
  NAND2_X1  g680(.A1(new_n875), .A2(new_n881), .ZN(G1343gat));
  AND2_X1   g681(.A1(new_n702), .A2(new_n859), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT57), .B1(new_n857), .B2(new_n261), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n261), .A2(KEYINPUT57), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n841), .A2(new_n573), .A3(new_n690), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n657), .B1(new_n844), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n621), .B1(new_n887), .B2(new_n843), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n885), .B1(new_n888), .B2(new_n823), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n574), .B(new_n883), .C1(new_n884), .C2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(G141gat), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT121), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n892), .B1(new_n469), .B2(new_n456), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n702), .A2(KEYINPUT121), .A3(new_n261), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n893), .A2(new_n401), .A3(new_n857), .A4(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n895), .A2(new_n363), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n724), .A2(G141gat), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT58), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n891), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  AOI22_X1  g699(.A1(new_n891), .A2(KEYINPUT120), .B1(new_n896), .B2(new_n897), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT120), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n890), .A2(new_n902), .A3(G141gat), .ZN(new_n903));
  AOI211_X1 g702(.A(KEYINPUT122), .B(new_n899), .C1(new_n901), .C2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n891), .A2(KEYINPUT120), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n906), .A2(new_n903), .A3(new_n898), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n905), .B1(new_n907), .B2(KEYINPUT58), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n900), .B1(new_n904), .B2(new_n908), .ZN(G1344gat));
  INV_X1    g708(.A(G148gat), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n896), .A2(new_n910), .A3(new_n690), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n883), .B1(new_n884), .B2(new_n889), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n912), .A2(new_n710), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT59), .ZN(new_n914));
  AND3_X1   g713(.A1(new_n913), .A2(new_n914), .A3(G148gat), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n857), .A2(KEYINPUT57), .A3(new_n261), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n888), .A2(new_n823), .ZN(new_n917));
  AOI21_X1  g716(.A(KEYINPUT57), .B1(new_n917), .B2(new_n261), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n920), .A2(new_n690), .A3(new_n883), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n914), .B1(new_n921), .B2(G148gat), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n911), .B1(new_n915), .B2(new_n922), .ZN(G1345gat));
  OAI21_X1  g722(.A(G155gat), .B1(new_n912), .B2(new_n621), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n896), .A2(new_n213), .A3(new_n783), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1346gat));
  OAI21_X1  g725(.A(G162gat), .B1(new_n912), .B2(new_n712), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n879), .A2(new_n214), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n895), .B2(new_n928), .ZN(G1347gat));
  NOR2_X1   g728(.A1(new_n457), .A2(new_n401), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n858), .A2(new_n930), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n931), .A2(new_n268), .A3(new_n724), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n857), .A2(new_n400), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n933), .A2(KEYINPUT123), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n457), .B1(new_n933), .B2(KEYINPUT123), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n934), .A2(new_n935), .A3(new_n862), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT124), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n934), .A2(new_n935), .A3(KEYINPUT124), .A4(new_n862), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n938), .A2(new_n574), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n932), .B1(new_n940), .B2(new_n268), .ZN(G1348gat));
  NAND4_X1  g740(.A1(new_n938), .A2(new_n269), .A3(new_n690), .A4(new_n939), .ZN(new_n942));
  OAI21_X1  g741(.A(G176gat), .B1(new_n931), .B2(new_n710), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1349gat));
  OAI21_X1  g743(.A(G183gat), .B1(new_n931), .B2(new_n621), .ZN(new_n945));
  OR2_X1    g744(.A1(new_n621), .A2(new_n286), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n945), .B1(new_n936), .B2(new_n946), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g747(.A(G190gat), .B1(new_n931), .B2(new_n712), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT61), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n712), .A2(G190gat), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n938), .A2(new_n939), .A3(new_n951), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n952), .A2(KEYINPUT125), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n952), .A2(KEYINPUT125), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n950), .B1(new_n953), .B2(new_n954), .ZN(G1351gat));
  AND2_X1   g754(.A1(new_n934), .A2(new_n935), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n469), .A2(new_n456), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g758(.A(G197gat), .B1(new_n959), .B2(new_n574), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n702), .A2(new_n930), .ZN(new_n961));
  OR3_X1    g760(.A1(new_n916), .A2(KEYINPUT126), .A3(new_n918), .ZN(new_n962));
  OAI21_X1  g761(.A(KEYINPUT126), .B1(new_n916), .B2(new_n918), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n574), .A2(G197gat), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n960), .B1(new_n964), .B2(new_n965), .ZN(G1352gat));
  INV_X1    g765(.A(KEYINPUT127), .ZN(new_n967));
  INV_X1    g766(.A(G204gat), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n968), .B1(new_n964), .B2(new_n690), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n710), .A2(G204gat), .ZN(new_n970));
  NAND4_X1  g769(.A1(new_n934), .A2(new_n935), .A3(new_n957), .A4(new_n970), .ZN(new_n971));
  OR2_X1    g770(.A1(new_n971), .A2(KEYINPUT62), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(KEYINPUT62), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n967), .B1(new_n969), .B2(new_n974), .ZN(new_n975));
  INV_X1    g774(.A(new_n961), .ZN(new_n976));
  INV_X1    g775(.A(new_n963), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n916), .A2(new_n918), .A3(KEYINPUT126), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g778(.A(G204gat), .B1(new_n979), .B2(new_n710), .ZN(new_n980));
  NAND4_X1  g779(.A1(new_n980), .A2(KEYINPUT127), .A3(new_n973), .A4(new_n972), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n975), .A2(new_n981), .ZN(G1353gat));
  INV_X1    g781(.A(G211gat), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n961), .A2(new_n621), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n983), .B1(new_n920), .B2(new_n984), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n985), .B(KEYINPUT63), .ZN(new_n986));
  OR2_X1    g785(.A1(new_n621), .A2(new_n225), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n986), .B1(new_n958), .B2(new_n987), .ZN(G1354gat));
  AOI21_X1  g787(.A(G218gat), .B1(new_n959), .B2(new_n657), .ZN(new_n989));
  AND2_X1   g788(.A1(new_n657), .A2(G218gat), .ZN(new_n990));
  AOI21_X1  g789(.A(new_n989), .B1(new_n964), .B2(new_n990), .ZN(G1355gat));
endmodule


