//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 0 0 0 1 1 0 0 0 1 1 0 0 0 0 1 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 0 0 0 0 1 1 1 0 1 0 0 0 0 0 1 1 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1261, new_n1262, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI211_X1 g0005(.A(G50), .B(G77), .C1(new_n203), .C2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(G250), .B1(G257), .B2(G264), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OR2_X1    g0015(.A1(new_n215), .A2(KEYINPUT0), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n203), .A2(new_n205), .ZN(new_n217));
  INV_X1    g0017(.A(G50), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n220), .A2(new_n209), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n215), .A2(KEYINPUT0), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n216), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT65), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT66), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n211), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT67), .ZN(new_n233));
  INV_X1    g0033(.A(KEYINPUT1), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AND2_X1   g0035(.A1(new_n233), .A2(new_n234), .ZN(new_n236));
  NOR3_X1   g0036(.A1(new_n225), .A2(new_n235), .A3(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G50), .B(G58), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G68), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XOR2_X1   g0050(.A(G107), .B(G116), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n249), .B(new_n252), .Z(G351));
  INV_X1    g0053(.A(KEYINPUT70), .ZN(new_n254));
  AND2_X1   g0054(.A1(KEYINPUT69), .A2(G1), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT69), .A2(G1), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G41), .A2(G45), .ZN(new_n257));
  NOR3_X1   g0057(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G1), .A3(G13), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n254), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT69), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n208), .ZN(new_n264));
  INV_X1    g0064(.A(G41), .ZN(new_n265));
  INV_X1    g0065(.A(G45), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(KEYINPUT69), .A2(G1), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n264), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(KEYINPUT70), .A3(new_n260), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n262), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G226), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n257), .A2(G1), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(new_n260), .A3(G274), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  OR2_X1    g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AND2_X1   g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NOR2_X1   g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI22_X1  g0081(.A1(new_n278), .A2(G223), .B1(new_n281), .B2(G77), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n276), .A2(new_n277), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(G222), .A3(new_n275), .ZN(new_n284));
  AND2_X1   g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n272), .B(new_n274), .C1(new_n260), .C2(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT73), .B(G200), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G190), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n289), .B1(new_n290), .B2(new_n286), .ZN(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n220), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n209), .B1(new_n217), .B2(new_n218), .ZN(new_n294));
  XNOR2_X1  g0094(.A(KEYINPUT8), .B(G58), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n209), .A2(G33), .ZN(new_n296));
  INV_X1    g0096(.A(G150), .ZN(new_n297));
  INV_X1    g0097(.A(G33), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n209), .A2(new_n298), .ZN(new_n299));
  OAI22_X1  g0099(.A1(new_n295), .A2(new_n296), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n293), .B1(new_n294), .B2(new_n300), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n264), .A2(G13), .A3(G20), .A4(new_n268), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n218), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n264), .A2(new_n268), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n304), .A2(new_n209), .ZN(new_n305));
  INV_X1    g0105(.A(new_n293), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT71), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n302), .A2(new_n306), .A3(KEYINPUT71), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n305), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n303), .B1(new_n311), .B2(new_n218), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT72), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n312), .A2(new_n313), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n301), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT9), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n291), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT10), .ZN(new_n319));
  OAI211_X1 g0119(.A(KEYINPUT9), .B(new_n301), .C1(new_n314), .C2(new_n315), .ZN(new_n320));
  AND3_X1   g0120(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n319), .B1(new_n318), .B2(new_n320), .ZN(new_n322));
  INV_X1    g0122(.A(new_n316), .ZN(new_n323));
  INV_X1    g0123(.A(G169), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n286), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(G179), .B2(new_n286), .ZN(new_n326));
  OAI22_X1  g0126(.A1(new_n321), .A2(new_n322), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n295), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n255), .A2(new_n256), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G20), .ZN(new_n330));
  AND3_X1   g0130(.A1(new_n302), .A2(new_n306), .A3(KEYINPUT71), .ZN(new_n331));
  AOI21_X1  g0131(.A(KEYINPUT71), .B1(new_n302), .B2(new_n306), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n328), .B(new_n330), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n302), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n295), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n276), .A2(new_n209), .A3(new_n277), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT7), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n276), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n277), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n202), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(G58), .A2(G68), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n203), .A2(new_n205), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(G20), .ZN(new_n344));
  INV_X1    g0144(.A(new_n299), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G159), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(KEYINPUT16), .B1(new_n341), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(KEYINPUT7), .B1(new_n281), .B2(new_n209), .ZN(new_n349));
  NOR4_X1   g0149(.A1(new_n279), .A2(new_n280), .A3(new_n338), .A4(G20), .ZN(new_n350));
  OAI21_X1  g0150(.A(G68), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT16), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n343), .A2(G20), .B1(G159), .B2(new_n345), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n348), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n336), .B1(new_n355), .B2(new_n293), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n269), .A2(G232), .A3(new_n260), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(KEYINPUT76), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT76), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n269), .A2(new_n359), .A3(G232), .A4(new_n260), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  AND3_X1   g0161(.A1(new_n273), .A2(new_n260), .A3(G274), .ZN(new_n362));
  OAI211_X1 g0162(.A(G223), .B(new_n275), .C1(new_n279), .C2(new_n280), .ZN(new_n363));
  OAI211_X1 g0163(.A(G226), .B(G1698), .C1(new_n279), .C2(new_n280), .ZN(new_n364));
  NAND2_X1  g0164(.A1(G33), .A2(G87), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n362), .B1(new_n366), .B2(new_n261), .ZN(new_n367));
  AND3_X1   g0167(.A1(new_n361), .A2(G190), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(G200), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n369), .B1(new_n361), .B2(new_n367), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n356), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT17), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n356), .A2(new_n371), .A3(KEYINPUT17), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n361), .A2(new_n367), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n324), .ZN(new_n378));
  INV_X1    g0178(.A(G179), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n361), .A2(new_n367), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(KEYINPUT18), .B1(new_n356), .B2(new_n381), .ZN(new_n382));
  AND3_X1   g0182(.A1(new_n361), .A2(new_n379), .A3(new_n367), .ZN(new_n383));
  AOI21_X1  g0183(.A(G169), .B1(new_n361), .B2(new_n367), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT18), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n306), .B1(new_n348), .B2(new_n354), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n385), .B(new_n386), .C1(new_n387), .C2(new_n336), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n382), .A2(new_n388), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n376), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n271), .A2(G244), .ZN(new_n391));
  NOR2_X1   g0191(.A1(G232), .A2(G1698), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n275), .A2(G238), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n283), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(G107), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n260), .B1(new_n281), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n362), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n391), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n398), .A2(new_n290), .ZN(new_n399));
  XOR2_X1   g0199(.A(KEYINPUT15), .B(G87), .Z(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n401), .A2(new_n296), .ZN(new_n402));
  INV_X1    g0202(.A(G77), .ZN(new_n403));
  OAI22_X1  g0203(.A1(new_n295), .A2(new_n299), .B1(new_n209), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n293), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n307), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n406), .A2(G77), .A3(new_n330), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n405), .B(new_n407), .C1(G77), .C2(new_n302), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n287), .B1(new_n391), .B2(new_n397), .ZN(new_n409));
  OR3_X1    g0209(.A1(new_n399), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n398), .A2(new_n324), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n391), .A2(new_n379), .A3(new_n397), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(new_n412), .A3(new_n408), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n302), .A2(G68), .ZN(new_n415));
  XNOR2_X1  g0215(.A(new_n415), .B(KEYINPUT12), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n406), .A2(G68), .A3(new_n330), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT11), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n202), .A2(G20), .ZN(new_n420));
  OAI221_X1 g0220(.A(new_n420), .B1(new_n296), .B2(new_n403), .C1(new_n218), .C2(new_n299), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n419), .B1(new_n421), .B2(new_n293), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n421), .A2(new_n419), .A3(new_n293), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n417), .B(new_n418), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(G238), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(new_n262), .B2(new_n270), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G33), .A2(G97), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT74), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT74), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n429), .A2(G33), .A3(G97), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(G226), .A2(G1698), .ZN(new_n432));
  INV_X1    g0232(.A(G232), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n432), .B1(new_n433), .B2(G1698), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n431), .B1(new_n283), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n274), .B1(new_n435), .B2(new_n260), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT13), .B1(new_n426), .B2(new_n436), .ZN(new_n437));
  AND3_X1   g0237(.A1(new_n269), .A2(KEYINPUT70), .A3(new_n260), .ZN(new_n438));
  AOI21_X1  g0238(.A(KEYINPUT70), .B1(new_n269), .B2(new_n260), .ZN(new_n439));
  OAI21_X1  g0239(.A(G238), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT13), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n433), .A2(G1698), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n442), .B1(G226), .B2(G1698), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n428), .B(new_n430), .C1(new_n443), .C2(new_n281), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n362), .B1(new_n444), .B2(new_n261), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n440), .A2(new_n441), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n437), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT14), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n447), .A2(new_n448), .A3(G169), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n437), .A2(G179), .A3(new_n446), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n448), .B1(new_n447), .B2(G169), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n424), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n437), .A2(G190), .A3(new_n446), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n418), .B1(new_n423), .B2(new_n422), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n455), .A2(new_n416), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n369), .B1(new_n437), .B2(new_n446), .ZN(new_n458));
  OAI21_X1  g0258(.A(KEYINPUT75), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n447), .A2(G200), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT75), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n460), .A2(new_n461), .A3(new_n456), .A4(new_n454), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n390), .A2(new_n414), .A3(new_n453), .A4(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n327), .A2(new_n464), .ZN(new_n465));
  OAI211_X1 g0265(.A(G264), .B(G1698), .C1(new_n279), .C2(new_n280), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT81), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT81), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n283), .A2(new_n468), .A3(G264), .A4(G1698), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(G257), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n471), .B1(new_n276), .B2(new_n277), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n472), .A2(new_n275), .B1(new_n281), .B2(G303), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n261), .ZN(new_n475));
  NOR3_X1   g0275(.A1(new_n255), .A2(new_n256), .A3(new_n266), .ZN(new_n476));
  XNOR2_X1  g0276(.A(KEYINPUT5), .B(G41), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n476), .A2(G274), .A3(new_n260), .A4(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n264), .A2(G45), .A3(new_n268), .ZN(new_n479));
  AND2_X1   g0279(.A1(KEYINPUT5), .A2(G41), .ZN(new_n480));
  NOR2_X1   g0280(.A1(KEYINPUT5), .A2(G41), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI211_X1 g0282(.A(G270), .B(new_n260), .C1(new_n479), .C2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n475), .A2(G179), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n260), .B1(new_n470), .B2(new_n473), .ZN(new_n487));
  OAI211_X1 g0287(.A(KEYINPUT21), .B(G169), .C1(new_n487), .C2(new_n484), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(G116), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n292), .A2(new_n220), .B1(G20), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(G33), .A2(G283), .ZN(new_n492));
  INV_X1    g0292(.A(G97), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n492), .B(new_n209), .C1(G33), .C2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n491), .A2(KEYINPUT20), .A3(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT82), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n491), .A2(KEYINPUT82), .A3(new_n494), .A4(KEYINPUT20), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n491), .A2(new_n494), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT20), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT83), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT83), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n500), .A2(new_n504), .A3(new_n501), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n499), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n264), .A2(G33), .A3(new_n268), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n302), .A2(new_n306), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G116), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(G116), .B2(new_n334), .ZN(new_n510));
  AOI21_X1  g0310(.A(KEYINPUT84), .B1(new_n506), .B2(new_n510), .ZN(new_n511));
  AND3_X1   g0311(.A1(new_n506), .A2(new_n510), .A3(KEYINPUT84), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n489), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n506), .A2(new_n510), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT84), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n475), .A2(G190), .A3(new_n485), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n506), .A2(new_n510), .A3(KEYINPUT84), .ZN(new_n518));
  OAI21_X1  g0318(.A(G200), .B1(new_n487), .B2(new_n484), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n516), .A2(new_n517), .A3(new_n518), .A4(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(G169), .B1(new_n487), .B2(new_n484), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n521), .B1(new_n516), .B2(new_n518), .ZN(new_n522));
  XNOR2_X1  g0322(.A(KEYINPUT85), .B(KEYINPUT21), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n513), .B(new_n520), .C1(new_n522), .C2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n334), .A2(new_n493), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n527), .B1(new_n508), .B2(new_n493), .ZN(new_n528));
  OAI21_X1  g0328(.A(G107), .B1(new_n349), .B2(new_n350), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n493), .A2(new_n395), .A3(KEYINPUT6), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT6), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(G97), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n395), .A2(KEYINPUT77), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT77), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G107), .ZN(new_n535));
  AND4_X1   g0335(.A1(new_n530), .A2(new_n532), .A3(new_n533), .A4(new_n535), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n530), .A2(new_n532), .B1(new_n533), .B2(new_n535), .ZN(new_n537));
  OAI21_X1  g0337(.A(G20), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n345), .A2(G77), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n529), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n528), .B1(new_n540), .B2(new_n293), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(G244), .B(new_n275), .C1(new_n279), .C2(new_n280), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT4), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n283), .A2(KEYINPUT4), .A3(G244), .A4(new_n275), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n283), .A2(G250), .A3(G1698), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n545), .A2(new_n546), .A3(new_n492), .A4(new_n547), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n548), .A2(new_n261), .ZN(new_n549));
  OAI211_X1 g0349(.A(G257), .B(new_n260), .C1(new_n479), .C2(new_n482), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n478), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n324), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n551), .B1(new_n261), .B2(new_n548), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n379), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n542), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n553), .A2(G190), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n556), .B(new_n541), .C1(new_n369), .C2(new_n553), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT87), .ZN(new_n559));
  OAI211_X1 g0359(.A(G264), .B(new_n260), .C1(new_n479), .C2(new_n482), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(G250), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n562), .A2(G1698), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(new_n279), .B2(new_n280), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT86), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n283), .A2(G257), .A3(G1698), .ZN(new_n567));
  NAND2_X1  g0367(.A1(G33), .A2(G294), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n563), .B(KEYINPUT86), .C1(new_n280), .C2(new_n279), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n566), .A2(new_n567), .A3(new_n568), .A4(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n561), .B1(new_n570), .B2(new_n261), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n571), .A2(new_n290), .A3(new_n478), .ZN(new_n572));
  AOI21_X1  g0372(.A(G200), .B1(new_n571), .B2(new_n478), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n209), .B(G87), .C1(new_n279), .C2(new_n280), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(KEYINPUT22), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT22), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n283), .A2(new_n577), .A3(new_n209), .A4(G87), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT24), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT23), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(new_n209), .B2(G107), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n395), .A2(KEYINPUT23), .A3(G20), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n298), .A2(G20), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n582), .A2(new_n583), .B1(new_n584), .B2(G116), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n579), .A2(new_n580), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n580), .B1(new_n579), .B2(new_n585), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n293), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n406), .A2(G107), .A3(new_n507), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n302), .A2(G107), .ZN(new_n590));
  XNOR2_X1  g0390(.A(new_n590), .B(KEYINPUT25), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n588), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n559), .B1(new_n574), .B2(new_n592), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n591), .A2(new_n589), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n588), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n571), .A2(new_n290), .A3(new_n478), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n570), .A2(new_n261), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n597), .A2(new_n478), .A3(new_n560), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n596), .B1(new_n598), .B2(G200), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n595), .A2(new_n599), .A3(KEYINPUT87), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n558), .B1(new_n593), .B2(new_n600), .ZN(new_n601));
  OAI211_X1 g0401(.A(G238), .B(new_n275), .C1(new_n279), .C2(new_n280), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT78), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT78), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n283), .A2(new_n604), .A3(G238), .A4(new_n275), .ZN(new_n605));
  NAND2_X1  g0405(.A1(G33), .A2(G116), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n283), .A2(G244), .A3(G1698), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n603), .A2(new_n605), .A3(new_n606), .A4(new_n607), .ZN(new_n608));
  OR2_X1    g0408(.A1(new_n479), .A2(G274), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n261), .B1(new_n479), .B2(new_n562), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n608), .A2(new_n261), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n379), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n608), .A2(new_n261), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n610), .A2(new_n609), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n324), .ZN(new_n616));
  INV_X1    g0416(.A(G87), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n617), .A2(new_n493), .A3(new_n395), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT19), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n619), .B1(new_n428), .B2(new_n430), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n618), .B1(new_n620), .B2(G20), .ZN(new_n621));
  AOI21_X1  g0421(.A(G20), .B1(new_n276), .B2(new_n277), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n584), .A2(G97), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n622), .A2(G68), .B1(new_n623), .B2(new_n619), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n306), .B1(new_n621), .B2(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n302), .A2(new_n400), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT80), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n302), .A2(new_n400), .A3(new_n306), .A4(new_n507), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT79), .ZN(new_n630));
  XNOR2_X1  g0430(.A(new_n629), .B(new_n630), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n627), .A2(new_n628), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n628), .B1(new_n627), .B2(new_n631), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n612), .B(new_n616), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n571), .A2(new_n478), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n324), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n571), .A2(new_n379), .A3(new_n478), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n592), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n611), .A2(G190), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n508), .A2(new_n617), .ZN(new_n640));
  NOR3_X1   g0440(.A1(new_n625), .A2(new_n640), .A3(new_n626), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n639), .B(new_n641), .C1(new_n287), .C2(new_n611), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n634), .A2(new_n638), .A3(new_n642), .ZN(new_n643));
  AND4_X1   g0443(.A1(new_n465), .A2(new_n526), .A3(new_n601), .A4(new_n643), .ZN(G372));
  NOR2_X1   g0444(.A1(new_n323), .A2(new_n326), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n382), .A2(new_n388), .ZN(new_n646));
  NOR3_X1   g0446(.A1(new_n426), .A2(new_n436), .A3(KEYINPUT13), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n441), .B1(new_n440), .B2(new_n445), .ZN(new_n648));
  OAI21_X1  g0448(.A(G169), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(KEYINPUT14), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n650), .A2(new_n450), .A3(new_n449), .ZN(new_n651));
  INV_X1    g0451(.A(new_n457), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n460), .ZN(new_n653));
  INV_X1    g0453(.A(new_n413), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n424), .A2(new_n651), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n646), .B1(new_n655), .B2(new_n376), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT90), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n322), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n656), .A2(new_n657), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n645), .B1(new_n658), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT89), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n637), .B1(new_n598), .B2(G169), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n663), .B1(new_n595), .B2(new_n664), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n592), .A2(KEYINPUT89), .A3(new_n636), .A4(new_n637), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n521), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(new_n512), .B2(new_n511), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n516), .A2(new_n518), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n669), .A2(new_n523), .B1(new_n670), .B2(new_n489), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n639), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n641), .B1(new_n287), .B2(new_n611), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n673), .B1(new_n674), .B2(KEYINPUT88), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT88), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n641), .B(new_n676), .C1(new_n287), .C2(new_n611), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n627), .A2(new_n631), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(KEYINPUT80), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n627), .A2(new_n628), .A3(new_n631), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n616), .A2(new_n612), .ZN(new_n682));
  AOI22_X1  g0482(.A1(new_n675), .A2(new_n677), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n672), .A2(new_n601), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n555), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n634), .A2(new_n685), .A3(new_n642), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(KEYINPUT26), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n674), .A2(KEYINPUT88), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n688), .A2(new_n639), .A3(new_n677), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT26), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n689), .A2(new_n634), .A3(new_n690), .A4(new_n685), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n687), .A2(new_n634), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n465), .B1(new_n684), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n662), .A2(new_n693), .ZN(G369));
  INV_X1    g0494(.A(G13), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G20), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT91), .B1(new_n304), .B2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT91), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n329), .A2(new_n699), .A3(new_n696), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT27), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n698), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(G213), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n701), .B1(new_n698), .B2(new_n700), .ZN(new_n704));
  OAI21_X1  g0504(.A(KEYINPUT92), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n698), .A2(new_n700), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(KEYINPUT27), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT92), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n707), .A2(new_n708), .A3(G213), .A4(new_n702), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(G343), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n670), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n526), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n671), .B2(new_n713), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(G330), .ZN(new_n716));
  INV_X1    g0516(.A(new_n638), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n717), .B1(new_n593), .B2(new_n600), .ZN(new_n718));
  INV_X1    g0518(.A(new_n712), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n718), .B1(new_n595), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n717), .A2(new_n712), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n716), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n671), .A2(new_n712), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n718), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n665), .A2(new_n666), .A3(new_n719), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n725), .A2(new_n729), .ZN(G399));
  NOR2_X1   g0530(.A1(new_n213), .A2(G41), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n618), .A2(G116), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n732), .A2(G1), .A3(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n219), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n734), .B1(new_n735), .B2(new_n732), .ZN(new_n736));
  XNOR2_X1  g0536(.A(new_n736), .B(KEYINPUT28), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n671), .A2(new_n638), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n738), .A2(new_n601), .A3(new_n683), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n689), .A2(new_n634), .A3(new_n685), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(KEYINPUT26), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n634), .A2(new_n685), .A3(new_n690), .A4(new_n642), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n742), .A2(new_n634), .A3(new_n743), .ZN(new_n744));
  OAI211_X1 g0544(.A(KEYINPUT29), .B(new_n719), .C1(new_n740), .C2(new_n744), .ZN(new_n745));
  AND3_X1   g0545(.A1(new_n687), .A2(new_n634), .A3(new_n691), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n672), .A2(new_n601), .A3(new_n683), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n712), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n745), .B1(new_n748), .B2(KEYINPUT29), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n553), .B1(new_n478), .B2(new_n571), .ZN(new_n750));
  AOI21_X1  g0550(.A(G179), .B1(new_n475), .B2(new_n485), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT93), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n615), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n611), .A2(KEYINPUT93), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n750), .A2(new_n751), .A3(new_n753), .A4(new_n754), .ZN(new_n755));
  AND2_X1   g0555(.A1(new_n553), .A2(new_n571), .ZN(new_n756));
  NOR3_X1   g0556(.A1(new_n487), .A2(new_n379), .A3(new_n484), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n756), .A2(KEYINPUT30), .A3(new_n757), .A4(new_n611), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT30), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n553), .A2(new_n611), .A3(new_n571), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n759), .B1(new_n760), .B2(new_n486), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n755), .A2(new_n758), .A3(new_n761), .ZN(new_n762));
  AND3_X1   g0562(.A1(new_n762), .A2(KEYINPUT31), .A3(new_n712), .ZN(new_n763));
  AOI21_X1  g0563(.A(KEYINPUT31), .B1(new_n762), .B2(new_n712), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n526), .A2(new_n601), .A3(new_n643), .A4(new_n719), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G330), .ZN(new_n768));
  AND2_X1   g0568(.A1(new_n749), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n737), .B1(new_n769), .B2(G1), .ZN(G364));
  INV_X1    g0570(.A(new_n716), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n208), .B1(new_n696), .B2(G45), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n731), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n775), .B1(G330), .B2(new_n715), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n212), .A2(new_n283), .ZN(new_n777));
  INV_X1    g0577(.A(G355), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n777), .A2(new_n778), .B1(G116), .B2(new_n212), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n249), .A2(new_n266), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n213), .A2(new_n283), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n782), .B1(new_n219), .B2(new_n266), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n779), .B1(new_n780), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G13), .A2(G33), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(G20), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n220), .B1(G20), .B2(new_n324), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n774), .B1(new_n784), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n788), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n209), .A2(new_n379), .ZN(new_n793));
  NOR2_X1   g0593(.A1(G190), .A2(G200), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n283), .B1(new_n795), .B2(new_n403), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n209), .A2(G179), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(new_n794), .ZN(new_n798));
  INV_X1    g0598(.A(G159), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  XOR2_X1   g0600(.A(KEYINPUT94), .B(KEYINPUT32), .Z(new_n801));
  XNOR2_X1  g0601(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n793), .A2(G190), .A3(new_n369), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n796), .B(new_n802), .C1(G58), .C2(new_n804), .ZN(new_n805));
  NOR3_X1   g0605(.A1(new_n290), .A2(G179), .A3(G200), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(new_n209), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(new_n493), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n793), .A2(G200), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(new_n290), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(new_n218), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n809), .A2(G190), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n808), .B(new_n812), .C1(G68), .C2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n288), .A2(new_n797), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(new_n290), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(G87), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n815), .A2(G190), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(G107), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n805), .A2(new_n814), .A3(new_n817), .A4(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n283), .B1(new_n816), .B2(G303), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT97), .ZN(new_n822));
  INV_X1    g0622(.A(new_n798), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n804), .A2(G322), .B1(new_n823), .B2(G329), .ZN(new_n824));
  INV_X1    g0624(.A(G311), .ZN(new_n825));
  INV_X1    g0625(.A(new_n813), .ZN(new_n826));
  XOR2_X1   g0626(.A(KEYINPUT33), .B(G317), .Z(new_n827));
  OAI221_X1 g0627(.A(new_n824), .B1(new_n825), .B2(new_n795), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(G283), .B2(new_n818), .ZN(new_n829));
  XNOR2_X1  g0629(.A(KEYINPUT95), .B(G326), .ZN(new_n830));
  INV_X1    g0630(.A(G294), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n811), .A2(new_n830), .B1(new_n831), .B2(new_n807), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(KEYINPUT96), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n822), .A2(new_n829), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n792), .B1(new_n820), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n791), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n787), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n836), .B1(new_n715), .B2(new_n837), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n776), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(G396));
  OAI211_X1 g0640(.A(new_n414), .B(new_n719), .C1(new_n684), .C2(new_n692), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n712), .A2(new_n408), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n410), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n413), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n719), .A2(new_n654), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n841), .B1(new_n748), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n774), .B1(new_n848), .B2(new_n768), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n768), .B2(new_n848), .ZN(new_n850));
  INV_X1    g0650(.A(new_n774), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n788), .A2(new_n785), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n851), .B1(new_n403), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n795), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n804), .A2(G143), .B1(new_n854), .B2(G159), .ZN(new_n855));
  INV_X1    g0655(.A(G137), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n855), .B1(new_n811), .B2(new_n856), .C1(new_n297), .C2(new_n826), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(KEYINPUT34), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n818), .A2(G68), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n816), .A2(G50), .ZN(new_n860));
  INV_X1    g0660(.A(new_n807), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(G58), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n281), .B1(new_n823), .B2(G132), .ZN(new_n863));
  AND4_X1   g0663(.A1(new_n859), .A2(new_n860), .A3(new_n862), .A4(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(G303), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n811), .A2(new_n865), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n808), .B(new_n866), .C1(G283), .C2(new_n813), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n818), .A2(G87), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n283), .B1(new_n804), .B2(G294), .ZN(new_n869));
  AOI22_X1  g0669(.A1(G116), .A2(new_n854), .B1(new_n823), .B2(G311), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(G107), .B2(new_n816), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n858), .A2(new_n864), .B1(new_n867), .B2(new_n872), .ZN(new_n873));
  OAI221_X1 g0673(.A(new_n853), .B1(new_n792), .B2(new_n873), .C1(new_n847), .C2(new_n786), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n850), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(G384));
  OAI211_X1 g0676(.A(new_n378), .B(new_n380), .C1(new_n387), .C2(new_n336), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n709), .B(new_n705), .C1(new_n387), .C2(new_n336), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n372), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT37), .ZN(new_n880));
  AOI211_X1 g0680(.A(KEYINPUT100), .B(new_n880), .C1(new_n878), .C2(KEYINPUT99), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT100), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT99), .B1(new_n356), .B2(new_n710), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n882), .B1(new_n883), .B2(KEYINPUT37), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n879), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT99), .ZN(new_n886));
  NOR3_X1   g0686(.A1(new_n341), .A2(new_n347), .A3(KEYINPUT16), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n352), .B1(new_n351), .B2(new_n353), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n293), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n336), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n705), .A2(new_n709), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n886), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(KEYINPUT100), .B1(new_n893), .B2(new_n880), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n883), .A2(new_n882), .A3(KEYINPUT37), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n372), .A2(new_n877), .A3(new_n878), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n878), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n376), .B2(new_n389), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n885), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT38), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n885), .A2(new_n897), .A3(new_n899), .A4(KEYINPUT38), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT39), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n356), .A2(new_n371), .A3(KEYINPUT17), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT17), .B1(new_n356), .B2(new_n371), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n878), .B1(new_n646), .B2(new_n908), .ZN(new_n909));
  XNOR2_X1  g0709(.A(KEYINPUT102), .B(KEYINPUT37), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n372), .A2(new_n877), .A3(new_n878), .A4(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n880), .A2(KEYINPUT102), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n911), .B1(new_n879), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n901), .B1(new_n909), .B2(new_n913), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n903), .A2(new_n914), .ZN(new_n915));
  XOR2_X1   g0715(.A(KEYINPUT103), .B(KEYINPUT39), .Z(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n905), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT101), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n453), .B2(new_n712), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n651), .A2(KEYINPUT101), .A3(new_n424), .A4(new_n719), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n918), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n892), .A2(new_n424), .A3(G343), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n451), .A2(new_n452), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n924), .B1(new_n463), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n924), .B1(new_n458), .B2(new_n457), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n424), .B2(new_n651), .ZN(new_n928));
  OAI21_X1  g0728(.A(KEYINPUT98), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT98), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n652), .A2(new_n460), .B1(new_n712), .B2(new_n424), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n453), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n651), .B1(new_n459), .B2(new_n462), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n930), .B(new_n932), .C1(new_n933), .C2(new_n924), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n929), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(new_n845), .B2(new_n841), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n904), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n389), .A2(new_n710), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n923), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n465), .B(new_n745), .C1(KEYINPUT29), .C2(new_n748), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n662), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n939), .B(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(G330), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n903), .A2(new_n914), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n929), .A2(new_n934), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n846), .B1(new_n765), .B2(new_n766), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(KEYINPUT40), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT40), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n904), .A2(new_n949), .A3(new_n945), .A4(new_n946), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n465), .A2(new_n767), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n943), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n952), .B2(new_n951), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n942), .A2(new_n954), .B1(new_n304), .B2(new_n697), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n942), .B2(new_n954), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n536), .A2(new_n537), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n958), .A2(KEYINPUT35), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(KEYINPUT35), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n959), .A2(G116), .A3(new_n221), .A4(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT36), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n219), .A2(G77), .A3(new_n342), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(G50), .B2(new_n202), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n964), .A2(new_n695), .A3(new_n304), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n956), .A2(new_n962), .A3(new_n965), .ZN(G367));
  INV_X1    g0766(.A(new_n769), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n555), .B(new_n557), .C1(new_n719), .C2(new_n541), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n685), .A2(new_n712), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n729), .A2(new_n970), .ZN(new_n971));
  XOR2_X1   g0771(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT107), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n971), .B(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n727), .A2(new_n728), .ZN(new_n975));
  INV_X1    g0775(.A(new_n970), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT44), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n977), .B(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n974), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n724), .A2(KEYINPUT108), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n980), .B(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n727), .B1(new_n722), .B2(new_n726), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n771), .B(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n967), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n731), .B(KEYINPUT41), .Z(new_n986));
  OAI21_X1  g0786(.A(new_n772), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT105), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n970), .A2(new_n726), .A3(new_n718), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(KEYINPUT42), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n555), .B1(new_n968), .B2(new_n638), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n719), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n990), .A2(KEYINPUT104), .A3(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(KEYINPUT42), .B2(new_n989), .ZN(new_n994));
  AOI21_X1  g0794(.A(KEYINPUT104), .B1(new_n990), .B2(new_n992), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n988), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n719), .A2(new_n641), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n998), .A2(new_n634), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(new_n683), .B2(new_n998), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n996), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n996), .A2(new_n1000), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(KEYINPUT43), .ZN(new_n1004));
  OAI21_X1  g0804(.A(KEYINPUT43), .B1(new_n994), .B2(new_n995), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1001), .A2(new_n1005), .A3(new_n1002), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1004), .B(new_n1006), .C1(new_n725), .C2(new_n976), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1008), .A2(new_n724), .A3(new_n970), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n987), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1000), .A2(new_n787), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n789), .B1(new_n212), .B2(new_n401), .C1(new_n782), .C2(new_n244), .ZN(new_n1012));
  AND2_X1   g0812(.A1(new_n1012), .A2(new_n774), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT46), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n816), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1014), .B1(new_n1015), .B2(new_n490), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n816), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1016), .B(new_n1017), .C1(new_n831), .C2(new_n826), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(KEYINPUT109), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n818), .A2(G97), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n283), .B1(new_n823), .B2(G317), .ZN(new_n1021));
  INV_X1    g0821(.A(G283), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1021), .B1(new_n1022), .B2(new_n795), .C1(new_n865), .C2(new_n803), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n811), .A2(new_n825), .B1(new_n395), .B2(new_n807), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1019), .A2(new_n1020), .A3(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1018), .A2(KEYINPUT109), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n807), .A2(new_n202), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n283), .B1(new_n798), .B2(new_n856), .C1(new_n803), .C2(new_n297), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1028), .B(new_n1029), .C1(G143), .C2(new_n810), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n818), .A2(G77), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1030), .B(new_n1031), .C1(new_n201), .C2(new_n1015), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n813), .A2(G159), .B1(new_n854), .B2(G50), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT110), .Z(new_n1034));
  OAI22_X1  g0834(.A1(new_n1026), .A2(new_n1027), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT47), .Z(new_n1036));
  OAI211_X1 g0836(.A(new_n1011), .B(new_n1013), .C1(new_n792), .C2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1010), .A2(new_n1037), .ZN(G387));
  INV_X1    g0838(.A(KEYINPUT117), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n984), .A2(new_n769), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n731), .B(KEYINPUT116), .Z(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1039), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1040), .A2(KEYINPUT117), .A3(new_n1042), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1044), .B(new_n1045), .C1(new_n769), .C2(new_n984), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n266), .B1(new_n202), .B2(new_n403), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n733), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT111), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1047), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AND3_X1   g0850(.A1(new_n328), .A2(KEYINPUT50), .A3(new_n218), .ZN(new_n1051));
  AOI21_X1  g0851(.A(KEYINPUT50), .B1(new_n328), .B2(new_n218), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1050), .B1(new_n1049), .B2(new_n1048), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n781), .B(new_n1053), .C1(new_n241), .C2(new_n266), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1054), .B1(G107), .B2(new_n212), .C1(new_n733), .C2(new_n777), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n851), .B1(new_n1055), .B2(new_n789), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n1015), .A2(new_n403), .B1(new_n297), .B2(new_n798), .ZN(new_n1057));
  OR2_X1    g0857(.A1(new_n1057), .A2(KEYINPUT112), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(KEYINPUT112), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1058), .A2(new_n283), .A3(new_n1020), .A4(new_n1059), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT113), .Z(new_n1061));
  AOI22_X1  g0861(.A1(new_n804), .A2(G50), .B1(new_n854), .B2(G68), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n295), .B2(new_n826), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n401), .A2(new_n807), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n799), .B2(new_n811), .ZN(new_n1066));
  NOR3_X1   g0866(.A1(new_n1061), .A2(new_n1063), .A3(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n281), .B1(new_n798), .B2(new_n830), .ZN(new_n1068));
  XOR2_X1   g0868(.A(KEYINPUT114), .B(G322), .Z(new_n1069));
  AOI22_X1  g0869(.A1(G311), .A2(new_n813), .B1(new_n810), .B2(new_n1069), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n1070), .A2(KEYINPUT115), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(KEYINPUT115), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n804), .A2(G317), .B1(new_n854), .B2(G303), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT48), .ZN(new_n1075));
  OR2_X1    g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n816), .A2(G294), .B1(G283), .B2(new_n861), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT49), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1068), .B(new_n1081), .C1(G116), .C2(new_n818), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1067), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1056), .B1(new_n1084), .B2(new_n792), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n723), .B2(new_n787), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n773), .B2(new_n984), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1046), .A2(new_n1087), .ZN(G393));
  AOI21_X1  g0888(.A(new_n1043), .B1(new_n982), .B2(new_n1041), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n725), .B1(new_n974), .B2(new_n979), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(KEYINPUT118), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n974), .A2(new_n979), .A3(new_n725), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1090), .A2(KEYINPUT118), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1040), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1089), .A2(new_n1095), .ZN(new_n1096));
  OR3_X1    g0896(.A1(new_n1093), .A2(new_n772), .A3(new_n1094), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(G317), .A2(new_n810), .B1(new_n804), .B2(G311), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT52), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n819), .B1(new_n1015), .B2(new_n1022), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1069), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n281), .B1(new_n831), .B2(new_n795), .C1(new_n1101), .C2(new_n798), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n826), .A2(new_n865), .B1(new_n490), .B2(new_n807), .ZN(new_n1103));
  OR4_X1    g0903(.A1(new_n1099), .A2(new_n1100), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n283), .B1(new_n795), .B2(new_n295), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n826), .A2(new_n218), .B1(new_n403), .B2(new_n807), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1105), .B(new_n1106), .C1(G143), .C2(new_n823), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n811), .A2(new_n297), .B1(new_n799), .B2(new_n803), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT51), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n816), .A2(G68), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1107), .A2(new_n868), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n792), .B1(new_n1104), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n781), .A2(new_n252), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n790), .B1(G97), .B2(new_n213), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n851), .B(new_n1112), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT119), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n837), .B2(new_n970), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1096), .A2(new_n1097), .A3(new_n1117), .ZN(G390));
  AOI22_X1  g0918(.A1(KEYINPUT39), .A2(new_n904), .B1(new_n915), .B2(new_n916), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n785), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n852), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1121), .A2(new_n328), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n817), .A2(new_n281), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT121), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n795), .A2(new_n493), .B1(new_n798), .B2(new_n831), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(G116), .B2(new_n804), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n813), .A2(G107), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(G77), .A2(new_n861), .B1(new_n810), .B2(G283), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n859), .A2(new_n1126), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n826), .A2(new_n856), .B1(new_n799), .B2(new_n807), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(G128), .B2(new_n810), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n818), .A2(G50), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n281), .B1(new_n804), .B2(G132), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(KEYINPUT54), .B(G143), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n854), .A2(new_n1135), .B1(new_n823), .B2(G125), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1131), .A2(new_n1132), .A3(new_n1133), .A4(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n816), .A2(G150), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT53), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n1124), .A2(new_n1129), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n851), .B(new_n1122), .C1(new_n1140), .C2(new_n788), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1120), .A2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n915), .A2(new_n922), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n845), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n690), .B1(new_n683), .B2(new_n685), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n743), .A2(new_n634), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n712), .B1(new_n1147), .B2(new_n739), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1144), .B1(new_n1148), .B2(new_n844), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1143), .B1(new_n1149), .B2(new_n935), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n841), .A2(new_n845), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n922), .B1(new_n1151), .B2(new_n945), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1150), .B1(new_n1152), .B2(new_n918), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n945), .A2(new_n946), .A3(G330), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1119), .B1(new_n936), .B2(new_n922), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1157), .A2(new_n1150), .A3(new_n1154), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1142), .B1(new_n1159), .B2(new_n772), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n465), .A2(new_n767), .A3(G330), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n940), .A2(new_n662), .A3(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n767), .A2(G330), .A3(new_n847), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n935), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n1154), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n1151), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1149), .A2(new_n1165), .A3(new_n1154), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1163), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1156), .A2(new_n1158), .A3(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1170), .A2(KEYINPUT120), .A3(new_n1042), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1163), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1159), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1171), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(KEYINPUT120), .B1(new_n1170), .B2(new_n1042), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1161), .B1(new_n1176), .B2(new_n1177), .ZN(G378));
  INV_X1    g0978(.A(KEYINPUT123), .ZN(new_n1179));
  AND2_X1   g0979(.A1(new_n945), .A2(new_n946), .ZN(new_n1180));
  AOI21_X1  g0980(.A(KEYINPUT40), .B1(new_n902), .B2(new_n903), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n1180), .A2(new_n1181), .B1(new_n947), .B2(KEYINPUT40), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1179), .B1(new_n1182), .B2(new_n943), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n951), .A2(KEYINPUT123), .A3(G330), .ZN(new_n1184));
  XOR2_X1   g0984(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n327), .B(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n323), .A2(new_n710), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT122), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1187), .B(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1183), .A2(new_n1184), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n939), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1187), .B(new_n1189), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n951), .A2(G330), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1194), .A2(new_n1195), .A3(new_n1179), .ZN(new_n1196));
  AND3_X1   g0996(.A1(new_n1192), .A2(new_n1193), .A3(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1193), .B1(new_n1192), .B2(new_n1196), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1191), .A2(new_n785), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n774), .B1(G50), .B2(new_n1121), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n218), .B1(G33), .B2(G41), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n281), .B2(new_n265), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n265), .B(new_n281), .C1(new_n798), .C2(new_n1022), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n401), .A2(new_n795), .B1(new_n395), .B2(new_n803), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1204), .B(new_n1205), .C1(new_n816), .C2(G77), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n810), .A2(G116), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1028), .B1(G97), .B2(new_n813), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n818), .A2(G58), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT58), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1203), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(G128), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n803), .A2(new_n1213), .B1(new_n795), .B2(new_n856), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(G132), .B2(new_n813), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(G150), .A2(new_n861), .B1(new_n810), .B2(G125), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1215), .B(new_n1216), .C1(new_n1015), .C2(new_n1134), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1217), .A2(KEYINPUT59), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(KEYINPUT59), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n818), .A2(G159), .ZN(new_n1220));
  AOI211_X1 g1020(.A(G33), .B(G41), .C1(new_n823), .C2(G124), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1212), .B1(new_n1211), .B2(new_n1210), .C1(new_n1218), .C2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1201), .B1(new_n1223), .B2(new_n788), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1199), .A2(new_n773), .B1(new_n1200), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1170), .A2(new_n1173), .ZN(new_n1226));
  AOI21_X1  g1026(.A(KEYINPUT57), .B1(new_n1199), .B2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT57), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(new_n1170), .B2(new_n1173), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1192), .A2(new_n1196), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(new_n939), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1192), .A2(new_n1193), .A3(new_n1196), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1229), .A2(new_n1231), .A3(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n1042), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1225), .B1(new_n1227), .B2(new_n1234), .ZN(G375));
  NAND2_X1  g1035(.A1(new_n1172), .A2(new_n773), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n851), .B1(new_n202), .B2(new_n852), .ZN(new_n1237));
  OAI221_X1 g1037(.A(new_n1065), .B1(new_n811), .B2(new_n831), .C1(new_n490), .C2(new_n826), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n283), .B1(new_n823), .B2(G303), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n804), .A2(G283), .B1(new_n854), .B2(G107), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1031), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n1238), .B(new_n1241), .C1(G97), .C2(new_n816), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  OR2_X1    g1043(.A1(new_n1243), .A2(KEYINPUT124), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n816), .A2(G159), .B1(G128), .B2(new_n823), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(KEYINPUT125), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n813), .A2(new_n1135), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(G50), .A2(new_n861), .B1(new_n810), .B2(G132), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n283), .B1(new_n795), .B2(new_n297), .C1(new_n856), .C2(new_n803), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(G58), .B2(new_n818), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .A4(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1243), .A2(KEYINPUT124), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1244), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n1237), .B1(new_n792), .B2(new_n1253), .C1(new_n945), .C2(new_n786), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1236), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n986), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1167), .A2(new_n1163), .A3(new_n1168), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1174), .A2(new_n1257), .A3(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1256), .A2(new_n1259), .ZN(G381));
  NAND3_X1  g1060(.A1(new_n1046), .A2(new_n839), .A3(new_n1087), .ZN(new_n1261));
  OR4_X1    g1061(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1261), .ZN(new_n1262));
  OR4_X1    g1062(.A1(G387), .A2(new_n1262), .A3(G378), .A4(G375), .ZN(G407));
  INV_X1    g1063(.A(G378), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n711), .A2(G213), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1267));
  OAI211_X1 g1067(.A(G407), .B(G213), .C1(G375), .C2(new_n1267), .ZN(G409));
  OAI211_X1 g1068(.A(G378), .B(new_n1225), .C1(new_n1227), .C2(new_n1234), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1231), .A2(new_n1257), .A3(new_n1226), .A4(new_n1232), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1231), .A2(new_n773), .A3(new_n1232), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1200), .A2(new_n1224), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1270), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1264), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1269), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1265), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT60), .ZN(new_n1277));
  NOR3_X1   g1077(.A1(new_n1172), .A2(new_n1173), .A3(new_n1277), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1278), .A2(new_n1043), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1258), .B1(new_n1169), .B2(new_n1277), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1281), .A2(G384), .A3(new_n1256), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(G384), .B1(new_n1281), .B2(new_n1256), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1266), .A2(G2897), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  OAI211_X1 g1087(.A(G2897), .B(new_n1266), .C1(new_n1283), .C2(new_n1284), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(KEYINPUT61), .B1(new_n1276), .B2(new_n1290), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1285), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1292), .B1(new_n1276), .B2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n839), .B1(new_n1046), .B2(new_n1087), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1296), .A2(G390), .A3(new_n1261), .ZN(new_n1297));
  AOI21_X1  g1097(.A(G390), .B1(new_n1296), .B2(new_n1261), .ZN(new_n1298));
  OAI21_X1  g1098(.A(G387), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  AND2_X1   g1099(.A1(new_n1010), .A2(new_n1037), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1097), .A2(new_n1117), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1261), .ZN(new_n1302));
  OAI211_X1 g1102(.A(new_n1096), .B(new_n1301), .C1(new_n1302), .C2(new_n1295), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1296), .A2(G390), .A3(new_n1261), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1300), .A2(new_n1303), .A3(new_n1304), .ZN(new_n1305));
  AND2_X1   g1105(.A1(new_n1299), .A2(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1266), .B1(new_n1269), .B2(new_n1274), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1307), .A2(KEYINPUT63), .A3(new_n1285), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1291), .A2(new_n1294), .A3(new_n1306), .A4(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT62), .ZN(new_n1310));
  AND3_X1   g1110(.A1(new_n1307), .A2(new_n1310), .A3(new_n1285), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT61), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1312), .B1(new_n1307), .B2(new_n1289), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1310), .B1(new_n1307), .B2(new_n1285), .ZN(new_n1314));
  NOR3_X1   g1114(.A1(new_n1311), .A2(new_n1313), .A3(new_n1314), .ZN(new_n1315));
  AND3_X1   g1115(.A1(new_n1299), .A2(new_n1305), .A3(KEYINPUT127), .ZN(new_n1316));
  AOI21_X1  g1116(.A(KEYINPUT127), .B1(new_n1299), .B2(new_n1305), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1309), .B1(new_n1315), .B2(new_n1318), .ZN(G405));
  NAND2_X1  g1119(.A1(G375), .A2(new_n1264), .ZN(new_n1320));
  AND3_X1   g1120(.A1(new_n1320), .A2(new_n1293), .A3(new_n1269), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1293), .B1(new_n1320), .B2(new_n1269), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1318), .A2(new_n1323), .ZN(new_n1324));
  OAI22_X1  g1124(.A1(new_n1316), .A2(new_n1317), .B1(new_n1322), .B2(new_n1321), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(G402));
endmodule


