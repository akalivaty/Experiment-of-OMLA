//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 0 1 0 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT28), .ZN(new_n188));
  INV_X1    g002(.A(G131), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G137), .ZN(new_n191));
  INV_X1    g005(.A(G137), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G134), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n189), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT66), .B1(new_n192), .B2(G134), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT66), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(new_n190), .A3(G137), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n198));
  AOI22_X1  g012(.A1(new_n195), .A2(new_n197), .B1(new_n198), .B2(KEYINPUT11), .ZN(new_n199));
  OAI22_X1  g013(.A1(new_n198), .A2(KEYINPUT11), .B1(new_n190), .B2(G137), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT11), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n201), .A2(new_n192), .A3(KEYINPUT65), .A4(G134), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n199), .A2(new_n189), .A3(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n194), .B1(new_n204), .B2(KEYINPUT67), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G143), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G128), .ZN(new_n211));
  NOR3_X1   g025(.A1(new_n210), .A2(KEYINPUT1), .A3(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT1), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n209), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(G143), .B(G146), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(G128), .ZN(new_n216));
  NOR3_X1   g030(.A1(new_n212), .A2(new_n214), .A3(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n205), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n194), .A2(KEYINPUT67), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n199), .A2(new_n203), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G131), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(new_n204), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n210), .B1(KEYINPUT0), .B2(G128), .ZN(new_n223));
  XOR2_X1   g037(.A(KEYINPUT0), .B(G128), .Z(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(new_n215), .ZN(new_n225));
  OR2_X1    g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  AOI22_X1  g040(.A1(new_n218), .A2(new_n219), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(G116), .B(G119), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XOR2_X1   g044(.A(KEYINPUT2), .B(G113), .Z(new_n231));
  XNOR2_X1  g045(.A(new_n230), .B(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n227), .A2(KEYINPUT70), .A3(new_n232), .ZN(new_n233));
  OR3_X1    g047(.A1(new_n212), .A2(new_n214), .A3(new_n216), .ZN(new_n234));
  AND2_X1   g048(.A1(new_n204), .A2(KEYINPUT67), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n219), .B(new_n234), .C1(new_n235), .C2(new_n194), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n222), .A2(new_n226), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(new_n232), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AND2_X1   g054(.A1(new_n233), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT64), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n226), .A2(new_n242), .ZN(new_n243));
  OR3_X1    g057(.A1(new_n223), .A2(new_n225), .A3(new_n242), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n243), .A2(new_n222), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n236), .ZN(new_n246));
  INV_X1    g060(.A(new_n232), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n188), .B1(new_n241), .B2(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT28), .B1(new_n227), .B2(new_n232), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n250), .B(KEYINPUT74), .ZN(new_n251));
  OR3_X1    g065(.A1(new_n249), .A2(new_n251), .A3(KEYINPUT29), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT26), .B(G101), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT72), .B(KEYINPUT27), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n253), .B(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT71), .ZN(new_n256));
  INV_X1    g070(.A(G953), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(KEYINPUT71), .A2(G953), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G237), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(G210), .A3(new_n261), .ZN(new_n262));
  XOR2_X1   g076(.A(new_n255), .B(new_n262), .Z(new_n263));
  OAI211_X1 g077(.A(new_n233), .B(new_n240), .C1(new_n232), .C2(new_n227), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT28), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT76), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT76), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n264), .A2(new_n267), .A3(KEYINPUT28), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n251), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT29), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n252), .B(new_n263), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT69), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n227), .A2(new_n272), .A3(KEYINPUT30), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT30), .ZN(new_n274));
  AOI21_X1  g088(.A(KEYINPUT69), .B1(new_n246), .B2(new_n274), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n227), .A2(KEYINPUT30), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n247), .B(new_n273), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n277), .A2(new_n241), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n263), .A2(KEYINPUT29), .ZN(new_n279));
  AOI21_X1  g093(.A(G902), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n187), .B1(new_n271), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n233), .A2(new_n240), .A3(new_n263), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT73), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT73), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n233), .A2(new_n240), .A3(new_n285), .A4(new_n263), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n284), .A2(new_n277), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT31), .ZN(new_n288));
  INV_X1    g102(.A(new_n263), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n289), .B1(new_n249), .B2(new_n251), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT31), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n284), .A2(new_n277), .A3(new_n291), .A4(new_n286), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n288), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(G472), .A2(G902), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT32), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT32), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n293), .A2(new_n297), .A3(new_n294), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n296), .A2(new_n298), .B1(KEYINPUT75), .B2(new_n295), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n295), .A2(KEYINPUT75), .A3(new_n297), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n282), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n226), .A2(G125), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n303), .B1(G125), .B2(new_n217), .ZN(new_n304));
  INV_X1    g118(.A(G224), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n305), .A2(G953), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n304), .B(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT92), .B(KEYINPUT93), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n307), .B(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT88), .B(KEYINPUT5), .ZN(new_n310));
  INV_X1    g124(.A(G116), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n311), .A2(G119), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT89), .ZN(new_n314));
  INV_X1    g128(.A(new_n310), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n228), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT89), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n310), .A2(new_n317), .A3(new_n312), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n314), .A2(new_n316), .A3(G113), .A4(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n231), .A2(new_n228), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(G104), .A2(G107), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT79), .B(G104), .ZN(new_n323));
  OAI211_X1 g137(.A(G101), .B(new_n322), .C1(new_n323), .C2(G107), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT84), .ZN(new_n325));
  NOR2_X1   g139(.A1(KEYINPUT3), .A2(G107), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT79), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n328), .A2(G104), .ZN(new_n329));
  INV_X1    g143(.A(G104), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n330), .A2(KEYINPUT79), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n327), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  XOR2_X1   g146(.A(KEYINPUT81), .B(G101), .Z(new_n333));
  AND2_X1   g147(.A1(KEYINPUT3), .A2(G107), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n334), .B1(G104), .B2(new_n326), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n332), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G107), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n337), .B1(new_n329), .B2(new_n331), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT84), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n338), .A2(new_n339), .A3(G101), .A4(new_n322), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n325), .A2(new_n336), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT85), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT85), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n325), .A2(new_n343), .A3(new_n340), .A4(new_n336), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n321), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT90), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT80), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n332), .A2(new_n348), .A3(new_n335), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n330), .A2(KEYINPUT79), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n328), .A2(G104), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n326), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT3), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n353), .A2(new_n337), .A3(G104), .ZN(new_n354));
  NAND2_X1  g168(.A1(KEYINPUT3), .A2(G107), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT80), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n349), .A2(new_n357), .A3(G101), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT4), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n352), .A2(new_n356), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n359), .B1(new_n360), .B2(new_n333), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(KEYINPUT82), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n349), .A2(new_n357), .A3(new_n359), .A4(G101), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT82), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n358), .A2(new_n361), .A3(new_n365), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n363), .A2(new_n247), .A3(new_n364), .A4(new_n366), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n321), .A2(new_n342), .A3(KEYINPUT90), .A4(new_n344), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n347), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT91), .ZN(new_n370));
  XOR2_X1   g184(.A(G110), .B(G122), .Z(new_n371));
  INV_X1    g185(.A(KEYINPUT91), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n347), .A2(new_n367), .A3(new_n372), .A4(new_n368), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n370), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT6), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n369), .ZN(new_n377));
  INV_X1    g191(.A(new_n371), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n375), .B1(new_n374), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n309), .B1(new_n376), .B2(new_n380), .ZN(new_n381));
  XOR2_X1   g195(.A(new_n371), .B(KEYINPUT8), .Z(new_n382));
  AND2_X1   g196(.A1(new_n342), .A2(new_n344), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n228), .A2(KEYINPUT5), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n314), .A2(G113), .A3(new_n318), .A4(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n383), .A2(new_n320), .A3(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n386), .B(KEYINPUT94), .ZN(new_n387));
  INV_X1    g201(.A(new_n321), .ZN(new_n388));
  AND2_X1   g202(.A1(new_n388), .A2(new_n341), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n382), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(KEYINPUT7), .B1(new_n305), .B2(G953), .ZN(new_n391));
  XOR2_X1   g205(.A(new_n304), .B(new_n391), .Z(new_n392));
  AOI21_X1  g206(.A(new_n392), .B1(new_n377), .B2(new_n378), .ZN(new_n393));
  AOI21_X1  g207(.A(G902), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n381), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g209(.A(G210), .B1(G237), .B2(G902), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n381), .A2(new_n396), .A3(new_n394), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(G214), .B1(G237), .B2(G902), .ZN(new_n401));
  INV_X1    g215(.A(G125), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n402), .A2(KEYINPUT16), .A3(G140), .ZN(new_n403));
  XNOR2_X1  g217(.A(G125), .B(G140), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n403), .B1(new_n404), .B2(KEYINPUT16), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n405), .B(G146), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n260), .A2(G214), .A3(new_n261), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT95), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n407), .B1(new_n408), .B2(new_n208), .ZN(new_n409));
  XNOR2_X1  g223(.A(KEYINPUT95), .B(G143), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n260), .A2(new_n410), .A3(G214), .A4(new_n261), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G131), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT17), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n409), .A2(new_n189), .A3(new_n411), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT98), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n406), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n189), .B1(new_n409), .B2(new_n411), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT17), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n413), .A2(KEYINPUT98), .A3(new_n414), .A4(new_n415), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n418), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(G113), .B(G122), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n423), .B(new_n330), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n404), .B(new_n206), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT18), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n409), .B(new_n411), .C1(new_n426), .C2(new_n189), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n425), .B(new_n427), .C1(new_n413), .C2(new_n426), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n422), .A2(new_n424), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n405), .A2(G146), .ZN(new_n430));
  XOR2_X1   g244(.A(G125), .B(G140), .Z(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT19), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT19), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n404), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n430), .B1(new_n435), .B2(G146), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(KEYINPUT96), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT96), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n438), .B(new_n430), .C1(new_n435), .C2(G146), .ZN(new_n439));
  INV_X1    g253(.A(new_n415), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n437), .B(new_n439), .C1(new_n440), .C2(new_n419), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n424), .B1(new_n441), .B2(new_n428), .ZN(new_n442));
  OR2_X1    g256(.A1(new_n442), .A2(KEYINPUT97), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(KEYINPUT97), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n429), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G475), .ZN(new_n446));
  INV_X1    g260(.A(G902), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT20), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT20), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n445), .A2(new_n450), .A3(new_n446), .A4(new_n447), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  XOR2_X1   g266(.A(KEYINPUT9), .B(G234), .Z(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G217), .ZN(new_n455));
  NOR3_X1   g269(.A1(new_n454), .A2(new_n455), .A3(G953), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n211), .A2(G143), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n458), .B(KEYINPUT100), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n211), .A2(G143), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(KEYINPUT99), .ZN(new_n462));
  NOR3_X1   g276(.A1(new_n460), .A2(G134), .A3(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(G116), .B(G122), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(G107), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n459), .B1(new_n462), .B2(KEYINPUT13), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT101), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n462), .A2(KEYINPUT13), .ZN(new_n469));
  OAI211_X1 g283(.A(KEYINPUT101), .B(new_n459), .C1(new_n462), .C2(KEYINPUT13), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AOI211_X1 g285(.A(new_n463), .B(new_n465), .C1(new_n471), .C2(G134), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n464), .A2(new_n337), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n311), .A2(KEYINPUT14), .A3(G122), .ZN(new_n474));
  INV_X1    g288(.A(new_n464), .ZN(new_n475));
  OAI211_X1 g289(.A(G107), .B(new_n474), .C1(new_n475), .C2(KEYINPUT14), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n460), .A2(new_n462), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n477), .A2(new_n190), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n473), .B(new_n476), .C1(new_n478), .C2(new_n463), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n457), .B1(new_n472), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n465), .B1(new_n471), .B2(G134), .ZN(new_n482));
  INV_X1    g296(.A(new_n463), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n484), .A2(new_n479), .A3(new_n456), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n481), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT15), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(G478), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n486), .A2(new_n447), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n488), .B1(new_n486), .B2(new_n447), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(G952), .ZN(new_n492));
  AOI211_X1 g306(.A(G953), .B(new_n492), .C1(G234), .C2(G237), .ZN(new_n493));
  AOI211_X1 g307(.A(new_n447), .B(new_n260), .C1(G234), .C2(G237), .ZN(new_n494));
  XOR2_X1   g308(.A(KEYINPUT21), .B(G898), .Z(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n493), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n422), .A2(new_n428), .ZN(new_n499));
  INV_X1    g313(.A(new_n424), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n429), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n447), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(G475), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n452), .A2(new_n491), .A3(new_n498), .A4(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n400), .A2(new_n401), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(G221), .B1(new_n454), .B2(G902), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n260), .A2(G227), .ZN(new_n510));
  XOR2_X1   g324(.A(G110), .B(G140), .Z(new_n511));
  XNOR2_X1  g325(.A(new_n510), .B(new_n511), .ZN(new_n512));
  NOR3_X1   g326(.A1(new_n341), .A2(KEYINPUT10), .A3(new_n217), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n342), .A2(new_n234), .A3(new_n344), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n513), .B1(new_n514), .B2(KEYINPUT10), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n363), .A2(new_n226), .A3(new_n364), .A4(new_n366), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT83), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n358), .A2(new_n365), .A3(new_n361), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n365), .B1(new_n358), .B2(new_n361), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n521), .A2(KEYINPUT83), .A3(new_n226), .A4(new_n364), .ZN(new_n522));
  AOI211_X1 g336(.A(new_n222), .B(new_n515), .C1(new_n518), .C2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n222), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n522), .A2(new_n518), .ZN(new_n525));
  INV_X1    g339(.A(new_n515), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n512), .B1(new_n523), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT87), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n523), .A2(new_n512), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n383), .A2(new_n234), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n341), .A2(new_n217), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n222), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT12), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI211_X1 g350(.A(KEYINPUT12), .B(new_n222), .C1(new_n532), .C2(new_n533), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n531), .A2(new_n538), .ZN(new_n539));
  OAI211_X1 g353(.A(KEYINPUT87), .B(new_n512), .C1(new_n523), .C2(new_n527), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n530), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(G469), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n542), .A2(KEYINPUT86), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(KEYINPUT86), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n541), .A2(new_n447), .A3(new_n544), .A4(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n525), .A2(new_n526), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n538), .B1(new_n222), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n527), .ZN(new_n549));
  AOI22_X1  g363(.A1(new_n548), .A2(new_n512), .B1(new_n549), .B2(new_n531), .ZN(new_n550));
  OAI21_X1  g364(.A(G469), .B1(new_n550), .B2(G902), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n509), .B1(new_n546), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(G119), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n553), .A2(G128), .ZN(new_n554));
  OR2_X1    g368(.A1(new_n554), .A2(KEYINPUT23), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n211), .A2(G119), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n554), .A2(KEYINPUT23), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n555), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n556), .A2(new_n554), .ZN(new_n560));
  XOR2_X1   g374(.A(KEYINPUT24), .B(G110), .Z(new_n561));
  OAI22_X1  g375(.A1(new_n559), .A2(G110), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n562), .B(new_n430), .C1(G146), .C2(new_n431), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n559), .A2(G110), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n560), .A2(new_n561), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n406), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT22), .B(G137), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(KEYINPUT77), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n260), .A2(G221), .A3(G234), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n569), .B(new_n570), .ZN(new_n571));
  XOR2_X1   g385(.A(new_n567), .B(new_n571), .Z(new_n572));
  OR3_X1    g386(.A1(new_n572), .A2(KEYINPUT25), .A3(G902), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n455), .B1(G234), .B2(new_n447), .ZN(new_n574));
  OAI21_X1  g388(.A(KEYINPUT25), .B1(new_n572), .B2(G902), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT78), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n573), .A2(new_n575), .A3(KEYINPUT78), .A4(new_n574), .ZN(new_n579));
  OR3_X1    g393(.A1(new_n572), .A2(G902), .A3(new_n574), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n302), .A2(new_n507), .A3(new_n552), .A4(new_n582), .ZN(new_n583));
  XOR2_X1   g397(.A(new_n583), .B(new_n333), .Z(G3));
  AND3_X1   g398(.A1(new_n381), .A2(new_n396), .A3(new_n394), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n396), .B1(new_n381), .B2(new_n394), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n401), .B(new_n498), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n486), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(G902), .ZN(new_n589));
  XNOR2_X1  g403(.A(KEYINPUT102), .B(G478), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n486), .A2(KEYINPUT33), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT33), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n481), .A2(new_n485), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(G902), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n591), .B1(new_n595), .B2(G478), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n449), .A2(new_n451), .B1(G475), .B2(new_n503), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n587), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n293), .A2(new_n447), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(G472), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n295), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n600), .A2(new_n552), .A3(new_n582), .A4(new_n604), .ZN(new_n605));
  XOR2_X1   g419(.A(KEYINPUT34), .B(G104), .Z(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(G6));
  NAND2_X1  g421(.A1(new_n546), .A2(new_n551), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n508), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n609), .A2(new_n581), .A3(new_n603), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT103), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n504), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n503), .A2(KEYINPUT103), .A3(G475), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n612), .A2(new_n452), .A3(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n491), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n617), .A2(new_n587), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n610), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT35), .B(G107), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G9));
  INV_X1    g435(.A(KEYINPUT36), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n571), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(new_n623), .B(KEYINPUT104), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(new_n567), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n625), .B(new_n447), .C1(new_n455), .C2(G234), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n578), .A2(new_n579), .A3(new_n626), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n608), .A2(new_n508), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n507), .A2(new_n628), .A3(new_n604), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G110), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT105), .B(KEYINPUT37), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G12));
  NAND2_X1  g446(.A1(new_n295), .A2(KEYINPUT75), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n293), .A2(new_n297), .A3(new_n294), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n297), .B1(new_n293), .B2(new_n294), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n281), .B1(new_n636), .B2(new_n300), .ZN(new_n637));
  INV_X1    g451(.A(G900), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n493), .B1(new_n494), .B2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n401), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n491), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n643), .B1(new_n398), .B2(new_n399), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n640), .A2(new_n615), .A3(new_n628), .A4(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G128), .ZN(G30));
  XOR2_X1   g460(.A(new_n639), .B(KEYINPUT39), .Z(new_n647));
  NAND2_X1  g461(.A1(new_n552), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n648), .B(KEYINPUT40), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n400), .B(KEYINPUT38), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n650), .A2(new_n642), .ZN(new_n651));
  INV_X1    g465(.A(new_n264), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n287), .B1(new_n652), .B2(new_n263), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n187), .B1(new_n653), .B2(new_n447), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n654), .B1(new_n636), .B2(new_n300), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n655), .A2(new_n597), .A3(new_n627), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n649), .A2(new_n651), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G143), .ZN(G45));
  AOI21_X1  g472(.A(new_n641), .B1(new_n398), .B2(new_n399), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n596), .A2(new_n597), .A3(new_n639), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n659), .A2(KEYINPUT106), .A3(new_n660), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n628), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(KEYINPUT106), .B1(new_n659), .B2(new_n660), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n663), .A2(new_n637), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G146), .ZN(G48));
  NOR2_X1   g480(.A1(new_n637), .A2(new_n581), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n541), .A2(new_n447), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(G469), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT107), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n668), .A2(KEYINPUT107), .A3(G469), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n673), .A2(KEYINPUT108), .A3(new_n508), .A4(new_n546), .ZN(new_n674));
  AOI21_X1  g488(.A(KEYINPUT107), .B1(new_n668), .B2(G469), .ZN(new_n675));
  AOI211_X1 g489(.A(new_n670), .B(new_n542), .C1(new_n541), .C2(new_n447), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n508), .B(new_n546), .C1(new_n675), .C2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT108), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n667), .A2(new_n674), .A3(new_n679), .A4(new_n600), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT41), .B(G113), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G15));
  AND4_X1   g496(.A1(new_n667), .A2(new_n674), .A3(new_n679), .A4(new_n618), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(new_n311), .ZN(G18));
  AND3_X1   g498(.A1(new_n674), .A2(new_n679), .A3(new_n659), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n685), .A2(new_n302), .A3(new_n506), .A4(new_n627), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G119), .ZN(G21));
  INV_X1    g501(.A(new_n597), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n644), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n689), .A2(new_n497), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n581), .B(KEYINPUT111), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n288), .B1(new_n269), .B2(new_n263), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n692), .A2(KEYINPUT109), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n292), .B1(new_n692), .B2(KEYINPUT109), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n294), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT110), .B(G472), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n601), .A2(new_n696), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n691), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n674), .A2(new_n679), .A3(new_n690), .A4(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G122), .ZN(G24));
  NAND3_X1  g514(.A1(new_n695), .A2(new_n660), .A3(new_n697), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n685), .A2(new_n627), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G125), .ZN(G27));
  NAND3_X1  g518(.A1(new_n398), .A2(new_n401), .A3(new_n399), .ZN(new_n705));
  NOR4_X1   g519(.A1(new_n637), .A2(new_n609), .A3(new_n581), .A4(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n660), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n707), .A2(KEYINPUT42), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n707), .A2(new_n705), .ZN(new_n709));
  OAI21_X1  g523(.A(KEYINPUT112), .B1(new_n634), .B2(new_n635), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT112), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n296), .A2(new_n711), .A3(new_n298), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n710), .A2(new_n712), .A3(new_n282), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n709), .A2(new_n713), .A3(new_n552), .A4(new_n691), .ZN(new_n714));
  AOI22_X1  g528(.A1(new_n706), .A2(new_n708), .B1(new_n714), .B2(KEYINPUT42), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G131), .ZN(G33));
  INV_X1    g530(.A(new_n705), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n302), .A2(new_n582), .A3(new_n552), .A4(new_n717), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n718), .A2(new_n617), .A3(new_n639), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(new_n190), .ZN(G36));
  AND2_X1   g534(.A1(new_n595), .A2(G478), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n597), .B1(new_n721), .B2(new_n591), .ZN(new_n722));
  XOR2_X1   g536(.A(new_n722), .B(KEYINPUT43), .Z(new_n723));
  AND3_X1   g537(.A1(new_n723), .A2(new_n603), .A3(new_n627), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n705), .B1(new_n724), .B2(KEYINPUT44), .ZN(new_n725));
  XOR2_X1   g539(.A(new_n550), .B(KEYINPUT45), .Z(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(G469), .ZN(new_n727));
  NAND2_X1  g541(.A1(G469), .A2(G902), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n727), .A2(KEYINPUT46), .A3(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT46), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n730), .B(G469), .C1(new_n726), .C2(G902), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n729), .A2(new_n546), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n508), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n723), .A2(new_n603), .A3(new_n627), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n725), .A2(new_n647), .A3(new_n734), .A4(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G137), .ZN(G39));
  INV_X1    g553(.A(KEYINPUT47), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(KEYINPUT113), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n733), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n302), .A2(new_n582), .ZN(new_n743));
  OR2_X1    g557(.A1(new_n740), .A2(KEYINPUT113), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n744), .A2(new_n741), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n732), .A2(new_n508), .A3(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n742), .A2(new_n709), .A3(new_n743), .A4(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G140), .ZN(G42));
  AND2_X1   g563(.A1(new_n674), .A2(new_n679), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n750), .A2(new_n717), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n582), .A2(new_n493), .ZN(new_n752));
  AND4_X1   g566(.A1(new_n597), .A2(new_n751), .A3(new_n655), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n596), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n723), .A2(new_n493), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n751), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n695), .A2(new_n627), .A3(new_n697), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  AND3_X1   g573(.A1(new_n698), .A2(new_n723), .A3(new_n493), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n650), .A2(new_n401), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n750), .A3(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT50), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT51), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n673), .A2(new_n546), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n509), .ZN(new_n769));
  INV_X1    g583(.A(new_n747), .ZN(new_n770));
  AOI22_X1  g584(.A1(new_n732), .A2(new_n508), .B1(KEYINPUT113), .B2(new_n740), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n760), .A2(new_n717), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n767), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n754), .A2(new_n759), .A3(new_n766), .A4(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT48), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n713), .A2(new_n691), .ZN(new_n777));
  OR3_X1    g591(.A1(new_n756), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n776), .B1(new_n756), .B2(new_n777), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n492), .A2(G953), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n751), .A2(new_n598), .A3(new_n655), .A4(new_n752), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n775), .A2(new_n778), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n758), .B1(new_n753), .B2(new_n596), .ZN(new_n784));
  INV_X1    g598(.A(new_n769), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n785), .A2(KEYINPUT116), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(KEYINPUT116), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n786), .B(new_n787), .C1(new_n770), .C2(new_n771), .ZN(new_n788));
  AOI22_X1  g602(.A1(new_n788), .A2(new_n773), .B1(new_n764), .B2(new_n765), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT51), .B1(new_n784), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n783), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n685), .A2(new_n760), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n680), .A2(new_n699), .ZN(new_n793));
  INV_X1    g607(.A(new_n683), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n686), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n583), .A2(new_n605), .A3(new_n629), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n688), .A2(new_n491), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(KEYINPUT114), .B1(new_n798), .B2(new_n587), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n659), .A2(new_n800), .A3(new_n498), .A4(new_n797), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n610), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n796), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n639), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n706), .A2(new_n616), .A3(new_n615), .A4(new_n804), .ZN(new_n805));
  NOR4_X1   g619(.A1(new_n637), .A2(new_n616), .A3(new_n614), .A4(new_n639), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n628), .B(new_n717), .C1(new_n806), .C2(new_n702), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n803), .A2(new_n715), .A3(new_n805), .A4(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n795), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n674), .A2(new_n679), .A3(new_n659), .A4(new_n627), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n645), .B(new_n665), .C1(new_n811), .C2(new_n701), .ZN(new_n812));
  OR2_X1    g626(.A1(new_n689), .A2(new_n627), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n552), .A2(new_n804), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n813), .A2(new_n655), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n810), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n552), .A2(new_n627), .ZN(new_n817));
  NOR4_X1   g631(.A1(new_n637), .A2(new_n817), .A3(new_n614), .A4(new_n639), .ZN(new_n818));
  AOI22_X1  g632(.A1(new_n818), .A2(new_n644), .B1(new_n662), .B2(new_n664), .ZN(new_n819));
  INV_X1    g633(.A(new_n815), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n703), .A2(new_n819), .A3(new_n820), .A4(KEYINPUT52), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n816), .A2(new_n821), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n809), .A2(new_n822), .A3(KEYINPUT53), .ZN(new_n823));
  XNOR2_X1  g637(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n824), .B1(new_n812), .B2(new_n815), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n821), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT53), .B1(new_n809), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(KEYINPUT54), .B1(new_n823), .B2(new_n827), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n825), .A2(new_n821), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n302), .A2(new_n491), .A3(new_n615), .A4(new_n804), .ZN(new_n830));
  AOI211_X1 g644(.A(new_n817), .B(new_n705), .C1(new_n830), .C2(new_n701), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n610), .A2(new_n799), .A3(new_n801), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n832), .A2(new_n583), .A3(new_n605), .A4(new_n629), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n831), .A2(new_n833), .A3(new_n719), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n811), .A2(new_n637), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n683), .B1(new_n835), .B2(new_n506), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n834), .A2(new_n836), .A3(new_n715), .A4(new_n793), .ZN(new_n837));
  OAI21_X1  g651(.A(KEYINPUT53), .B1(new_n829), .B2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n809), .A2(new_n822), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n791), .A2(new_n792), .A3(new_n828), .A4(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n844), .B1(G952), .B2(G953), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n768), .B(KEYINPUT49), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n655), .A2(new_n508), .A3(new_n691), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n650), .A2(new_n641), .A3(new_n722), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n845), .A2(new_n849), .ZN(G75));
  INV_X1    g664(.A(new_n260), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(new_n492), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(KEYINPUT118), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n309), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n838), .A2(G210), .A3(G902), .A4(new_n840), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT56), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n376), .A2(new_n380), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(KEYINPUT117), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(KEYINPUT55), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n856), .A2(new_n857), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n860), .B1(new_n856), .B2(new_n857), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n855), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n856), .A2(new_n857), .ZN(new_n864));
  INV_X1    g678(.A(new_n860), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n856), .A2(new_n857), .A3(new_n860), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n866), .A2(new_n309), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n854), .B1(new_n863), .B2(new_n868), .ZN(G51));
  XOR2_X1   g683(.A(new_n728), .B(KEYINPUT57), .Z(new_n870));
  NOR2_X1   g684(.A1(new_n841), .A2(new_n842), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT54), .B1(new_n838), .B2(new_n840), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(new_n541), .ZN(new_n874));
  INV_X1    g688(.A(new_n727), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n838), .A2(G902), .A3(new_n875), .A4(new_n840), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT119), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n854), .B1(new_n874), .B2(new_n877), .ZN(G54));
  INV_X1    g692(.A(KEYINPUT120), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n809), .A2(new_n822), .A3(new_n839), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n839), .B1(new_n809), .B2(new_n826), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n882), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n883));
  INV_X1    g697(.A(new_n445), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n879), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n883), .A2(new_n884), .ZN(new_n886));
  AND4_X1   g700(.A1(KEYINPUT58), .A2(new_n838), .A3(G902), .A4(new_n840), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n887), .A2(KEYINPUT120), .A3(G475), .A4(new_n445), .ZN(new_n888));
  AND4_X1   g702(.A1(new_n853), .A2(new_n885), .A3(new_n886), .A4(new_n888), .ZN(G60));
  INV_X1    g703(.A(new_n592), .ZN(new_n890));
  INV_X1    g704(.A(new_n594), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(G478), .A2(G902), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT59), .Z(new_n894));
  NOR2_X1   g708(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n895), .B1(new_n871), .B2(new_n872), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n894), .B1(new_n843), .B2(new_n828), .ZN(new_n897));
  INV_X1    g711(.A(new_n892), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n896), .B(new_n853), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(G63));
  NAND2_X1  g714(.A1(G217), .A2(G902), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT60), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n838), .A2(new_n625), .A3(new_n840), .A4(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n853), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT61), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n572), .B1(new_n841), .B2(new_n902), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n906), .A2(KEYINPUT121), .A3(new_n907), .A4(new_n908), .ZN(new_n909));
  OR2_X1    g723(.A1(new_n907), .A2(KEYINPUT121), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n907), .A2(KEYINPUT121), .ZN(new_n911));
  INV_X1    g725(.A(new_n572), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n912), .B1(new_n882), .B2(new_n903), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n910), .B(new_n911), .C1(new_n913), .C2(new_n905), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n909), .A2(new_n914), .ZN(G66));
  OAI21_X1  g729(.A(G953), .B1(new_n496), .B2(new_n305), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n836), .A2(new_n793), .A3(new_n803), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n916), .B1(new_n918), .B2(new_n851), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n859), .B1(G898), .B2(new_n260), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n919), .B(new_n920), .ZN(G69));
  NAND2_X1  g735(.A1(new_n738), .A2(new_n748), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT62), .ZN(new_n923));
  INV_X1    g737(.A(new_n657), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n923), .B1(new_n924), .B2(new_n812), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n703), .A2(new_n657), .A3(new_n819), .A4(KEYINPUT62), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n922), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n648), .A2(new_n705), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n667), .B(new_n928), .C1(new_n598), .C2(new_n797), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n851), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n273), .B1(new_n275), .B2(new_n276), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n435), .B(KEYINPUT122), .Z(new_n932));
  XNOR2_X1  g746(.A(new_n931), .B(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  OR3_X1    g748(.A1(new_n930), .A2(KEYINPUT123), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n851), .A2(G900), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n734), .A2(new_n647), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n937), .A2(new_n689), .A3(new_n777), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n922), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n812), .A2(new_n719), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n939), .A2(new_n715), .A3(new_n940), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n934), .B(new_n936), .C1(new_n941), .C2(new_n851), .ZN(new_n942));
  OAI21_X1  g756(.A(KEYINPUT123), .B1(new_n930), .B2(new_n934), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n935), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(G227), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n851), .B1(new_n945), .B2(new_n638), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT124), .Z(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n944), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n935), .A2(new_n942), .A3(new_n943), .A4(new_n947), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(G72));
  NAND2_X1  g765(.A1(G472), .A2(G902), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT63), .Z(new_n953));
  OAI21_X1  g767(.A(new_n953), .B1(new_n941), .B2(new_n917), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n278), .B(KEYINPUT125), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n954), .A2(new_n289), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n287), .B1(new_n278), .B2(new_n263), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n953), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT126), .Z(new_n959));
  OAI21_X1  g773(.A(new_n959), .B1(new_n823), .B2(new_n827), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n956), .A2(new_n853), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n927), .A2(new_n918), .A3(new_n929), .ZN(new_n962));
  AOI211_X1 g776(.A(new_n289), .B(new_n955), .C1(new_n962), .C2(new_n953), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n961), .A2(new_n963), .ZN(G57));
endmodule


