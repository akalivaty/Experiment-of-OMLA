//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 0 1 0 1 1 1 0 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 0 1 0 0 0 1 0 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1275, new_n1276, new_n1277, new_n1278, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  AOI22_X1  g0007(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n208));
  INV_X1    g0008(.A(G68), .ZN(new_n209));
  INV_X1    g0009(.A(G238), .ZN(new_n210));
  OAI21_X1  g0010(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n212));
  INV_X1    g0012(.A(G116), .ZN(new_n213));
  INV_X1    g0013(.A(G270), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n211), .B(new_n215), .C1(G97), .C2(G257), .ZN(new_n216));
  INV_X1    g0016(.A(G58), .ZN(new_n217));
  INV_X1    g0017(.A(G232), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G20), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT64), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n220), .A2(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT0), .Z(new_n227));
  NOR2_X1   g0027(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G20), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n217), .A2(new_n209), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G50), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n223), .B(new_n228), .C1(new_n231), .C2(new_n233), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(new_n218), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT2), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT65), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G264), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n214), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n239), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(G107), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(new_n213), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  INV_X1    g0051(.A(G1), .ZN(new_n252));
  OAI211_X1 g0052(.A(new_n252), .B(G274), .C1(G41), .C2(G45), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G1), .A3(G13), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n252), .B1(G41), .B2(G45), .ZN(new_n257));
  AND3_X1   g0057(.A1(new_n256), .A2(G238), .A3(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  AND2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  OAI211_X1 g0061(.A(G226), .B(new_n259), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  OAI211_X1 g0062(.A(G232), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  INV_X1    g0064(.A(G97), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n262), .B(new_n263), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n256), .A2(KEYINPUT66), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT66), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n230), .A2(new_n268), .A3(new_n255), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  AOI211_X1 g0070(.A(new_n254), .B(new_n258), .C1(new_n266), .C2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT13), .ZN(new_n272));
  OAI21_X1  g0072(.A(KEYINPUT71), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT71), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n266), .A2(new_n270), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n253), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n274), .B(KEYINPUT13), .C1(new_n276), .C2(new_n258), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n271), .A2(new_n272), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n273), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G169), .ZN(new_n280));
  OR2_X1    g0080(.A1(new_n280), .A2(KEYINPUT14), .ZN(new_n281));
  AND2_X1   g0081(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n282));
  AND2_X1   g0082(.A1(new_n271), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n271), .A2(new_n282), .ZN(new_n284));
  OAI21_X1  g0084(.A(G179), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n280), .A2(KEYINPUT14), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n281), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G20), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G33), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(G20), .A2(G33), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n290), .A2(G77), .B1(new_n291), .B2(G50), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n292), .B1(new_n288), .B2(G68), .ZN(new_n293));
  NAND3_X1  g0093(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n229), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n293), .A2(KEYINPUT11), .A3(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n295), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n252), .A2(G20), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G68), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n296), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n252), .A2(G13), .A3(G20), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n303), .A2(G68), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n304), .B(KEYINPUT12), .ZN(new_n305));
  AOI21_X1  g0105(.A(KEYINPUT11), .B1(new_n293), .B2(new_n295), .ZN(new_n306));
  OR3_X1    g0106(.A1(new_n302), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n287), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT74), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n307), .B1(new_n279), .B2(G200), .ZN(new_n310));
  OAI21_X1  g0110(.A(G190), .B1(new_n283), .B2(new_n284), .ZN(new_n311));
  AND3_X1   g0111(.A1(new_n310), .A2(KEYINPUT73), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(KEYINPUT73), .B1(new_n310), .B2(new_n311), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n309), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n279), .A2(G200), .ZN(new_n315));
  INV_X1    g0115(.A(new_n307), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n315), .A2(new_n311), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT73), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n310), .A2(KEYINPUT73), .A3(new_n311), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n319), .A2(KEYINPUT74), .A3(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n308), .A2(new_n314), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n203), .A2(G20), .ZN(new_n323));
  INV_X1    g0123(.A(G150), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n288), .A2(new_n264), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n217), .A2(KEYINPUT8), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT8), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G58), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n326), .A2(new_n328), .A3(KEYINPUT67), .ZN(new_n329));
  OR3_X1    g0129(.A1(new_n327), .A2(KEYINPUT67), .A3(G58), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI221_X1 g0131(.A(new_n323), .B1(new_n324), .B2(new_n325), .C1(new_n331), .C2(new_n289), .ZN(new_n332));
  INV_X1    g0132(.A(new_n303), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n332), .A2(new_n295), .B1(new_n202), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n300), .A2(G50), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  OR2_X1    g0137(.A1(new_n337), .A2(KEYINPUT9), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT3), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n264), .ZN(new_n340));
  NAND2_X1  g0140(.A1(KEYINPUT3), .A2(G33), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(G223), .A3(G1698), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n342), .A2(G222), .A3(new_n259), .ZN(new_n344));
  INV_X1    g0144(.A(G77), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n343), .B(new_n344), .C1(new_n345), .C2(new_n342), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n270), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n256), .A2(new_n257), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(G226), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n347), .A2(new_n253), .A3(new_n349), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n337), .A2(KEYINPUT9), .B1(G200), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G190), .ZN(new_n352));
  OR2_X1    g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n338), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT10), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT10), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n338), .A2(new_n351), .A3(new_n356), .A4(new_n353), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NOR3_X1   g0158(.A1(new_n327), .A2(KEYINPUT67), .A3(G58), .ZN(new_n359));
  XNOR2_X1  g0159(.A(KEYINPUT8), .B(G58), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n359), .B1(new_n360), .B2(KEYINPUT67), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n361), .A2(KEYINPUT77), .A3(new_n298), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n329), .A2(new_n330), .A3(new_n298), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT77), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n362), .A2(new_n365), .A3(new_n297), .A4(new_n303), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n331), .A2(new_n333), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n256), .A2(G232), .A3(new_n257), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n253), .ZN(new_n370));
  OAI211_X1 g0170(.A(G226), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n371));
  OAI211_X1 g0171(.A(G223), .B(new_n259), .C1(new_n260), .C2(new_n261), .ZN(new_n372));
  NAND2_X1  g0172(.A1(G33), .A2(G87), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n370), .B1(new_n374), .B2(new_n270), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n352), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n376), .B1(G200), .B2(new_n375), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT75), .ZN(new_n378));
  NAND2_X1  g0178(.A1(G58), .A2(G68), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n288), .B1(new_n232), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n291), .A2(G159), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n378), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  AND2_X1   g0183(.A1(G58), .A2(G68), .ZN(new_n384));
  OAI21_X1  g0184(.A(G20), .B1(new_n384), .B2(new_n201), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n385), .A2(KEYINPUT75), .A3(new_n381), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n260), .A2(new_n261), .ZN(new_n388));
  AOI21_X1  g0188(.A(KEYINPUT7), .B1(new_n388), .B2(new_n288), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n340), .A2(KEYINPUT7), .A3(new_n288), .A4(new_n341), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(G68), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n387), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n340), .A2(new_n288), .A3(new_n341), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT7), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n396), .A2(KEYINPUT76), .A3(new_n390), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT76), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n394), .A2(new_n398), .A3(new_n395), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(G68), .A3(new_n399), .ZN(new_n400));
  NOR3_X1   g0200(.A1(new_n380), .A2(new_n382), .A3(KEYINPUT16), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n393), .A2(KEYINPUT16), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n368), .B(new_n377), .C1(new_n402), .C2(new_n297), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n403), .A2(KEYINPUT17), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT79), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  AND3_X1   g0206(.A1(new_n385), .A2(KEYINPUT75), .A3(new_n381), .ZN(new_n407));
  AOI21_X1  g0207(.A(KEYINPUT75), .B1(new_n385), .B2(new_n381), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n209), .B1(new_n396), .B2(new_n390), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT16), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n400), .A2(new_n401), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n295), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n414), .A2(KEYINPUT79), .A3(new_n368), .A4(new_n377), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n406), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n404), .B1(new_n416), .B2(KEYINPUT17), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT18), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n366), .A2(new_n367), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n420), .B1(new_n413), .B2(new_n295), .ZN(new_n421));
  AOI211_X1 g0221(.A(G179), .B(new_n370), .C1(new_n270), .C2(new_n374), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n374), .A2(new_n270), .ZN(new_n423));
  INV_X1    g0223(.A(new_n370), .ZN(new_n424));
  AOI21_X1  g0224(.A(G169), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT78), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(G179), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n423), .A2(new_n427), .A3(new_n424), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT78), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n428), .B(new_n429), .C1(G169), .C2(new_n375), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n419), .B1(new_n421), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n368), .B1(new_n402), .B2(new_n297), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n433), .A2(KEYINPUT18), .A3(new_n426), .A4(new_n430), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n358), .A2(new_n418), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT70), .ZN(new_n437));
  NAND2_X1  g0237(.A1(G20), .A2(G77), .ZN(new_n438));
  XNOR2_X1  g0238(.A(KEYINPUT15), .B(G87), .ZN(new_n439));
  OAI221_X1 g0239(.A(new_n438), .B1(new_n439), .B2(new_n289), .C1(new_n325), .C2(new_n360), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n440), .A2(new_n295), .B1(new_n345), .B2(new_n333), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n300), .A2(G77), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n342), .A2(G238), .A3(G1698), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n342), .A2(G232), .A3(new_n259), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n388), .A2(G107), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT69), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n444), .A2(new_n445), .A3(KEYINPUT69), .A4(new_n446), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n449), .A2(new_n270), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n348), .A2(G244), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n451), .A2(new_n253), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(G169), .ZN(new_n454));
  AOI211_X1 g0254(.A(new_n437), .B(new_n443), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n454), .ZN(new_n456));
  INV_X1    g0256(.A(new_n443), .ZN(new_n457));
  AOI21_X1  g0257(.A(KEYINPUT70), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n453), .A2(G179), .ZN(new_n459));
  NOR3_X1   g0259(.A1(new_n455), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n350), .A2(new_n454), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n336), .B(new_n462), .C1(G179), .C2(new_n350), .ZN(new_n463));
  XNOR2_X1  g0263(.A(new_n463), .B(KEYINPUT68), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n457), .B1(new_n453), .B2(G200), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n465), .B1(new_n352), .B2(new_n453), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n461), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  NOR3_X1   g0267(.A1(new_n322), .A2(new_n436), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n252), .A2(G33), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n303), .A2(new_n469), .A3(new_n229), .A4(new_n294), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT80), .ZN(new_n471));
  XNOR2_X1  g0271(.A(new_n470), .B(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G107), .ZN(new_n473));
  INV_X1    g0273(.A(G107), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n333), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g0275(.A(new_n475), .B(KEYINPUT25), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT22), .ZN(new_n478));
  OAI211_X1 g0278(.A(KEYINPUT86), .B(new_n288), .C1(new_n260), .C2(new_n261), .ZN(new_n479));
  INV_X1    g0279(.A(G87), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(G20), .B1(new_n340), .B2(new_n341), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n482), .A2(KEYINPUT86), .A3(KEYINPUT22), .A4(G87), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n290), .A2(G116), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n288), .A2(G107), .ZN(new_n485));
  XNOR2_X1  g0285(.A(new_n485), .B(KEYINPUT23), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n481), .A2(new_n483), .A3(new_n484), .A4(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT24), .ZN(new_n488));
  XNOR2_X1  g0288(.A(new_n487), .B(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n473), .B(new_n477), .C1(new_n489), .C2(new_n297), .ZN(new_n490));
  OAI211_X1 g0290(.A(G257), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n491));
  OAI211_X1 g0291(.A(G250), .B(new_n259), .C1(new_n260), .C2(new_n261), .ZN(new_n492));
  INV_X1    g0292(.A(G294), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n491), .B(new_n492), .C1(new_n264), .C2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n270), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT82), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT5), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n496), .B1(new_n497), .B2(G41), .ZN(new_n498));
  INV_X1    g0298(.A(G41), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n499), .A2(KEYINPUT82), .A3(KEYINPUT5), .ZN(new_n500));
  INV_X1    g0300(.A(G45), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(G1), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n497), .A2(G41), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n498), .A2(new_n500), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n504), .A2(G264), .A3(new_n256), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT87), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(G274), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n504), .A2(KEYINPUT87), .A3(G264), .A4(new_n256), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n495), .A2(new_n507), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(G200), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT90), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n512), .A2(KEYINPUT90), .A3(new_n513), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n495), .A2(new_n505), .A3(new_n510), .ZN(new_n519));
  OR2_X1    g0319(.A1(new_n519), .A2(G190), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n490), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n495), .A2(new_n507), .A3(new_n511), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT88), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n522), .A2(new_n523), .A3(G179), .A4(new_n510), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n519), .A2(G169), .ZN(new_n525));
  OAI21_X1  g0325(.A(KEYINPUT88), .B1(new_n512), .B2(new_n427), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT89), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n524), .A2(new_n526), .A3(KEYINPUT89), .A4(new_n525), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n521), .B1(new_n490), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n439), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n472), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n342), .A2(new_n288), .A3(G68), .ZN(new_n535));
  NAND3_X1  g0335(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n288), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(new_n206), .B2(G87), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT19), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(new_n289), .B2(new_n265), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n535), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n541), .A2(new_n295), .B1(new_n333), .B2(new_n439), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n534), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(G244), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n544));
  OAI211_X1 g0344(.A(G238), .B(new_n259), .C1(new_n260), .C2(new_n261), .ZN(new_n545));
  NAND2_X1  g0345(.A1(G33), .A2(G116), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n270), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n252), .A2(G45), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n549), .A2(new_n508), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n256), .A2(G250), .A3(new_n549), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n548), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n454), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n543), .B(new_n554), .C1(G179), .C2(new_n553), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n548), .A2(G190), .A3(new_n551), .A4(new_n552), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n470), .A2(new_n471), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n470), .A2(new_n471), .ZN(new_n558));
  OAI21_X1  g0358(.A(G87), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n559), .A2(KEYINPUT83), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT83), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n561), .B1(new_n472), .B2(G87), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n556), .B(new_n542), .C1(new_n560), .C2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n552), .ZN(new_n564));
  AOI211_X1 g0364(.A(new_n550), .B(new_n564), .C1(new_n547), .C2(new_n270), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n565), .A2(new_n513), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n555), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n303), .A2(G97), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n472), .A2(G97), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n397), .A2(G107), .A3(new_n399), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n291), .A2(G77), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n474), .A2(KEYINPUT6), .A3(G97), .ZN(new_n574));
  XOR2_X1   g0374(.A(G97), .B(G107), .Z(new_n575));
  OAI21_X1  g0375(.A(new_n574), .B1(new_n575), .B2(KEYINPUT6), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n572), .B(new_n573), .C1(new_n577), .C2(new_n288), .ZN(new_n578));
  AOI211_X1 g0378(.A(new_n569), .B(new_n571), .C1(new_n578), .C2(new_n295), .ZN(new_n579));
  OAI211_X1 g0379(.A(G244), .B(new_n259), .C1(new_n260), .C2(new_n261), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT4), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n342), .A2(KEYINPUT4), .A3(G244), .A4(new_n259), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n342), .A2(G250), .A3(G1698), .ZN(new_n584));
  NAND2_X1  g0384(.A1(G33), .A2(G283), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(KEYINPUT81), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT81), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n587), .A2(G33), .A3(G283), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n582), .A2(new_n583), .A3(new_n584), .A4(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n509), .B1(new_n590), .B2(new_n270), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n504), .A2(new_n256), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G257), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n513), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n591), .A2(new_n593), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n594), .B1(G190), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n579), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n578), .A2(new_n295), .ZN(new_n598));
  INV_X1    g0398(.A(new_n569), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n598), .A2(new_n570), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(G169), .B1(new_n591), .B2(new_n593), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n595), .A2(new_n427), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n568), .A2(new_n597), .A3(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT85), .ZN(new_n606));
  OAI211_X1 g0406(.A(G257), .B(new_n259), .C1(new_n260), .C2(new_n261), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT84), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n342), .A2(KEYINPUT84), .A3(G257), .A4(new_n259), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n388), .A2(G303), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n342), .A2(G264), .A3(G1698), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n609), .A2(new_n610), .A3(new_n611), .A4(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n270), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n504), .A2(G270), .A3(new_n256), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n614), .A2(G179), .A3(new_n616), .A4(new_n510), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n303), .A2(G116), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n470), .A2(new_n213), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT20), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n288), .B1(new_n265), .B2(G33), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n621), .B1(new_n586), .B2(new_n588), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n294), .A2(new_n229), .B1(G20), .B2(new_n213), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n620), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n586), .A2(new_n588), .ZN(new_n626));
  OAI211_X1 g0426(.A(KEYINPUT20), .B(new_n623), .C1(new_n626), .C2(new_n621), .ZN(new_n627));
  AOI211_X1 g0427(.A(new_n618), .B(new_n619), .C1(new_n625), .C2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n606), .B1(new_n617), .B2(new_n628), .ZN(new_n629));
  AOI211_X1 g0429(.A(new_n509), .B(new_n615), .C1(new_n613), .C2(new_n270), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n618), .B1(new_n625), .B2(new_n627), .ZN(new_n631));
  INV_X1    g0431(.A(new_n619), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n630), .A2(new_n633), .A3(KEYINPUT85), .A4(G179), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n629), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n614), .A2(new_n510), .A3(new_n616), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n636), .A2(new_n633), .A3(G169), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(KEYINPUT21), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT21), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n636), .A2(new_n633), .A3(new_n639), .A4(G169), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n636), .A2(G200), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n642), .B(new_n628), .C1(new_n352), .C2(new_n636), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n635), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n605), .A2(new_n644), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n468), .A2(new_n532), .A3(new_n645), .ZN(G372));
  OAI21_X1  g0446(.A(KEYINPUT91), .B1(new_n565), .B2(new_n513), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT91), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n553), .A2(new_n648), .A3(G200), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n555), .B1(new_n650), .B2(new_n563), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(KEYINPUT92), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT92), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n653), .B(new_n555), .C1(new_n650), .C2(new_n563), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n604), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(KEYINPUT93), .B1(new_n655), .B2(KEYINPUT26), .ZN(new_n656));
  INV_X1    g0456(.A(new_n604), .ZN(new_n657));
  INV_X1    g0457(.A(new_n654), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n541), .A2(new_n295), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n439), .A2(new_n333), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n559), .A2(KEYINPUT83), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n472), .A2(new_n561), .A3(G87), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n664), .A2(new_n556), .A3(new_n647), .A4(new_n649), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n653), .B1(new_n665), .B2(new_n555), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n657), .B1(new_n658), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT93), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT26), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n657), .A2(KEYINPUT26), .A3(new_n568), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n656), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n652), .A2(new_n654), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n490), .A2(new_n527), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n674), .A2(new_n635), .A3(new_n641), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n571), .B1(new_n578), .B2(new_n295), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n601), .B1(new_n676), .B2(new_n599), .ZN(new_n677));
  AOI22_X1  g0477(.A1(new_n677), .A2(new_n603), .B1(new_n579), .B2(new_n596), .ZN(new_n678));
  INV_X1    g0478(.A(new_n490), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n516), .A2(new_n520), .A3(new_n517), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n673), .A2(new_n675), .A3(new_n678), .A4(new_n681), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n682), .A2(new_n555), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n672), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n468), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n460), .B1(new_n312), .B2(new_n313), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n417), .B1(new_n308), .B2(new_n686), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n432), .A2(new_n434), .A3(KEYINPUT94), .ZN(new_n688));
  AOI21_X1  g0488(.A(KEYINPUT94), .B1(new_n432), .B2(new_n434), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n358), .B1(new_n687), .B2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n685), .A2(new_n464), .A3(new_n692), .ZN(G369));
  INV_X1    g0493(.A(G13), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(G20), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n252), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G213), .A3(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(G343), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(KEYINPUT95), .B1(new_n679), .B2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT95), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n490), .A2(new_n704), .A3(new_n701), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n532), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n701), .B1(new_n635), .B2(new_n641), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n490), .A2(new_n527), .A3(new_n702), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n679), .B1(new_n529), .B2(new_n530), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n701), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n706), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(G330), .ZN(new_n716));
  INV_X1    g0516(.A(new_n644), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(new_n628), .B2(new_n702), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n635), .A2(new_n641), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n719), .A2(new_n633), .A3(new_n701), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n716), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n715), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n712), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT96), .ZN(G399));
  INV_X1    g0525(.A(new_n225), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G41), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n728), .A2(G1), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(new_n233), .B2(new_n728), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n731), .B(KEYINPUT28), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n669), .B1(new_n604), .B2(new_n567), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT98), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI211_X1 g0535(.A(KEYINPUT98), .B(new_n669), .C1(new_n604), .C2(new_n567), .ZN(new_n736));
  OAI211_X1 g0536(.A(new_n735), .B(new_n736), .C1(new_n669), .C2(new_n667), .ZN(new_n737));
  AOI22_X1  g0537(.A1(new_n652), .A2(new_n654), .B1(new_n679), .B2(new_n680), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n738), .B(new_n678), .C1(new_n713), .C2(new_n719), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n737), .A2(new_n739), .A3(new_n555), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(new_n702), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(KEYINPUT29), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT30), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n595), .A2(new_n522), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n630), .A2(G179), .A3(new_n565), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(KEYINPUT97), .ZN(new_n747));
  OR3_X1    g0547(.A1(new_n744), .A2(new_n745), .A3(new_n743), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n565), .A2(G179), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n591), .A2(new_n593), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n749), .A2(new_n750), .A3(new_n636), .A4(new_n512), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT97), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n752), .B(new_n743), .C1(new_n744), .C2(new_n745), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n747), .A2(new_n748), .A3(new_n751), .A4(new_n753), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n754), .A2(new_n701), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n645), .A2(new_n532), .A3(new_n702), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n755), .B1(new_n756), .B2(KEYINPUT31), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n748), .A2(new_n751), .A3(new_n746), .ZN(new_n758));
  AND3_X1   g0558(.A1(new_n758), .A2(KEYINPUT31), .A3(new_n701), .ZN(new_n759));
  OAI21_X1  g0559(.A(G330), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT29), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n684), .A2(new_n761), .A3(new_n702), .ZN(new_n762));
  AND3_X1   g0562(.A1(new_n742), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n732), .B1(new_n763), .B2(G1), .ZN(G364));
  AOI21_X1  g0564(.A(new_n252), .B1(new_n695), .B2(G45), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n727), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n288), .A2(new_n352), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n427), .A2(G200), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n288), .A2(G190), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n513), .A2(G179), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI22_X1  g0575(.A1(G58), .A2(new_n771), .B1(new_n775), .B2(G107), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n772), .A2(new_n769), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n776), .B1(new_n345), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n768), .A2(new_n773), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n388), .B(new_n779), .C1(G87), .C2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G179), .A2(G200), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n772), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G159), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n784), .A2(KEYINPUT32), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(KEYINPUT32), .B1(new_n784), .B2(new_n785), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n288), .A2(new_n427), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n788), .A2(new_n352), .A3(G200), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n787), .B1(new_n209), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n788), .A2(G200), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n352), .ZN(new_n792));
  AOI211_X1 g0592(.A(new_n786), .B(new_n790), .C1(G50), .C2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n288), .B1(new_n783), .B2(G190), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n782), .B(new_n793), .C1(new_n265), .C2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G311), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n778), .A2(new_n796), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n342), .B(new_n797), .C1(G326), .C2(new_n792), .ZN(new_n798));
  INV_X1    g0598(.A(new_n784), .ZN(new_n799));
  AOI22_X1  g0599(.A1(G322), .A2(new_n771), .B1(new_n799), .B2(G329), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n781), .A2(G303), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(G283), .B2(new_n775), .ZN(new_n803));
  INV_X1    g0603(.A(new_n794), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(G294), .ZN(new_n805));
  INV_X1    g0605(.A(new_n789), .ZN(new_n806));
  INV_X1    g0606(.A(G317), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(KEYINPUT33), .ZN(new_n808));
  OR2_X1    g0608(.A1(new_n807), .A2(KEYINPUT33), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n806), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n798), .A2(new_n803), .A3(new_n805), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n795), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n229), .B1(G20), .B2(new_n454), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n247), .A2(G45), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n726), .A2(new_n342), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n814), .B(new_n815), .C1(G45), .C2(new_n233), .ZN(new_n816));
  NAND3_X1  g0616(.A1(G355), .A2(new_n342), .A3(new_n225), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n816), .B(new_n817), .C1(G116), .C2(new_n225), .ZN(new_n818));
  NOR2_X1   g0618(.A1(G13), .A2(G33), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT99), .Z(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(G20), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(new_n813), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n812), .A2(new_n813), .B1(new_n818), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n718), .A2(new_n720), .ZN(new_n825));
  INV_X1    g0625(.A(new_n822), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n767), .B(new_n824), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n721), .A2(new_n767), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n825), .A2(G330), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(G396));
  NAND2_X1  g0630(.A1(new_n684), .A2(new_n702), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n457), .A2(new_n701), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n455), .A2(new_n458), .ZN(new_n834));
  INV_X1    g0634(.A(new_n459), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NOR4_X1   g0636(.A1(new_n455), .A2(new_n458), .A3(new_n459), .A4(new_n832), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n466), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n831), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n838), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n684), .A2(new_n702), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  OR2_X1    g0642(.A1(new_n842), .A2(new_n760), .ZN(new_n843));
  INV_X1    g0643(.A(new_n767), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n842), .A2(new_n760), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  AOI22_X1  g0646(.A1(G137), .A2(new_n792), .B1(new_n806), .B2(G150), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT102), .ZN(new_n848));
  INV_X1    g0648(.A(G143), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n848), .B1(new_n849), .B2(new_n770), .C1(new_n785), .C2(new_n778), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(KEYINPUT34), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n775), .A2(G68), .ZN(new_n852));
  INV_X1    g0652(.A(G132), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n342), .B1(new_n784), .B2(new_n853), .C1(new_n202), .C2(new_n780), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(G58), .B2(new_n804), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n851), .A2(new_n852), .A3(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n774), .A2(new_n480), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n342), .B1(new_n781), .B2(G107), .ZN(new_n858));
  INV_X1    g0658(.A(new_n792), .ZN(new_n859));
  INV_X1    g0659(.A(G303), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n858), .B1(new_n796), .B2(new_n784), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n770), .A2(new_n493), .B1(new_n794), .B2(new_n265), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n861), .B1(KEYINPUT101), .B2(new_n862), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n806), .A2(G283), .B1(new_n777), .B2(G116), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n864), .B(KEYINPUT100), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n863), .B(new_n865), .C1(KEYINPUT101), .C2(new_n862), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n856), .B1(new_n857), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n813), .A2(new_n819), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n867), .A2(new_n813), .B1(new_n345), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n840), .B2(new_n821), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n846), .B1(new_n844), .B2(new_n870), .ZN(G384));
  INV_X1    g0671(.A(KEYINPUT38), .ZN(new_n872));
  INV_X1    g0672(.A(new_n699), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n297), .B1(new_n411), .B2(new_n412), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n873), .B1(new_n874), .B2(new_n420), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(new_n690), .B2(new_n418), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n426), .B(new_n430), .C1(new_n874), .C2(new_n420), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n877), .A2(new_n403), .A3(new_n875), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n878), .A2(KEYINPUT37), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT108), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n406), .A2(new_n415), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT37), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n877), .A2(new_n882), .A3(new_n875), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n880), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n877), .A2(new_n882), .A3(new_n875), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n885), .A2(KEYINPUT108), .A3(new_n416), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n879), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n872), .B1(new_n876), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(KEYINPUT111), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT105), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n890), .A2(KEYINPUT16), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(new_n409), .B2(new_n410), .ZN(new_n892));
  INV_X1    g0692(.A(new_n891), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n387), .A2(new_n392), .A3(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n892), .A2(new_n295), .A3(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT106), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n895), .A2(new_n896), .A3(new_n368), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n896), .B1(new_n895), .B2(new_n368), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n435), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n873), .B(new_n899), .C1(new_n417), .C2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT107), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n873), .B1(new_n426), .B2(new_n430), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n899), .A2(new_n904), .B1(new_n406), .B2(new_n415), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n902), .B1(new_n905), .B2(new_n882), .ZN(new_n906));
  NOR3_X1   g0706(.A1(new_n897), .A2(new_n903), .A3(new_n898), .ZN(new_n907));
  OAI211_X1 g0707(.A(KEYINPUT107), .B(KEYINPUT37), .C1(new_n881), .C2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NOR3_X1   g0709(.A1(new_n881), .A2(new_n880), .A3(new_n883), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT108), .B1(new_n885), .B2(new_n416), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g0712(.A(KEYINPUT38), .B(new_n901), .C1(new_n909), .C2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT111), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n914), .B(new_n872), .C1(new_n876), .C2(new_n887), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n889), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n754), .A2(KEYINPUT31), .A3(new_n701), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n756), .A2(KEYINPUT31), .ZN(new_n918));
  INV_X1    g0718(.A(new_n755), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AND3_X1   g0720(.A1(new_n281), .A2(new_n285), .A3(new_n286), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n314), .A2(new_n321), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n316), .A2(new_n702), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(new_n319), .B2(new_n320), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n922), .A2(new_n923), .B1(new_n308), .B2(new_n924), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n920), .A2(new_n925), .A3(new_n838), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n916), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(KEYINPUT40), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT109), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n913), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n901), .B1(new_n909), .B2(new_n912), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n872), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n906), .B(new_n908), .C1(new_n911), .C2(new_n910), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n933), .A2(KEYINPUT109), .A3(KEYINPUT38), .A4(new_n901), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n930), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT40), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n935), .A2(new_n926), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n928), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n920), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n468), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n938), .B(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(G330), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n690), .A2(new_n873), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  AND3_X1   g0744(.A1(new_n930), .A2(new_n932), .A3(new_n934), .ZN(new_n945));
  INV_X1    g0745(.A(new_n925), .ZN(new_n946));
  AOI211_X1 g0746(.A(new_n701), .B(new_n838), .C1(new_n672), .C2(new_n683), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n460), .A2(new_n702), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT104), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n946), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n944), .B1(new_n945), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(KEYINPUT110), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT39), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n916), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n308), .A2(new_n701), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n930), .A2(new_n932), .A3(KEYINPUT39), .A4(new_n934), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n949), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n925), .B1(new_n841), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n935), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT110), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n960), .A2(new_n961), .A3(new_n944), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n952), .A2(new_n957), .A3(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n942), .B(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n468), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n965), .B1(new_n742), .B2(new_n762), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n692), .A2(new_n464), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n964), .B(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n252), .B2(new_n695), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT35), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n231), .B1(new_n577), .B2(new_n971), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n972), .B(G116), .C1(new_n971), .C2(new_n577), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT36), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n379), .A2(G77), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n233), .A2(new_n975), .B1(G50), .B2(new_n209), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n976), .A2(G1), .A3(new_n694), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT103), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n970), .A2(new_n974), .A3(new_n978), .ZN(G367));
  NAND2_X1  g0779(.A1(new_n657), .A2(new_n701), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT112), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n678), .B1(new_n579), .B2(new_n702), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(KEYINPUT42), .B1(new_n984), .B2(new_n710), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n657), .B1(new_n983), .B2(new_n713), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n986), .A2(new_n701), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT42), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n983), .A2(new_n709), .A3(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n985), .A2(new_n987), .A3(new_n989), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n664), .A2(new_n702), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n991), .A2(new_n555), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(new_n673), .B2(new_n991), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT43), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n993), .A2(new_n994), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n990), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  AND2_X1   g0797(.A1(new_n985), .A2(new_n989), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n998), .A2(new_n994), .A3(new_n993), .A4(new_n987), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n722), .B2(new_n984), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n984), .A2(new_n722), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n997), .A2(new_n1002), .A3(new_n999), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT113), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n727), .B(KEYINPUT41), .Z(new_n1005));
  NAND3_X1  g0805(.A1(new_n710), .A2(new_n711), .A3(new_n983), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT45), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(KEYINPUT44), .B1(new_n712), .B2(new_n984), .ZN(new_n1009));
  AND3_X1   g0809(.A1(new_n712), .A2(KEYINPUT44), .A3(new_n984), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1008), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n723), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1008), .B(new_n722), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n710), .B1(new_n715), .B2(new_n707), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(new_n721), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1012), .A2(new_n763), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1005), .B1(new_n1016), .B2(new_n763), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1001), .B(new_n1004), .C1(new_n1017), .C2(new_n766), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n993), .A2(new_n822), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n388), .B1(new_n789), .B2(new_n493), .ZN(new_n1020));
  INV_X1    g0820(.A(G283), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n778), .A2(new_n1021), .B1(new_n265), .B2(new_n774), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n1020), .B(new_n1022), .C1(G317), .C2(new_n799), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n781), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT46), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n780), .B2(new_n213), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1024), .B(new_n1026), .C1(new_n474), .C2(new_n794), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(G311), .B2(new_n792), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1023), .B(new_n1028), .C1(new_n860), .C2(new_n770), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n859), .A2(new_n849), .B1(new_n785), .B2(new_n789), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G58), .B2(new_n781), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n804), .A2(G68), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n774), .A2(new_n345), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(KEYINPUT114), .B(G137), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n770), .A2(new_n324), .B1(new_n784), .B2(new_n1034), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n1033), .B(new_n1035), .C1(G50), .C2(new_n777), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1031), .A2(new_n342), .A3(new_n1032), .A4(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1029), .A2(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT47), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n844), .B1(new_n1039), .B2(new_n813), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n243), .A2(new_n815), .B1(new_n726), .B2(new_n533), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n823), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1019), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1018), .A2(new_n1043), .ZN(G387));
  OR2_X1    g0844(.A1(new_n1015), .A2(new_n763), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1015), .A2(new_n763), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1045), .A2(new_n727), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1015), .A2(new_n766), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n794), .A2(new_n439), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n342), .B1(new_n859), .B2(new_n785), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(G97), .C2(new_n775), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n771), .A2(G50), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n361), .A2(new_n806), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n778), .A2(new_n209), .B1(new_n784), .B2(new_n324), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n780), .A2(new_n345), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .A4(new_n1056), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n792), .A2(G322), .B1(G303), .B2(new_n777), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1058), .B1(new_n796), .B2(new_n789), .C1(new_n807), .C2(new_n770), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT48), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1060), .B1(new_n1021), .B2(new_n794), .C1(new_n493), .C2(new_n780), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT116), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(KEYINPUT115), .B(KEYINPUT49), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n342), .B1(new_n799), .B2(G326), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n774), .A2(new_n213), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1057), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n729), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(G68), .B2(G77), .ZN(new_n1072));
  OR3_X1    g0872(.A1(new_n360), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1073));
  OAI21_X1  g0873(.A(KEYINPUT50), .B1(new_n360), .B2(G50), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1072), .A2(new_n501), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n815), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n239), .B2(G45), .ZN(new_n1077));
  NOR3_X1   g0877(.A1(new_n729), .A2(new_n726), .A3(new_n388), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1075), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(G107), .B2(new_n225), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n1070), .A2(new_n813), .B1(new_n823), .B2(new_n1080), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1081), .B(new_n767), .C1(new_n715), .C2(new_n826), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1047), .A2(new_n1048), .A3(new_n1082), .ZN(G393));
  NAND3_X1  g0883(.A1(new_n1012), .A2(new_n766), .A3(new_n1013), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n823), .B1(new_n265), .B2(new_n225), .C1(new_n250), .C2(new_n1076), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n792), .A2(G150), .B1(new_n771), .B2(G159), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT51), .Z(new_n1087));
  NOR2_X1   g0887(.A1(new_n778), .A2(new_n360), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n794), .A2(new_n345), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n780), .A2(new_n209), .B1(new_n784), .B2(new_n849), .ZN(new_n1090));
  NOR3_X1   g0890(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n388), .B(new_n857), .C1(G50), .C2(new_n806), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1087), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n792), .A2(G317), .B1(new_n771), .B2(G311), .ZN(new_n1094));
  XOR2_X1   g0894(.A(new_n1094), .B(KEYINPUT52), .Z(new_n1095));
  AOI22_X1  g0895(.A1(G283), .A2(new_n781), .B1(new_n799), .B2(G322), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n789), .A2(new_n860), .B1(new_n774), .B2(new_n474), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n342), .B(new_n1097), .C1(G116), .C2(new_n804), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1095), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n778), .A2(new_n493), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1093), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n844), .B1(new_n1101), .B2(new_n813), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1085), .B(new_n1102), .C1(new_n983), .C2(new_n826), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1084), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n728), .B1(new_n1105), .B2(new_n1046), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1104), .B1(new_n1106), .B2(new_n1016), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(G390));
  NAND2_X1  g0908(.A1(new_n954), .A2(new_n956), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n955), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n950), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n740), .A2(new_n840), .A3(new_n702), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n948), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n946), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1115), .A2(new_n916), .A3(new_n1110), .ZN(new_n1116));
  OAI211_X1 g0916(.A(G330), .B(new_n840), .C1(new_n757), .C2(new_n759), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1117), .A2(new_n925), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1112), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n939), .A2(G330), .A3(new_n840), .A4(new_n946), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n954), .A2(new_n956), .B1(new_n950), .B2(new_n1110), .ZN(new_n1121));
  AND3_X1   g0921(.A1(new_n1115), .A2(new_n916), .A3(new_n1110), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1120), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n765), .B1(new_n1119), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n868), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1125), .A2(new_n361), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n342), .B1(new_n789), .B2(new_n1034), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n792), .A2(G128), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n785), .B2(new_n794), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n1127), .B(new_n1129), .C1(G50), .C2(new_n775), .ZN(new_n1130));
  XOR2_X1   g0930(.A(KEYINPUT54), .B(G143), .Z(new_n1131));
  NAND2_X1  g0931(.A1(new_n777), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n853), .B2(new_n770), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT53), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1134), .B1(new_n780), .B2(new_n324), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n781), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1133), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(G125), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1130), .B(new_n1137), .C1(new_n1138), .C2(new_n784), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT118), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(G283), .A2(new_n792), .B1(new_n806), .B2(G107), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1141), .B1(new_n265), .B2(new_n778), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT119), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n852), .B1(new_n213), .B2(new_n770), .C1(new_n493), .C2(new_n784), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1089), .B(new_n1144), .C1(G87), .C2(new_n781), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1143), .A2(new_n1145), .A3(new_n388), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1140), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n844), .B1(new_n1147), .B2(new_n813), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n1126), .B(new_n1149), .C1(new_n1109), .C2(new_n820), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1124), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT117), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n468), .B(G330), .C1(new_n757), .C2(new_n917), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  NOR3_X1   g0954(.A1(new_n966), .A2(new_n1154), .A3(new_n967), .ZN(new_n1155));
  OAI211_X1 g0955(.A(G330), .B(new_n840), .C1(new_n757), .C2(new_n917), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n1156), .A2(new_n925), .ZN(new_n1157));
  NOR3_X1   g0957(.A1(new_n1157), .A2(new_n1118), .A3(new_n1114), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1117), .A2(new_n925), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1120), .A2(new_n1159), .B1(new_n841), .B2(new_n958), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1155), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n1119), .A2(new_n1123), .A3(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1161), .B1(new_n1119), .B2(new_n1123), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1152), .B1(new_n1164), .B2(new_n727), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1161), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1120), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(new_n1112), .B2(new_n1116), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1118), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(new_n1121), .A2(new_n1122), .A3(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1166), .B1(new_n1168), .B2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1119), .A2(new_n1123), .A3(new_n1161), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1171), .A2(new_n727), .A3(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1173), .A2(KEYINPUT117), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1151), .B1(new_n1165), .B2(new_n1174), .ZN(G378));
  AND3_X1   g0975(.A1(new_n935), .A2(new_n926), .A3(new_n936), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n936), .B1(new_n916), .B2(new_n926), .ZN(new_n1177));
  OAI21_X1  g0977(.A(G330), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n337), .A2(new_n699), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n358), .A2(new_n463), .A3(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1180), .B1(new_n358), .B2(new_n463), .ZN(new_n1183));
  OAI21_X1  g0983(.A(KEYINPUT55), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1183), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT55), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1185), .A2(new_n1186), .A3(new_n1181), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1184), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT56), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1184), .A2(new_n1187), .A3(KEYINPUT56), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1178), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1192), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n938), .A2(G330), .A3(new_n1194), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n1193), .A2(new_n963), .A3(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n963), .B1(new_n1195), .B2(new_n1193), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n766), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(G128), .A2(new_n771), .B1(new_n781), .B2(new_n1131), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT120), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n777), .A2(G137), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n859), .B2(new_n1138), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G150), .B2(new_n804), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1200), .B(new_n1203), .C1(new_n853), .C2(new_n789), .ZN(new_n1204));
  XOR2_X1   g1004(.A(new_n1204), .B(KEYINPUT59), .Z(new_n1205));
  AOI21_X1  g1005(.A(G41), .B1(new_n799), .B2(G124), .ZN(new_n1206));
  AOI21_X1  g1006(.A(G33), .B1(new_n775), .B2(G159), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1032), .B1(new_n265), .B2(new_n789), .C1(new_n859), .C2(new_n213), .ZN(new_n1209));
  NOR4_X1   g1009(.A1(new_n1209), .A2(G41), .A3(new_n342), .A4(new_n1055), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n778), .A2(new_n439), .B1(new_n217), .B2(new_n774), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(G107), .B2(new_n771), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1210), .B(new_n1212), .C1(new_n1021), .C2(new_n784), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT58), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n202), .B1(new_n260), .B2(G41), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1208), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n844), .B1(new_n1216), .B2(new_n813), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(G50), .B2(new_n1125), .C1(new_n1192), .C2(new_n821), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1198), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n963), .A2(new_n1193), .A3(new_n1195), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n957), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n961), .B1(new_n960), .B2(new_n944), .ZN(new_n1223));
  AOI211_X1 g1023(.A(KEYINPUT110), .B(new_n943), .C1(new_n959), .C2(new_n935), .ZN(new_n1224));
  NOR3_X1   g1024(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1194), .B1(new_n938), .B2(G330), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n716), .B(new_n1192), .C1(new_n928), .C2(new_n937), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1225), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n1221), .A2(new_n1228), .B1(new_n1171), .B2(new_n1155), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n727), .B1(new_n1229), .B2(KEYINPUT57), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n968), .A2(new_n1153), .ZN(new_n1231));
  OAI21_X1  g1031(.A(KEYINPUT57), .B1(new_n1163), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT121), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1228), .A2(KEYINPUT121), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1232), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1220), .B1(new_n1230), .B2(new_n1236), .ZN(G375));
  NOR2_X1   g1037(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1238), .A2(new_n765), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n792), .A2(G132), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n806), .A2(new_n1131), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n804), .A2(G50), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1240), .A2(new_n1241), .A3(new_n342), .A4(new_n1242), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(G159), .A2(new_n781), .B1(new_n799), .B2(G128), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n1244), .B1(new_n324), .B2(new_n778), .C1(new_n770), .C2(new_n1034), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1243), .B(new_n1245), .C1(G58), .C2(new_n775), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(G283), .A2(new_n771), .B1(new_n781), .B2(G97), .ZN(new_n1247));
  OAI221_X1 g1047(.A(new_n1247), .B1(new_n474), .B2(new_n778), .C1(new_n860), .C2(new_n784), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1033), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n1249), .B1(new_n213), .B2(new_n789), .C1(new_n859), .C2(new_n493), .ZN(new_n1250));
  NOR4_X1   g1050(.A1(new_n1248), .A2(new_n1250), .A3(new_n342), .A4(new_n1049), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n813), .B1(new_n1246), .B2(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(G68), .B2(new_n1125), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(new_n925), .B2(new_n819), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1239), .B1(new_n767), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1238), .A2(new_n1231), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(new_n1005), .B(KEYINPUT122), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1256), .A2(new_n1161), .A3(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1255), .A2(new_n1258), .ZN(G381));
  OAI22_X1  g1059(.A1(new_n1196), .A2(new_n1197), .B1(new_n1231), .B2(new_n1163), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT57), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n728), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1261), .B1(new_n1171), .B2(new_n1155), .ZN(new_n1263));
  AOI21_X1  g1063(.A(KEYINPUT121), .B1(new_n1228), .B2(new_n1221), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1197), .A2(new_n1233), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1263), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1219), .B1(new_n1262), .B2(new_n1266), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1267), .B(KEYINPUT123), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1173), .A2(new_n1151), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1018), .A2(new_n1107), .A3(new_n1043), .ZN(new_n1271));
  NOR3_X1   g1071(.A1(new_n1271), .A2(G384), .A3(G381), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(G393), .A2(G396), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1270), .A2(new_n1272), .A3(new_n1273), .ZN(G407));
  NAND2_X1  g1074(.A1(new_n700), .A2(G213), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(new_n1275), .B(KEYINPUT124), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1270), .A2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(G407), .A2(G213), .A3(new_n1278), .ZN(G409));
  INV_X1    g1079(.A(new_n1275), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1266), .A2(new_n1281), .A3(new_n727), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1282), .A2(G378), .A3(new_n1220), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1269), .ZN(new_n1284));
  OAI221_X1 g1084(.A(new_n1257), .B1(new_n1163), .B2(new_n1231), .C1(new_n1196), .C2(new_n1197), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n1218), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n765), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1284), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1280), .B1(new_n1283), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT60), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n728), .B1(new_n1256), .B2(new_n1290), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1291), .B(new_n1161), .C1(new_n1290), .C2(new_n1256), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(G384), .B(KEYINPUT125), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1292), .A2(new_n1293), .A3(new_n1255), .ZN(new_n1294));
  AND2_X1   g1094(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1295), .B1(new_n1292), .B2(new_n1255), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1294), .A2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1280), .A2(G2897), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  OAI211_X1 g1099(.A(G2897), .B(new_n1277), .C1(new_n1294), .C2(new_n1296), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(KEYINPUT126), .B1(new_n1289), .B2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1292), .A2(new_n1255), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1295), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1292), .A2(new_n1293), .A3(new_n1255), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1276), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  AOI22_X1  g1107(.A1(new_n1307), .A2(G2897), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT126), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n766), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1310), .A2(new_n1218), .A3(new_n1285), .ZN(new_n1311));
  AOI22_X1  g1111(.A1(new_n1267), .A2(G378), .B1(new_n1311), .B2(new_n1284), .ZN(new_n1312));
  OAI211_X1 g1112(.A(new_n1308), .B(new_n1309), .C1(new_n1312), .C2(new_n1280), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1302), .A2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT61), .ZN(new_n1315));
  XOR2_X1   g1115(.A(G393), .B(G396), .Z(new_n1316));
  INV_X1    g1116(.A(new_n1271), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1107), .B1(new_n1018), .B2(new_n1043), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1316), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1318), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1316), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1320), .A2(new_n1271), .A3(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1319), .A2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1151), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1174), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1173), .A2(KEYINPUT117), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1324), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1288), .B1(G375), .B2(new_n1327), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1328), .A2(new_n1275), .A3(new_n1297), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT63), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1323), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1312), .A2(new_n1277), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1332), .A2(KEYINPUT63), .A3(new_n1297), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1314), .A2(new_n1315), .A3(new_n1331), .A4(new_n1333), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1308), .B1(new_n1312), .B2(new_n1277), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT62), .ZN(new_n1336));
  NAND4_X1  g1136(.A1(new_n1328), .A2(new_n1336), .A3(new_n1275), .A4(new_n1297), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1335), .A2(new_n1337), .A3(new_n1315), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1336), .B1(new_n1332), .B2(new_n1297), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1323), .B1(new_n1338), .B2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1334), .A2(new_n1340), .ZN(G405));
  NAND2_X1  g1141(.A1(G375), .A2(new_n1284), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(new_n1283), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT127), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  INV_X1    g1145(.A(new_n1323), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1345), .A2(new_n1346), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1342), .A2(KEYINPUT127), .A3(new_n1283), .ZN(new_n1348));
  AND2_X1   g1148(.A1(new_n1348), .A2(new_n1297), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1323), .A2(new_n1343), .A3(new_n1344), .ZN(new_n1350));
  AND3_X1   g1150(.A1(new_n1347), .A2(new_n1349), .A3(new_n1350), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1349), .B1(new_n1347), .B2(new_n1350), .ZN(new_n1352));
  NOR2_X1   g1152(.A1(new_n1351), .A2(new_n1352), .ZN(G402));
endmodule


