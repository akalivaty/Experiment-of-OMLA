//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 0 1 1 0 0 1 1 1 1 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 1 1 0 0 0 0 1 0 1 0 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n753, new_n754, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989;
  INV_X1    g000(.A(KEYINPUT77), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G116), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT2), .B(G113), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  AND2_X1   g009(.A1(KEYINPUT64), .A2(G146), .ZN(new_n196));
  NOR2_X1   g010(.A1(KEYINPUT64), .A2(G146), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  NOR3_X1   g012(.A1(new_n196), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT1), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT69), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  OR2_X1    g015(.A1(KEYINPUT64), .A2(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT64), .A2(G146), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(G143), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT69), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(KEYINPUT1), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n201), .A2(G128), .A3(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n198), .A2(G146), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n196), .A2(new_n197), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n209), .B1(new_n210), .B2(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n207), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n204), .A2(new_n213), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n202), .A2(KEYINPUT65), .A3(G143), .A4(new_n203), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G146), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT66), .B1(new_n217), .B2(G143), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(new_n198), .A3(G146), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n200), .A2(G128), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n216), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n212), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G131), .ZN(new_n227));
  INV_X1    g041(.A(G137), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G134), .ZN(new_n229));
  INV_X1    g043(.A(G134), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G137), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n227), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n228), .A2(KEYINPUT11), .A3(G134), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(new_n231), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT11), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n235), .B1(new_n230), .B2(G137), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT67), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n229), .A2(new_n238), .A3(new_n235), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n234), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  XOR2_X1   g054(.A(KEYINPUT68), .B(G131), .Z(new_n241));
  AOI21_X1  g055(.A(new_n232), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n233), .A2(new_n231), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n238), .B1(new_n229), .B2(new_n235), .ZN(new_n244));
  AOI211_X1 g058(.A(KEYINPUT67), .B(KEYINPUT11), .C1(new_n228), .C2(G134), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n243), .B(new_n241), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n246), .B1(new_n227), .B2(new_n240), .ZN(new_n247));
  NAND2_X1  g061(.A1(KEYINPUT0), .A2(G128), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n216), .A2(new_n222), .A3(new_n249), .ZN(new_n250));
  OR2_X1    g064(.A1(KEYINPUT0), .A2(G128), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n211), .A2(new_n248), .A3(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n247), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT71), .ZN(new_n254));
  AOI22_X1  g068(.A1(new_n226), .A2(new_n242), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n247), .A2(new_n250), .A3(KEYINPUT71), .A4(new_n252), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n195), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n253), .A2(new_n254), .ZN(new_n258));
  INV_X1    g072(.A(new_n211), .ZN(new_n259));
  INV_X1    g073(.A(G128), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n204), .A2(KEYINPUT1), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n260), .B1(new_n261), .B2(KEYINPUT69), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n259), .B1(new_n262), .B2(new_n206), .ZN(new_n263));
  AOI211_X1 g077(.A(new_n221), .B(new_n223), .C1(new_n214), .C2(new_n215), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n242), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n258), .A2(new_n265), .A3(new_n195), .A4(new_n256), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT28), .B1(new_n257), .B2(new_n267), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n247), .A2(new_n250), .A3(new_n252), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n269), .A2(new_n194), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT28), .B1(new_n270), .B2(new_n265), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n273));
  INV_X1    g087(.A(G237), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(KEYINPUT72), .A2(G237), .ZN(new_n276));
  AOI21_X1  g090(.A(G953), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G210), .ZN(new_n278));
  XNOR2_X1  g092(.A(KEYINPUT26), .B(G101), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n278), .B(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(KEYINPUT73), .B(KEYINPUT27), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n280), .B(new_n281), .ZN(new_n282));
  AND2_X1   g096(.A1(new_n282), .A2(KEYINPUT29), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n268), .A2(KEYINPUT76), .A3(new_n272), .A4(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G902), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n258), .A2(new_n265), .A3(new_n256), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n194), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n266), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n271), .B1(new_n289), .B2(KEYINPUT28), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT76), .B1(new_n290), .B2(new_n283), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n187), .B1(new_n286), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n268), .A2(new_n272), .A3(new_n283), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT76), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n295), .A2(KEYINPUT77), .A3(new_n285), .A4(new_n284), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n221), .B1(new_n214), .B2(new_n215), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n207), .A2(new_n211), .B1(new_n297), .B2(new_n224), .ZN(new_n298));
  INV_X1    g112(.A(new_n242), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT70), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT70), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n242), .B(new_n301), .C1(new_n263), .C2(new_n264), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n300), .A2(new_n302), .A3(new_n253), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT30), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n255), .A2(KEYINPUT30), .A3(new_n256), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(new_n194), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n266), .ZN(new_n308));
  INV_X1    g122(.A(new_n282), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT29), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n269), .B1(new_n265), .B2(KEYINPUT70), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n195), .B1(new_n311), .B2(new_n302), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT28), .B1(new_n312), .B2(new_n267), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(new_n282), .A3(new_n272), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n292), .A2(new_n296), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G472), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n267), .A2(new_n309), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n307), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT74), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT74), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n307), .A2(new_n321), .A3(new_n318), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n320), .A2(KEYINPUT31), .A3(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT31), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n307), .A2(new_n324), .A3(new_n318), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n282), .B1(new_n313), .B2(new_n272), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(G472), .A2(G902), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(KEYINPUT32), .A3(new_n329), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n307), .A2(new_n321), .A3(new_n318), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n321), .B1(new_n307), .B2(new_n318), .ZN(new_n332));
  NOR3_X1   g146(.A1(new_n331), .A2(new_n332), .A3(new_n324), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n313), .A2(new_n272), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(new_n309), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n307), .A2(new_n324), .A3(new_n318), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n329), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT75), .B(KEYINPUT32), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n317), .A2(new_n330), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G217), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n343), .B1(G234), .B2(new_n285), .ZN(new_n344));
  INV_X1    g158(.A(G953), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(G221), .A3(G234), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(KEYINPUT79), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT22), .B(G137), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n347), .B(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n188), .A2(G128), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n260), .A2(KEYINPUT23), .A3(G119), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n188), .A2(G128), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n351), .B(new_n352), .C1(new_n353), .C2(KEYINPUT23), .ZN(new_n354));
  XNOR2_X1  g168(.A(G119), .B(G128), .ZN(new_n355));
  INV_X1    g169(.A(G110), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(KEYINPUT24), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT24), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G110), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  AOI22_X1  g174(.A1(new_n354), .A2(G110), .B1(new_n355), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G140), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G125), .ZN(new_n363));
  INV_X1    g177(.A(G125), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G140), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n363), .A2(new_n365), .A3(KEYINPUT16), .ZN(new_n366));
  OR3_X1    g180(.A1(new_n364), .A2(KEYINPUT16), .A3(G140), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n366), .A2(G146), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(G146), .B1(new_n366), .B2(new_n367), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n361), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT78), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n260), .A2(G119), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n351), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT24), .B(G110), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n375), .B1(new_n354), .B2(G110), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n366), .A2(new_n367), .A3(G146), .ZN(new_n377));
  XNOR2_X1  g191(.A(G125), .B(G140), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n210), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n376), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n370), .A2(new_n371), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n371), .B1(new_n370), .B2(new_n380), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n350), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n370), .A2(new_n380), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n349), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(KEYINPUT25), .B1(new_n386), .B2(new_n285), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT25), .ZN(new_n388));
  AOI211_X1 g202(.A(new_n388), .B(G902), .C1(new_n383), .C2(new_n385), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n344), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT80), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI211_X1 g206(.A(KEYINPUT80), .B(new_n344), .C1(new_n387), .C2(new_n389), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n344), .A2(G902), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n386), .A2(new_n394), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n392), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(KEYINPUT9), .B(G234), .ZN(new_n397));
  OAI21_X1  g211(.A(G221), .B1(new_n397), .B2(G902), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G469), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n400), .A2(new_n285), .ZN(new_n401));
  INV_X1    g215(.A(G104), .ZN(new_n402));
  OAI21_X1  g216(.A(KEYINPUT3), .B1(new_n402), .B2(G107), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT3), .ZN(new_n404));
  INV_X1    g218(.A(G107), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n404), .A2(new_n405), .A3(G104), .ZN(new_n406));
  INV_X1    g220(.A(G101), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n402), .A2(G107), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n403), .A2(new_n406), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n402), .A2(G107), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n405), .A2(G104), .ZN(new_n411));
  OAI21_X1  g225(.A(G101), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n260), .B1(new_n209), .B2(KEYINPUT1), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n297), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n414), .B1(new_n416), .B2(new_n264), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT10), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n413), .A2(KEYINPUT82), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT82), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n409), .A2(new_n412), .A3(new_n421), .ZN(new_n422));
  AND2_X1   g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n423), .B(KEYINPUT10), .C1(new_n263), .C2(new_n264), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n403), .A2(new_n406), .A3(new_n408), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT4), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n426), .A3(G101), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n425), .A2(G101), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(KEYINPUT4), .A3(new_n409), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n250), .A2(new_n252), .A3(new_n427), .A4(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n419), .A2(new_n424), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n247), .ZN(new_n432));
  INV_X1    g246(.A(new_n247), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n419), .A2(new_n433), .A3(new_n424), .A4(new_n430), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  XNOR2_X1  g249(.A(G110), .B(G140), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n436), .B(KEYINPUT81), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n345), .A2(G227), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n437), .B(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n435), .A2(new_n440), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n434), .A2(new_n439), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT83), .ZN(new_n443));
  AOI21_X1  g257(.A(KEYINPUT12), .B1(new_n247), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n420), .A2(new_n422), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n225), .B1(new_n297), .B2(new_n415), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n298), .A2(new_n445), .B1(new_n446), .B2(new_n414), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n444), .B1(new_n447), .B2(new_n433), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n212), .A2(new_n225), .A3(new_n445), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n417), .ZN(new_n450));
  INV_X1    g264(.A(new_n444), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n450), .A2(new_n247), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n442), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(G902), .B1(new_n441), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n401), .B1(new_n455), .B2(new_n400), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n434), .A2(new_n439), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT85), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n434), .A2(KEYINPUT85), .A3(new_n439), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n432), .A3(new_n460), .ZN(new_n461));
  AOI211_X1 g275(.A(new_n433), .B(new_n444), .C1(new_n449), .C2(new_n417), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n451), .B1(new_n450), .B2(new_n247), .ZN(new_n463));
  OAI211_X1 g277(.A(KEYINPUT84), .B(new_n434), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n440), .ZN(new_n465));
  AOI21_X1  g279(.A(KEYINPUT84), .B1(new_n453), .B2(new_n434), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n461), .B(G469), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n399), .B1(new_n456), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n190), .A2(G122), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n190), .A2(G122), .ZN(new_n471));
  OAI21_X1  g285(.A(G107), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(G122), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(G116), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n474), .A2(new_n469), .A3(new_n405), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n198), .A2(G128), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n260), .A2(G143), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(new_n478), .A3(new_n230), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT13), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n198), .A2(KEYINPUT13), .A3(G128), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n481), .A2(new_n482), .A3(new_n478), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n476), .B(new_n479), .C1(new_n483), .C2(new_n230), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n477), .A2(new_n478), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(G134), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n486), .A2(new_n479), .B1(KEYINPUT94), .B2(new_n475), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n487), .B1(KEYINPUT94), .B2(new_n475), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n469), .B1(new_n471), .B2(KEYINPUT14), .ZN(new_n489));
  OR2_X1    g303(.A1(new_n489), .A2(KEYINPUT95), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n469), .A2(KEYINPUT14), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n491), .B1(new_n489), .B2(KEYINPUT95), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n405), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n484), .B1(new_n488), .B2(new_n493), .ZN(new_n494));
  OR3_X1    g308(.A1(new_n397), .A2(new_n343), .A3(G953), .ZN(new_n495));
  OR2_X1    g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n495), .ZN(new_n497));
  AOI21_X1  g311(.A(G902), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G478), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n499), .A2(KEYINPUT15), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  AND2_X1   g315(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n498), .A2(new_n501), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(G113), .B(G122), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n505), .B(new_n402), .ZN(new_n506));
  INV_X1    g320(.A(new_n276), .ZN(new_n507));
  NOR2_X1   g321(.A1(KEYINPUT72), .A2(G237), .ZN(new_n508));
  OAI211_X1 g322(.A(G214), .B(new_n345), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(KEYINPUT88), .A3(new_n198), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n198), .A2(KEYINPUT88), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n277), .A2(G214), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n510), .A2(new_n241), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT92), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n510), .A2(new_n512), .ZN(new_n515));
  INV_X1    g329(.A(new_n241), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT92), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n510), .A2(new_n512), .A3(new_n518), .A4(new_n241), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n514), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n378), .B(KEYINPUT19), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n368), .B1(new_n521), .B2(new_n210), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(KEYINPUT18), .A2(G131), .ZN(new_n524));
  XOR2_X1   g338(.A(new_n524), .B(KEYINPUT90), .Z(new_n525));
  NAND3_X1  g339(.A1(new_n510), .A2(new_n512), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT91), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n510), .A2(new_n512), .A3(KEYINPUT91), .A4(new_n525), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n524), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n378), .A2(new_n217), .ZN(new_n532));
  OR2_X1    g346(.A1(new_n532), .A2(KEYINPUT89), .ZN(new_n533));
  AOI22_X1  g347(.A1(new_n532), .A2(KEYINPUT89), .B1(new_n210), .B2(new_n378), .ZN(new_n534));
  AOI22_X1  g348(.A1(new_n515), .A2(new_n531), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n506), .B1(new_n523), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT17), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n514), .A2(new_n517), .A3(new_n538), .A4(new_n519), .ZN(new_n539));
  OR2_X1    g353(.A1(new_n368), .A2(new_n369), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n241), .B1(new_n510), .B2(new_n512), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n540), .B1(KEYINPUT17), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(new_n506), .A3(new_n536), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT93), .ZN(new_n545));
  AOI22_X1  g359(.A1(new_n539), .A2(new_n542), .B1(new_n530), .B2(new_n535), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT93), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(new_n547), .A3(new_n506), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n537), .B1(new_n545), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(G475), .A2(G902), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(KEYINPUT20), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n537), .ZN(new_n553));
  AND4_X1   g367(.A1(new_n547), .A2(new_n543), .A3(new_n506), .A4(new_n536), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n547), .B1(new_n546), .B2(new_n506), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT20), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n556), .A2(new_n557), .A3(new_n550), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n552), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(G234), .A2(G237), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n560), .A2(G902), .A3(G953), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(KEYINPUT96), .ZN(new_n562));
  XOR2_X1   g376(.A(KEYINPUT21), .B(G898), .Z(new_n563));
  NOR2_X1   g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(G952), .ZN(new_n565));
  AOI211_X1 g379(.A(G953), .B(new_n565), .C1(G234), .C2(G237), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(KEYINPUT97), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n554), .A2(new_n555), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n546), .A2(new_n506), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n285), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(G475), .ZN(new_n572));
  AND4_X1   g386(.A1(new_n504), .A2(new_n559), .A3(new_n568), .A4(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(G214), .B1(G237), .B2(G902), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n263), .A2(G125), .A3(new_n264), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n345), .A2(G224), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n364), .B1(new_n250), .B2(new_n252), .ZN(new_n579));
  NOR3_X1   g393(.A1(new_n576), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n298), .A2(new_n364), .ZN(new_n581));
  INV_X1    g395(.A(new_n579), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n577), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n192), .A2(new_n193), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n189), .A2(new_n191), .A3(KEYINPUT5), .ZN(new_n585));
  OR3_X1    g399(.A1(new_n190), .A2(KEYINPUT5), .A3(G119), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(new_n586), .A3(G113), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT86), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n584), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n585), .A2(new_n586), .A3(KEYINPUT86), .A4(G113), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n589), .A2(new_n420), .A3(new_n422), .A4(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n429), .A2(new_n194), .A3(new_n427), .ZN(new_n592));
  XNOR2_X1  g406(.A(G110), .B(G122), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n591), .A2(new_n592), .ZN(new_n595));
  INV_X1    g409(.A(new_n593), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n596), .A2(KEYINPUT87), .ZN(new_n597));
  AOI22_X1  g411(.A1(new_n594), .A2(KEYINPUT6), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n595), .A2(KEYINPUT6), .A3(new_n597), .ZN(new_n599));
  OAI22_X1  g413(.A1(new_n580), .A2(new_n583), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n594), .ZN(new_n601));
  XOR2_X1   g415(.A(new_n593), .B(KEYINPUT8), .Z(new_n602));
  NAND2_X1  g416(.A1(new_n589), .A2(new_n590), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n413), .ZN(new_n604));
  INV_X1    g418(.A(new_n584), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n420), .A2(new_n605), .A3(new_n422), .A4(new_n587), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n602), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n601), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n578), .B1(new_n576), .B2(new_n579), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n581), .A2(new_n582), .A3(KEYINPUT7), .A4(new_n577), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT7), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n611), .B1(new_n576), .B2(new_n579), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n608), .A2(new_n609), .A3(new_n610), .A4(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n600), .A2(new_n613), .A3(new_n285), .ZN(new_n614));
  OAI21_X1  g428(.A(G210), .B1(G237), .B2(G902), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n600), .A2(new_n613), .A3(new_n285), .A4(new_n615), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n575), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AND3_X1   g433(.A1(new_n468), .A2(new_n573), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n342), .A2(new_n396), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G101), .ZN(G3));
  AOI21_X1  g436(.A(G902), .B1(new_n323), .B2(new_n327), .ZN(new_n623));
  INV_X1    g437(.A(G472), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n338), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n457), .B1(new_n452), .B2(new_n448), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n439), .B1(new_n432), .B2(new_n434), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n400), .B(new_n285), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n401), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n467), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n630), .A2(new_n396), .A3(new_n398), .ZN(new_n631));
  OAI21_X1  g445(.A(KEYINPUT98), .B1(new_n625), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n285), .B1(new_n333), .B2(new_n337), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(G472), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n630), .A2(new_n396), .A3(new_n398), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT98), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n634), .A2(new_n635), .A3(new_n636), .A4(new_n338), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n498), .A2(new_n499), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n499), .A2(new_n285), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n496), .A2(new_n497), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT33), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n642), .B1(new_n497), .B2(KEYINPUT99), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n641), .B(new_n643), .ZN(new_n644));
  OAI211_X1 g458(.A(new_n638), .B(new_n640), .C1(new_n644), .C2(new_n499), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n645), .B1(new_n559), .B2(new_n572), .ZN(new_n646));
  INV_X1    g460(.A(new_n568), .ZN(new_n647));
  AOI211_X1 g461(.A(new_n647), .B(new_n575), .C1(new_n617), .C2(new_n618), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n632), .A2(new_n637), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT100), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT34), .B(G104), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G6));
  INV_X1    g467(.A(new_n504), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n619), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n559), .A2(new_n572), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n655), .A2(new_n656), .A3(new_n647), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n632), .A2(new_n637), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT35), .B(G107), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G9));
  INV_X1    g474(.A(new_n625), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n381), .A2(new_n382), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT36), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n662), .A2(new_n663), .A3(new_n349), .ZN(new_n664));
  OAI22_X1  g478(.A1(new_n381), .A2(new_n382), .B1(KEYINPUT36), .B2(new_n350), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n666), .A2(KEYINPUT101), .A3(new_n394), .ZN(new_n667));
  AOI21_X1  g481(.A(KEYINPUT101), .B1(new_n666), .B2(new_n394), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n392), .A2(new_n669), .A3(new_n393), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n670), .A2(new_n619), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n661), .A2(new_n573), .A3(new_n468), .A4(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT37), .B(G110), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G12));
  NOR2_X1   g488(.A1(new_n656), .A2(new_n504), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n562), .A2(G900), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n676), .A2(new_n566), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT102), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n468), .A2(new_n675), .A3(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n342), .A2(new_n671), .A3(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT103), .B(G128), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G30));
  NAND2_X1  g497(.A1(new_n289), .A2(new_n309), .ZN(new_n684));
  OR2_X1    g498(.A1(new_n684), .A2(KEYINPUT104), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(KEYINPUT104), .ZN(new_n686));
  AND4_X1   g500(.A1(new_n320), .A2(new_n685), .A3(new_n322), .A4(new_n686), .ZN(new_n687));
  OAI21_X1  g501(.A(G472), .B1(new_n687), .B2(G902), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n341), .A2(new_n330), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT105), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n617), .A2(new_n618), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT38), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  AOI22_X1  g507(.A1(new_n552), .A2(new_n558), .B1(new_n571), .B2(G475), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n654), .A2(new_n574), .ZN(new_n695));
  NOR4_X1   g509(.A1(new_n693), .A2(new_n694), .A3(new_n670), .A4(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n630), .A2(new_n398), .ZN(new_n697));
  XOR2_X1   g511(.A(new_n678), .B(KEYINPUT39), .Z(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(KEYINPUT40), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n696), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n701), .A2(KEYINPUT40), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n690), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(new_n198), .ZN(G45));
  NAND2_X1  g520(.A1(new_n646), .A2(new_n679), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n707), .A2(new_n697), .ZN(new_n708));
  INV_X1    g522(.A(new_n329), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n709), .B1(new_n323), .B2(new_n327), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n330), .B1(new_n710), .B2(new_n339), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n295), .A2(new_n285), .A3(new_n284), .ZN(new_n712));
  AOI22_X1  g526(.A1(new_n712), .A2(new_n187), .B1(new_n314), .B2(new_n310), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n624), .B1(new_n713), .B2(new_n296), .ZN(new_n714));
  OAI211_X1 g528(.A(new_n671), .B(new_n708), .C1(new_n711), .C2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G146), .ZN(G48));
  AOI22_X1  g530(.A1(new_n440), .A2(new_n435), .B1(new_n442), .B2(new_n453), .ZN(new_n717));
  OAI21_X1  g531(.A(G469), .B1(new_n717), .B2(G902), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n718), .A2(new_n398), .A3(new_n628), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT106), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n718), .A2(KEYINPUT106), .A3(new_n398), .A4(new_n628), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n342), .A2(new_n396), .A3(new_n649), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT41), .B(G113), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G15));
  INV_X1    g540(.A(new_n396), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n339), .B1(new_n328), .B2(new_n329), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT32), .ZN(new_n729));
  AOI211_X1 g543(.A(new_n729), .B(new_n709), .C1(new_n323), .C2(new_n327), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n727), .B1(new_n731), .B2(new_n317), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT107), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n732), .A2(new_n733), .A3(new_n657), .A4(new_n723), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n342), .A2(new_n396), .A3(new_n657), .A4(new_n723), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(KEYINPUT107), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G116), .ZN(G18));
  AND3_X1   g552(.A1(new_n721), .A2(new_n619), .A3(new_n722), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n342), .A2(new_n739), .A3(new_n573), .A4(new_n670), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G119), .ZN(G21));
  INV_X1    g555(.A(KEYINPUT109), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n742), .B1(new_n655), .B2(new_n694), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n656), .A2(KEYINPUT109), .A3(new_n654), .A4(new_n619), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n647), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n290), .A2(new_n282), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(new_n325), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n709), .B1(new_n323), .B2(new_n747), .ZN(new_n748));
  XOR2_X1   g562(.A(KEYINPUT108), .B(G472), .Z(new_n749));
  AOI21_X1  g563(.A(new_n748), .B1(new_n633), .B2(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n745), .A2(new_n396), .A3(new_n723), .A4(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G122), .ZN(G24));
  INV_X1    g566(.A(new_n707), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n739), .A2(new_n670), .A3(new_n753), .A4(new_n750), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G125), .ZN(G27));
  NAND2_X1  g569(.A1(new_n338), .A2(new_n729), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n317), .A2(new_n330), .A3(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n691), .A2(new_n575), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n697), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n757), .A2(new_n396), .A3(new_n753), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(KEYINPUT42), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n707), .A2(KEYINPUT42), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n342), .A2(new_n396), .A3(new_n760), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(new_n227), .ZN(G33));
  INV_X1    g580(.A(new_n675), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(new_n678), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n342), .A2(new_n768), .A3(new_n396), .A4(new_n760), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G134), .ZN(G36));
  OAI21_X1  g584(.A(new_n461), .B1(new_n465), .B2(new_n466), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT45), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n400), .B1(new_n771), .B2(new_n772), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n775), .A2(new_n401), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n776), .A2(KEYINPUT46), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(KEYINPUT46), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(new_n628), .A3(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(new_n398), .A3(new_n698), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(KEYINPUT110), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n656), .A2(new_n645), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT111), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n782), .B1(new_n783), .B2(KEYINPUT43), .ZN(new_n784));
  XNOR2_X1  g598(.A(KEYINPUT111), .B(KEYINPUT43), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n784), .B1(new_n782), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n786), .A2(new_n625), .A3(new_n670), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT44), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n758), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n789), .B1(new_n788), .B2(new_n787), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n781), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G137), .ZN(G39));
  NAND2_X1  g606(.A1(new_n779), .A2(new_n398), .ZN(new_n793));
  XOR2_X1   g607(.A(new_n793), .B(KEYINPUT47), .Z(new_n794));
  NOR4_X1   g608(.A1(new_n342), .A2(new_n396), .A3(new_n707), .A4(new_n759), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G140), .ZN(G42));
  NAND3_X1  g611(.A1(new_n724), .A2(new_n740), .A3(new_n751), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n798), .B1(new_n734), .B2(new_n736), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT119), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n799), .B(new_n800), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n681), .A2(new_n754), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n743), .A2(new_n744), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n697), .A2(new_n670), .A3(new_n678), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n689), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n715), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n802), .A2(new_n806), .A3(KEYINPUT117), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n681), .A2(new_n754), .A3(new_n715), .A4(new_n805), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT117), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT52), .B1(new_n807), .B2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n812), .B1(new_n802), .B2(new_n806), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT113), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n646), .A2(new_n648), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n815), .B1(new_n646), .B2(new_n648), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n632), .A2(new_n637), .A3(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT114), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n819), .A2(new_n820), .A3(new_n621), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n820), .B1(new_n819), .B2(new_n621), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n658), .A2(new_n672), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n750), .A2(new_n760), .A3(new_n753), .A4(new_n670), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n502), .A2(new_n503), .A3(new_n678), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n758), .A2(new_n694), .A3(KEYINPUT115), .A4(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n826), .A2(new_n617), .A3(new_n574), .A4(new_n618), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n828), .B1(new_n656), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n697), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n342), .A2(new_n670), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n769), .A2(new_n825), .A3(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n765), .A2(new_n833), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n824), .A2(KEYINPUT53), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n801), .A2(new_n814), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT118), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n807), .A2(KEYINPUT52), .A3(new_n810), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n838), .B1(new_n839), .B2(new_n811), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT117), .B1(new_n802), .B2(new_n806), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n808), .A2(new_n809), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n812), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n807), .A2(new_n810), .A3(KEYINPUT52), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n843), .A2(KEYINPUT118), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n342), .A2(new_n396), .A3(new_n760), .ZN(new_n848));
  AOI22_X1  g662(.A1(new_n848), .A2(new_n763), .B1(new_n761), .B2(KEYINPUT42), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n724), .A2(new_n740), .A3(new_n751), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n769), .A2(new_n825), .A3(new_n832), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n737), .A2(new_n849), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n819), .A2(new_n621), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT114), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n819), .A2(new_n820), .A3(new_n621), .ZN(new_n855));
  INV_X1    g669(.A(new_n823), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n847), .B1(new_n852), .B2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n824), .A2(KEYINPUT116), .A3(new_n799), .A4(new_n834), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n846), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n837), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n858), .A2(new_n859), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n866), .B1(new_n840), .B2(new_n845), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n814), .A2(new_n862), .ZN(new_n868));
  OAI22_X1  g682(.A1(new_n867), .A2(new_n862), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n865), .B1(new_n864), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n786), .A2(new_n566), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n872), .A2(new_n396), .A3(new_n750), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n718), .A2(new_n628), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT112), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(new_n398), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n758), .B(new_n873), .C1(new_n794), .C2(new_n876), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n871), .A2(new_n574), .A3(new_n692), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n878), .A2(new_n396), .A3(new_n723), .A4(new_n750), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT50), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n723), .A2(new_n758), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT120), .ZN(new_n882));
  AND4_X1   g696(.A1(new_n670), .A2(new_n882), .A3(new_n750), .A4(new_n872), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n882), .A2(new_n396), .A3(new_n566), .A4(new_n690), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n694), .A2(new_n645), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n877), .B(new_n884), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT51), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n887), .A2(new_n888), .ZN(new_n890));
  AND4_X1   g704(.A1(new_n396), .A2(new_n882), .A3(new_n757), .A4(new_n872), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT48), .ZN(new_n892));
  INV_X1    g706(.A(new_n646), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n885), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n873), .A2(new_n739), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n895), .A2(G952), .A3(new_n345), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n892), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n889), .A2(new_n890), .A3(new_n897), .ZN(new_n898));
  OAI22_X1  g712(.A1(new_n870), .A2(new_n898), .B1(G952), .B2(G953), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n875), .B(KEYINPUT49), .Z(new_n900));
  AND4_X1   g714(.A1(new_n398), .A2(new_n693), .A3(new_n574), .A4(new_n782), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n900), .A2(new_n690), .A3(new_n396), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n899), .A2(new_n902), .ZN(G75));
  NAND2_X1  g717(.A1(new_n565), .A2(G953), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT122), .Z(new_n905));
  AOI21_X1  g719(.A(KEYINPUT53), .B1(new_n846), .B2(new_n860), .ZN(new_n906));
  OAI211_X1 g720(.A(G210), .B(G902), .C1(new_n906), .C2(new_n837), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT56), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n598), .A2(new_n599), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n909), .B(KEYINPUT121), .Z(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT55), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n580), .A2(new_n583), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n911), .B(new_n912), .Z(new_n913));
  AND3_X1   g727(.A1(new_n907), .A2(new_n908), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n913), .B1(new_n907), .B2(new_n908), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n905), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT123), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI211_X1 g732(.A(KEYINPUT123), .B(new_n905), .C1(new_n914), .C2(new_n915), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(G51));
  INV_X1    g734(.A(new_n905), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n836), .B1(new_n867), .B2(KEYINPUT53), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n922), .A2(G902), .A3(new_n775), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT124), .Z(new_n924));
  XNOR2_X1  g738(.A(new_n863), .B(KEYINPUT54), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n401), .B(KEYINPUT57), .Z(new_n926));
  OAI22_X1  g740(.A1(new_n925), .A2(new_n926), .B1(new_n627), .B2(new_n626), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n921), .B1(new_n924), .B2(new_n927), .ZN(G54));
  NAND4_X1  g742(.A1(new_n922), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n929));
  OR2_X1    g743(.A1(new_n929), .A2(new_n556), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n556), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n921), .B1(new_n930), .B2(new_n931), .ZN(G60));
  XOR2_X1   g746(.A(new_n639), .B(KEYINPUT59), .Z(new_n933));
  NAND2_X1  g747(.A1(new_n644), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n905), .B1(new_n925), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n644), .B1(new_n870), .B2(new_n933), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n935), .A2(new_n936), .ZN(G63));
  NAND2_X1  g751(.A1(G217), .A2(G902), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT60), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n666), .B(new_n940), .C1(new_n906), .C2(new_n837), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n905), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n386), .B1(new_n922), .B2(new_n940), .ZN(new_n943));
  OAI21_X1  g757(.A(KEYINPUT126), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT125), .ZN(new_n945));
  AOI21_X1  g759(.A(KEYINPUT61), .B1(new_n941), .B2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n386), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n947), .B1(new_n863), .B2(new_n939), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT126), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n948), .A2(new_n949), .A3(new_n905), .A4(new_n941), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n944), .A2(new_n946), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n946), .B1(new_n944), .B2(new_n950), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n951), .A2(new_n952), .ZN(G66));
  AOI21_X1  g767(.A(new_n345), .B1(new_n563), .B2(G224), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n824), .A2(new_n799), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n954), .B1(new_n955), .B2(new_n345), .ZN(new_n956));
  INV_X1    g770(.A(G898), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n910), .B1(new_n957), .B2(G953), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n956), .B(new_n958), .ZN(G69));
  NAND2_X1  g773(.A1(new_n305), .A2(new_n306), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(new_n521), .Z(new_n961));
  NAND2_X1  g775(.A1(G900), .A2(G953), .ZN(new_n962));
  AND3_X1   g776(.A1(new_n757), .A2(new_n396), .A3(new_n803), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n781), .B1(new_n790), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n802), .A2(new_n715), .ZN(new_n965));
  AOI211_X1 g779(.A(new_n765), .B(new_n965), .C1(new_n768), .C2(new_n848), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n964), .A2(new_n796), .A3(new_n966), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n961), .B(new_n962), .C1(new_n967), .C2(G953), .ZN(new_n968));
  AOI211_X1 g782(.A(new_n759), .B(new_n701), .C1(new_n893), .C2(new_n767), .ZN(new_n969));
  AOI22_X1  g783(.A1(new_n794), .A2(new_n795), .B1(new_n732), .B2(new_n969), .ZN(new_n970));
  OR3_X1    g784(.A1(new_n705), .A2(new_n965), .A3(KEYINPUT62), .ZN(new_n971));
  OAI21_X1  g785(.A(KEYINPUT62), .B1(new_n705), .B2(new_n965), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n970), .A2(new_n791), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n973), .A2(new_n345), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n968), .B1(new_n974), .B2(new_n961), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n345), .B1(G227), .B2(G900), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(G72));
  NAND2_X1  g791(.A1(G472), .A2(G902), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT63), .Z(new_n979));
  OAI21_X1  g793(.A(new_n979), .B1(new_n973), .B2(new_n955), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n980), .A2(new_n282), .A3(new_n308), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n979), .B1(new_n967), .B2(new_n955), .ZN(new_n982));
  INV_X1    g796(.A(new_n308), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n982), .A2(new_n309), .A3(new_n983), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n981), .A2(new_n905), .A3(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n869), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n320), .B(new_n322), .C1(new_n983), .C2(new_n282), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n979), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT127), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n985), .B1(new_n986), .B2(new_n989), .ZN(G57));
endmodule


