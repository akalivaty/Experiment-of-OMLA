//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 1 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 1 1 1 1 1 1 1 0 1 0 1 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:12 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990;
  INV_X1    g000(.A(G116), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT67), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT67), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G116), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n188), .A2(new_n190), .A3(G119), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT66), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT66), .A2(G119), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(G116), .A3(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G113), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT2), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT2), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G113), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  AND3_X1   g015(.A1(new_n191), .A2(new_n196), .A3(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n201), .B1(new_n191), .B2(new_n196), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G143), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(KEYINPUT0), .A2(G128), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT64), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(G143), .B(G146), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n213));
  AND2_X1   g027(.A1(KEYINPUT0), .A2(G128), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(KEYINPUT0), .A2(G128), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g031(.A1(new_n211), .A2(new_n215), .B1(new_n209), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT11), .ZN(new_n219));
  INV_X1    g033(.A(G134), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n219), .B1(new_n220), .B2(G137), .ZN(new_n221));
  INV_X1    g035(.A(G137), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n222), .A2(KEYINPUT11), .A3(G134), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n220), .A2(G137), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n221), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G131), .ZN(new_n226));
  INV_X1    g040(.A(G131), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n221), .A2(new_n223), .A3(new_n227), .A4(new_n224), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(KEYINPUT1), .B1(new_n207), .B2(G146), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n209), .A2(G128), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G128), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n206), .B(new_n208), .C1(KEYINPUT1), .C2(new_n232), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(new_n222), .A3(G134), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT65), .B1(new_n220), .B2(G137), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n222), .A2(G134), .ZN(new_n238));
  OAI211_X1 g052(.A(G131), .B(new_n236), .C1(new_n237), .C2(new_n238), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n239), .A2(new_n228), .ZN(new_n240));
  AOI22_X1  g054(.A1(new_n218), .A2(new_n229), .B1(new_n234), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT30), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n231), .A2(new_n239), .A3(new_n228), .A4(new_n233), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n226), .A2(new_n228), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n209), .A2(new_n217), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n213), .B1(new_n212), .B2(new_n214), .ZN(new_n247));
  AND4_X1   g061(.A1(new_n213), .A2(new_n206), .A3(new_n208), .A4(new_n214), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n244), .B1(new_n245), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT30), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n204), .B1(new_n243), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n211), .A2(new_n215), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n229), .A2(new_n253), .A3(new_n246), .ZN(new_n254));
  AND3_X1   g068(.A1(new_n254), .A2(new_n204), .A3(new_n244), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G237), .ZN(new_n257));
  INV_X1    g071(.A(G953), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(new_n258), .A3(G210), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n259), .B(KEYINPUT27), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT26), .B(G101), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n260), .B(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(KEYINPUT31), .B1(new_n256), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT31), .ZN(new_n264));
  INV_X1    g078(.A(new_n262), .ZN(new_n265));
  NOR4_X1   g079(.A1(new_n252), .A2(new_n264), .A3(new_n255), .A4(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(KEYINPUT28), .B1(new_n241), .B2(new_n204), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n191), .A2(new_n196), .ZN(new_n268));
  INV_X1    g082(.A(new_n201), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n191), .A2(new_n196), .A3(new_n201), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n250), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n254), .A2(new_n204), .A3(new_n244), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n267), .B1(new_n275), .B2(KEYINPUT28), .ZN(new_n276));
  OAI22_X1  g090(.A1(new_n263), .A2(new_n266), .B1(new_n276), .B2(new_n262), .ZN(new_n277));
  NOR2_X1   g091(.A1(G472), .A2(G902), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT32), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT32), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n277), .A2(new_n281), .A3(new_n278), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT69), .B1(new_n241), .B2(new_n204), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n284), .B1(new_n275), .B2(KEYINPUT69), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT28), .ZN(new_n286));
  OAI21_X1  g100(.A(KEYINPUT70), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n267), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT70), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT69), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n290), .B1(new_n273), .B2(new_n274), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n289), .B(KEYINPUT28), .C1(new_n291), .C2(new_n284), .ZN(new_n292));
  AND2_X1   g106(.A1(new_n262), .A2(KEYINPUT29), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n287), .A2(new_n288), .A3(new_n292), .A4(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT71), .ZN(new_n295));
  INV_X1    g109(.A(G902), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n204), .B1(new_n254), .B2(new_n244), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT69), .B1(new_n255), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n274), .A2(new_n290), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n286), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n267), .B1(new_n300), .B2(new_n289), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT71), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n301), .A2(new_n302), .A3(new_n287), .A4(new_n293), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n243), .A2(new_n251), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n272), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n274), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n306), .A2(KEYINPUT68), .A3(new_n265), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT68), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n308), .B1(new_n256), .B2(new_n262), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT29), .B1(new_n276), .B2(new_n262), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n307), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n295), .A2(new_n296), .A3(new_n303), .A4(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G472), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n283), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G217), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n315), .B1(G234), .B2(new_n296), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT22), .B(G137), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n258), .A2(G221), .A3(G234), .ZN(new_n319));
  XOR2_X1   g133(.A(new_n318), .B(new_n319), .Z(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT23), .ZN(new_n322));
  AND2_X1   g136(.A1(KEYINPUT66), .A2(G119), .ZN(new_n323));
  NOR2_X1   g137(.A1(KEYINPUT66), .A2(G119), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n322), .B1(new_n325), .B2(G128), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n194), .A2(G128), .A3(new_n195), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n232), .A2(G119), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n326), .B(new_n327), .C1(new_n322), .C2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G110), .ZN(new_n330));
  INV_X1    g144(.A(G140), .ZN(new_n331));
  INV_X1    g145(.A(G125), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT75), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G125), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n331), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(G125), .A2(G140), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT16), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n333), .A2(new_n335), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT16), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(new_n340), .A3(new_n331), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n338), .A2(G146), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(G146), .B1(new_n338), .B2(new_n341), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n330), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT24), .B(G110), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT72), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n347), .B1(G119), .B2(new_n232), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n327), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT73), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n194), .A2(new_n347), .A3(G128), .A4(new_n195), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n350), .B1(new_n349), .B2(new_n351), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n346), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT74), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n328), .A2(KEYINPUT72), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n356), .B1(new_n325), .B2(G128), .ZN(new_n357));
  INV_X1    g171(.A(new_n351), .ZN(new_n358));
  OAI21_X1  g172(.A(KEYINPUT73), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT74), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n362), .A3(new_n346), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n344), .B1(new_n355), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n327), .B1(new_n322), .B2(new_n328), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n194), .A2(new_n195), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT23), .B1(new_n366), .B2(new_n232), .ZN(new_n367));
  NOR3_X1   g181(.A1(new_n365), .A2(new_n367), .A3(G110), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n352), .A2(new_n353), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n368), .B1(new_n369), .B2(new_n345), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n338), .A2(G146), .A3(new_n341), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT76), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n338), .A2(KEYINPUT76), .A3(G146), .A4(new_n341), .ZN(new_n374));
  XNOR2_X1  g188(.A(G125), .B(G140), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n205), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n373), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n370), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n321), .B1(new_n364), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n343), .ZN(new_n380));
  AOI22_X1  g194(.A1(new_n380), .A2(new_n371), .B1(G110), .B2(new_n329), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n362), .B1(new_n361), .B2(new_n346), .ZN(new_n382));
  AOI211_X1 g196(.A(KEYINPUT74), .B(new_n345), .C1(new_n359), .C2(new_n360), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n368), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n385), .B1(new_n361), .B2(new_n346), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n386), .A2(new_n373), .A3(new_n374), .A4(new_n376), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n384), .A2(new_n387), .A3(new_n320), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n379), .A2(new_n296), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT25), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n379), .A2(new_n388), .A3(KEYINPUT25), .A4(new_n296), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n317), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n316), .A2(G902), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n395), .B(KEYINPUT77), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n379), .A2(new_n396), .A3(new_n388), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n314), .A2(new_n398), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n191), .A2(new_n196), .A3(KEYINPUT5), .ZN(new_n400));
  OAI21_X1  g214(.A(G113), .B1(new_n196), .B2(KEYINPUT5), .ZN(new_n401));
  OAI21_X1  g215(.A(KEYINPUT81), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n191), .A2(new_n196), .A3(KEYINPUT5), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT81), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT5), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n325), .A2(new_n405), .A3(G116), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n403), .A2(new_n404), .A3(G113), .A4(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n402), .A2(new_n271), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(G104), .ZN(new_n409));
  OAI21_X1  g223(.A(KEYINPUT3), .B1(new_n409), .B2(G107), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT3), .ZN(new_n411));
  INV_X1    g225(.A(G107), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(new_n412), .A3(G104), .ZN(new_n413));
  INV_X1    g227(.A(G101), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n409), .A2(G107), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n410), .A2(new_n413), .A3(new_n414), .A4(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n409), .A2(G107), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n412), .A2(G104), .ZN(new_n418));
  OAI21_X1  g232(.A(G101), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n202), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n403), .A2(G113), .A3(new_n406), .ZN(new_n422));
  AOI22_X1  g236(.A1(new_n408), .A2(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(G110), .B(G122), .ZN(new_n424));
  XOR2_X1   g238(.A(new_n424), .B(KEYINPUT8), .Z(new_n425));
  NAND2_X1  g239(.A1(new_n231), .A2(new_n233), .ZN(new_n426));
  XNOR2_X1  g240(.A(KEYINPUT75), .B(G125), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n428), .B1(new_n218), .B2(new_n427), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT7), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n258), .A2(G224), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT90), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n430), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n434), .B1(new_n433), .B2(new_n432), .ZN(new_n435));
  OAI22_X1  g249(.A1(new_n423), .A2(new_n425), .B1(new_n429), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n428), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT88), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n437), .A2(new_n438), .B1(KEYINPUT7), .B2(new_n431), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n439), .B1(new_n438), .B2(new_n429), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT89), .ZN(new_n441));
  OR2_X1    g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(new_n441), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n436), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n402), .A2(new_n421), .A3(new_n407), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n410), .A2(new_n413), .A3(new_n415), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(G101), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(KEYINPUT4), .A3(new_n416), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT4), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n446), .A2(new_n449), .A3(G101), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n272), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n445), .A2(new_n451), .A3(new_n424), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT84), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT84), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n445), .A2(new_n454), .A3(new_n451), .A4(new_n424), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(G902), .B1(new_n444), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(KEYINPUT82), .B1(new_n445), .B2(new_n451), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n445), .A2(KEYINPUT82), .A3(new_n451), .ZN(new_n460));
  XOR2_X1   g274(.A(new_n424), .B(KEYINPUT83), .Z(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n459), .A2(KEYINPUT6), .A3(new_n460), .A4(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT6), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n464), .B1(new_n453), .B2(new_n455), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n445), .A2(KEYINPUT82), .A3(new_n451), .ZN(new_n466));
  NOR3_X1   g280(.A1(new_n466), .A2(new_n458), .A3(new_n461), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n463), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n431), .B(KEYINPUT85), .ZN(new_n469));
  XOR2_X1   g283(.A(new_n469), .B(KEYINPUT86), .Z(new_n470));
  XNOR2_X1  g284(.A(new_n429), .B(new_n470), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n468), .A2(KEYINPUT87), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(KEYINPUT87), .B1(new_n468), .B2(new_n471), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n457), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(G210), .B1(G237), .B2(G902), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n475), .B(KEYINPUT91), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n476), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n478), .B(new_n457), .C1(new_n472), .C2(new_n473), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(G214), .B1(G237), .B2(G902), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(G221), .ZN(new_n485));
  XNOR2_X1  g299(.A(KEYINPUT9), .B(G234), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n485), .B1(new_n487), .B2(new_n296), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n258), .A2(G227), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(KEYINPUT78), .ZN(new_n491));
  XNOR2_X1  g305(.A(G110), .B(G140), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n491), .B(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT12), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n426), .A2(new_n420), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n231), .A2(new_n233), .A3(new_n416), .A4(new_n419), .ZN(new_n497));
  AOI221_X4 g311(.A(new_n495), .B1(new_n228), .B2(new_n226), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n497), .ZN(new_n499));
  AOI21_X1  g313(.A(KEYINPUT12), .B1(new_n499), .B2(new_n229), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n218), .A2(new_n448), .A3(new_n450), .ZN(new_n502));
  INV_X1    g316(.A(new_n420), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n234), .A2(new_n503), .A3(KEYINPUT10), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT10), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n497), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n502), .A2(new_n504), .A3(new_n245), .A4(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n494), .B1(new_n501), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT79), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n502), .A2(new_n506), .A3(new_n504), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n229), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n512), .A2(new_n507), .A3(new_n493), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n509), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n510), .B1(new_n509), .B2(new_n513), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n296), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n516), .A2(G469), .ZN(new_n517));
  INV_X1    g331(.A(G469), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n507), .A2(new_n493), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n501), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n493), .B1(new_n512), .B2(new_n507), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n518), .B(new_n296), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT80), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n497), .B(KEYINPUT10), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n245), .B1(new_n525), .B2(new_n502), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n494), .B1(new_n526), .B2(new_n508), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n507), .B(new_n493), .C1(new_n498), .C2(new_n500), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n529), .A2(KEYINPUT80), .A3(new_n518), .A4(new_n296), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n524), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n489), .B1(new_n517), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n342), .A2(new_n343), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n257), .A2(new_n258), .A3(G214), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n535), .B(new_n207), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n536), .A2(KEYINPUT17), .A3(G131), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(G131), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n535), .B(G143), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n227), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n534), .B(new_n537), .C1(KEYINPUT17), .C2(new_n541), .ZN(new_n542));
  XNOR2_X1  g356(.A(G113), .B(G122), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(new_n409), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT18), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n539), .B1(new_n545), .B2(new_n227), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n536), .A2(KEYINPUT18), .A3(G131), .ZN(new_n547));
  INV_X1    g361(.A(new_n337), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n548), .B1(new_n427), .B2(new_n331), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n376), .B1(new_n549), .B2(new_n205), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n546), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n542), .A2(new_n544), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n544), .B1(new_n542), .B2(new_n551), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n296), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(G475), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n373), .A2(new_n374), .A3(new_n541), .ZN(new_n557));
  OAI211_X1 g371(.A(KEYINPUT19), .B(new_n548), .C1(new_n427), .C2(new_n331), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT19), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n375), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n558), .A2(new_n205), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT92), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n558), .A2(KEYINPUT92), .A3(new_n205), .A4(new_n560), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI211_X1 g379(.A(KEYINPUT93), .B(new_n551), .C1(new_n557), .C2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n544), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n563), .A2(new_n564), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n569), .A2(new_n373), .A3(new_n374), .A4(new_n541), .ZN(new_n570));
  AOI21_X1  g384(.A(KEYINPUT93), .B1(new_n570), .B2(new_n551), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n552), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT20), .ZN(new_n573));
  NOR2_X1   g387(.A1(G475), .A2(G902), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n573), .B1(new_n572), .B2(new_n574), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n556), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(G128), .B(G143), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(new_n220), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n188), .A2(new_n190), .A3(G122), .ZN(new_n580));
  INV_X1    g394(.A(G122), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(G116), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n579), .B1(G107), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n580), .A2(KEYINPUT14), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT14), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n580), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n585), .B1(KEYINPUT94), .B2(new_n588), .ZN(new_n589));
  OR2_X1    g403(.A1(new_n588), .A2(KEYINPUT94), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n584), .B1(new_n591), .B2(G107), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n583), .B(new_n412), .ZN(new_n593));
  AOI21_X1  g407(.A(KEYINPUT13), .B1(new_n232), .B2(G143), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n594), .A2(new_n220), .ZN(new_n595));
  XOR2_X1   g409(.A(new_n595), .B(new_n578), .Z(new_n596));
  NOR2_X1   g410(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  NOR3_X1   g411(.A1(new_n486), .A2(new_n315), .A3(G953), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  OR3_X1    g413(.A1(new_n592), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n599), .B1(new_n592), .B2(new_n597), .ZN(new_n601));
  AOI21_X1  g415(.A(G902), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(G478), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(KEYINPUT15), .ZN(new_n604));
  XOR2_X1   g418(.A(new_n602), .B(new_n604), .Z(new_n605));
  OR2_X1    g419(.A1(new_n577), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(G952), .ZN(new_n607));
  AOI211_X1 g421(.A(G953), .B(new_n607), .C1(G234), .C2(G237), .ZN(new_n608));
  AOI211_X1 g422(.A(new_n296), .B(new_n258), .C1(G234), .C2(G237), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT21), .B(G898), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n533), .A2(new_n606), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n399), .A2(new_n484), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(G101), .ZN(G3));
  INV_X1    g428(.A(KEYINPUT95), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n477), .A2(new_n615), .A3(new_n479), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n600), .A2(new_n601), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(KEYINPUT33), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n600), .A2(new_n619), .A3(new_n601), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n618), .A2(G478), .A3(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n603), .A2(new_n296), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n602), .B2(new_n603), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n577), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n474), .A2(KEYINPUT95), .A3(new_n476), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n616), .A2(new_n482), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n611), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n276), .A2(new_n262), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n305), .A2(new_n274), .A3(new_n262), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n264), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n256), .A2(KEYINPUT31), .A3(new_n262), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n631), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g449(.A(G472), .B1(new_n635), .B2(G902), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n279), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n533), .A2(new_n398), .A3(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n630), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT34), .B(G104), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G6));
  OAI211_X1 g456(.A(new_n605), .B(new_n556), .C1(new_n576), .C2(new_n575), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n616), .A2(new_n482), .A3(new_n626), .A4(new_n644), .ZN(new_n645));
  OR2_X1    g459(.A1(new_n645), .A2(new_n611), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n646), .A2(new_n639), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT96), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT35), .B(G107), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  OAI22_X1  g464(.A1(new_n364), .A2(new_n378), .B1(KEYINPUT36), .B2(new_n321), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n321), .A2(KEYINPUT36), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n384), .A2(new_n387), .A3(new_n652), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n651), .A2(new_n396), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n391), .A2(new_n392), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n654), .B1(new_n655), .B2(new_n316), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n637), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n484), .A2(new_n612), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT37), .B(G110), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G12));
  NAND2_X1  g474(.A1(new_n283), .A2(new_n313), .ZN(new_n661));
  INV_X1    g475(.A(new_n656), .ZN(new_n662));
  INV_X1    g476(.A(G900), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n609), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n608), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n516), .A2(G469), .ZN(new_n668));
  AOI211_X1 g482(.A(new_n488), .B(new_n667), .C1(new_n668), .C2(new_n531), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n661), .A2(new_n662), .A3(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n645), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(new_n232), .ZN(G30));
  XNOR2_X1  g486(.A(new_n666), .B(KEYINPUT39), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  OR2_X1    g488(.A1(new_n533), .A2(new_n674), .ZN(new_n675));
  OR2_X1    g489(.A1(new_n675), .A2(KEYINPUT40), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(KEYINPUT40), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n577), .A2(new_n605), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n306), .A2(new_n262), .ZN(new_n679));
  AOI21_X1  g493(.A(G902), .B1(new_n285), .B2(new_n265), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(G472), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n283), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n684), .A2(new_n483), .A3(new_n662), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n676), .A2(new_n677), .A3(new_n678), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n480), .B(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT98), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G143), .ZN(G45));
  INV_X1    g507(.A(new_n670), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n628), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G146), .ZN(G48));
  AOI21_X1  g510(.A(new_n518), .B1(new_n529), .B2(new_n296), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT99), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n531), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n488), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n399), .A2(new_n700), .ZN(new_n701));
  OR2_X1    g515(.A1(new_n630), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT41), .B(G113), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G15));
  OR2_X1    g518(.A1(new_n646), .A2(new_n701), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G116), .ZN(G18));
  NAND2_X1  g520(.A1(new_n468), .A2(new_n471), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT87), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n468), .A2(KEYINPUT87), .A3(new_n471), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n478), .B1(new_n711), .B2(new_n457), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n483), .B1(new_n712), .B2(KEYINPUT95), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n713), .A2(new_n616), .A3(new_n700), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n606), .A2(new_n611), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n314), .A2(new_n656), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT100), .ZN(new_n718));
  OR2_X1    g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n717), .A2(new_n718), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G119), .ZN(G21));
  INV_X1    g536(.A(KEYINPUT101), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n577), .A2(new_n723), .A3(new_n605), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n723), .B1(new_n577), .B2(new_n605), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n398), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n262), .B1(new_n301), .B2(new_n287), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n263), .A2(new_n266), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n278), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n727), .A2(new_n636), .A3(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n714), .A2(new_n629), .A3(new_n726), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G122), .ZN(G24));
  OAI211_X1 g547(.A(new_n730), .B(new_n636), .C1(new_n393), .C2(new_n654), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n577), .A2(new_n624), .A3(new_n666), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n713), .A2(new_n736), .A3(new_n616), .A4(new_n700), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G125), .ZN(G27));
  XNOR2_X1  g552(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n739));
  NAND2_X1  g553(.A1(KEYINPUT102), .A2(KEYINPUT42), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n480), .A2(new_n483), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n509), .A2(new_n513), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n296), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(G469), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n488), .B1(new_n531), .B2(new_n744), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n735), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(new_n399), .A3(new_n747), .ZN(new_n748));
  MUX2_X1   g562(.A(new_n739), .B(new_n740), .S(new_n748), .Z(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G131), .ZN(G33));
  NAND4_X1  g564(.A1(new_n746), .A2(new_n399), .A3(new_n644), .A4(new_n666), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G134), .ZN(G36));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n753));
  OAI21_X1  g567(.A(G469), .B1(new_n742), .B2(new_n753), .ZN(new_n754));
  OR2_X1    g568(.A1(new_n514), .A2(new_n515), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n754), .B1(new_n755), .B2(new_n753), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n518), .A2(new_n296), .ZN(new_n757));
  OR2_X1    g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT46), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n532), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n760), .B1(new_n759), .B2(new_n758), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n489), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n673), .A3(new_n741), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT44), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n624), .B(new_n556), .C1(new_n576), .C2(new_n575), .ZN(new_n766));
  XOR2_X1   g580(.A(new_n766), .B(KEYINPUT43), .Z(new_n767));
  OR2_X1    g581(.A1(new_n767), .A2(KEYINPUT103), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(KEYINPUT103), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n768), .A2(new_n637), .A3(new_n662), .A4(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n764), .B1(new_n765), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n771), .B1(new_n765), .B2(new_n770), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G137), .ZN(G39));
  OR2_X1    g587(.A1(KEYINPUT104), .A2(KEYINPUT47), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n762), .A2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n741), .ZN(new_n776));
  NOR4_X1   g590(.A1(new_n776), .A2(new_n661), .A3(new_n727), .A4(new_n735), .ZN(new_n777));
  XOR2_X1   g591(.A(KEYINPUT104), .B(KEYINPUT47), .Z(new_n778));
  OAI211_X1 g592(.A(new_n775), .B(new_n777), .C1(new_n762), .C2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G140), .ZN(G42));
  XOR2_X1   g594(.A(new_n699), .B(KEYINPUT49), .Z(new_n781));
  NOR3_X1   g595(.A1(new_n398), .A2(new_n483), .A3(new_n488), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n781), .A2(new_n684), .A3(new_n782), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n783), .A2(new_n688), .A3(new_n766), .ZN(new_n784));
  XOR2_X1   g598(.A(new_n784), .B(KEYINPUT105), .Z(new_n785));
  AND2_X1   g599(.A1(new_n767), .A2(new_n608), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n731), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  AOI211_X1 g602(.A(new_n607), .B(G953), .C1(new_n788), .C2(new_n714), .ZN(new_n789));
  INV_X1    g603(.A(new_n700), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n776), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n786), .A2(new_n399), .A3(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(KEYINPUT48), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n789), .A2(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n791), .A2(new_n684), .A3(new_n727), .A4(new_n608), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT114), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n794), .B1(new_n625), .B2(new_n797), .ZN(new_n798));
  OR3_X1    g612(.A1(new_n796), .A2(new_n577), .A3(new_n624), .ZN(new_n799));
  NOR4_X1   g613(.A1(new_n787), .A2(new_n482), .A3(new_n688), .A4(new_n790), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT50), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n786), .A2(new_n791), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n799), .B(new_n801), .C1(new_n734), .C2(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n775), .B1(new_n762), .B2(new_n778), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n804), .B1(new_n489), .B2(new_n699), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n741), .A3(new_n788), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(KEYINPUT51), .ZN(new_n807));
  XOR2_X1   g621(.A(new_n806), .B(KEYINPUT113), .Z(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(new_n803), .ZN(new_n809));
  OAI221_X1 g623(.A(new_n798), .B1(new_n803), .B2(new_n807), .C1(new_n809), .C2(KEYINPUT51), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n719), .A2(new_n720), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n702), .A2(new_n705), .A3(new_n732), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OR2_X1    g627(.A1(new_n644), .A2(new_n625), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n484), .A2(new_n629), .A3(new_n638), .A4(new_n814), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n815), .A2(new_n613), .A3(new_n658), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n776), .A2(new_n606), .ZN(new_n817));
  AOI22_X1  g631(.A1(new_n817), .A2(new_n694), .B1(new_n746), .B2(new_n736), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n816), .A2(new_n751), .A3(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n813), .A2(new_n749), .A3(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n726), .A2(new_n713), .A3(new_n616), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT106), .ZN(new_n823));
  AND4_X1   g637(.A1(new_n823), .A2(new_n745), .A3(new_n656), .A4(new_n666), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n393), .A2(new_n654), .A3(new_n667), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n823), .B1(new_n825), .B2(new_n745), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n683), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  OAI22_X1  g641(.A1(new_n822), .A2(new_n827), .B1(new_n627), .B2(new_n670), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  AND4_X1   g643(.A1(new_n616), .A2(new_n713), .A3(new_n736), .A4(new_n700), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n671), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT107), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n829), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT52), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n737), .B1(new_n645), .B2(new_n670), .ZN(new_n835));
  OAI21_X1  g649(.A(KEYINPUT107), .B1(new_n828), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n833), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n837), .A2(KEYINPUT108), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT108), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n833), .A2(new_n839), .A3(new_n834), .A4(new_n836), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n829), .A2(new_n831), .A3(KEYINPUT52), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT109), .B1(new_n838), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n837), .A2(KEYINPUT108), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT109), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n844), .A2(new_n845), .A3(new_n841), .A4(new_n840), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n821), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n812), .ZN(new_n848));
  AND4_X1   g662(.A1(new_n721), .A2(new_n848), .A3(new_n820), .A4(new_n749), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n833), .A2(new_n836), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT52), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(new_n837), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  XOR2_X1   g667(.A(KEYINPUT110), .B(KEYINPUT53), .Z(new_n854));
  OAI22_X1  g668(.A1(new_n847), .A2(KEYINPUT53), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT54), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n857), .B1(new_n819), .B2(KEYINPUT112), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT112), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n816), .A2(new_n859), .A3(new_n751), .A4(new_n818), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n813), .A2(new_n858), .A3(new_n749), .A4(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n840), .A2(new_n841), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n845), .B1(new_n863), .B2(new_n844), .ZN(new_n864));
  AND4_X1   g678(.A1(new_n845), .A2(new_n844), .A3(new_n841), .A4(new_n840), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n862), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n853), .A2(new_n854), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n856), .B(KEYINPUT111), .C1(KEYINPUT54), .C2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT111), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n855), .A2(new_n870), .A3(KEYINPUT54), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n810), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(G952), .A2(G953), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(KEYINPUT115), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n785), .B1(new_n872), .B2(new_n874), .ZN(G75));
  NOR2_X1   g689(.A1(new_n258), .A2(G952), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n868), .A2(G902), .A3(new_n476), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT117), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n468), .B(new_n471), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n880), .B(KEYINPUT55), .Z(new_n881));
  INV_X1    g695(.A(KEYINPUT56), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n878), .A2(new_n879), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n879), .B1(new_n878), .B2(new_n883), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n877), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n878), .A2(KEYINPUT116), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT56), .B1(new_n878), .B2(KEYINPUT116), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n881), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n886), .A2(new_n889), .ZN(G51));
  AOI21_X1  g704(.A(new_n861), .B1(new_n843), .B2(new_n846), .ZN(new_n891));
  INV_X1    g705(.A(new_n854), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n892), .B1(new_n849), .B2(new_n852), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT54), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n894), .B(new_n895), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n757), .B(KEYINPUT57), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n529), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n894), .A2(new_n296), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(new_n756), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n876), .B1(new_n899), .B2(new_n901), .ZN(G54));
  NAND3_X1  g716(.A1(new_n900), .A2(KEYINPUT58), .A3(G475), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT118), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n904), .A2(new_n905), .A3(new_n572), .ZN(new_n906));
  INV_X1    g720(.A(new_n572), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT118), .B1(new_n903), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n876), .B1(new_n903), .B2(new_n907), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n906), .A2(new_n908), .A3(new_n909), .ZN(G60));
  AND2_X1   g724(.A1(new_n618), .A2(new_n620), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n622), .B(KEYINPUT59), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n896), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n877), .ZN(new_n915));
  INV_X1    g729(.A(new_n912), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n869), .A2(new_n871), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n915), .B1(new_n911), .B2(new_n917), .ZN(G63));
  XNOR2_X1  g732(.A(KEYINPUT119), .B(KEYINPUT60), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n315), .A2(new_n296), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n919), .B(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n921), .B1(new_n891), .B2(new_n893), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n379), .A2(new_n388), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n876), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n651), .A2(new_n653), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n925), .B(new_n921), .C1(new_n891), .C2(new_n893), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n924), .A2(KEYINPUT61), .A3(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT120), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n868), .A2(new_n928), .A3(new_n925), .A4(new_n921), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n926), .A2(KEYINPUT120), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n924), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT121), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT61), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n932), .B1(new_n931), .B2(new_n933), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n927), .B1(new_n934), .B2(new_n935), .ZN(G66));
  INV_X1    g750(.A(new_n610), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n258), .B1(new_n937), .B2(G224), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n813), .A2(new_n816), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT122), .Z(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n938), .B1(new_n941), .B2(new_n258), .ZN(new_n942));
  INV_X1    g756(.A(new_n468), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n943), .B1(G898), .B2(new_n258), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n942), .B(new_n944), .Z(G69));
  NAND2_X1  g759(.A1(new_n558), .A2(new_n560), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT123), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n304), .B(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n831), .A2(new_n695), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n692), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(KEYINPUT62), .ZN(new_n952));
  INV_X1    g766(.A(new_n675), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n953), .A2(new_n399), .A3(new_n741), .A4(new_n814), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n779), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n952), .A2(new_n772), .A3(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT62), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n692), .A2(new_n957), .A3(new_n950), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(KEYINPUT124), .ZN(new_n959));
  OR2_X1    g773(.A1(new_n958), .A2(KEYINPUT124), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n956), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n948), .B1(new_n961), .B2(G953), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n258), .B1(G227), .B2(G900), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n822), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n763), .A2(new_n399), .A3(new_n673), .A4(new_n965), .ZN(new_n966));
  AND4_X1   g780(.A1(new_n749), .A2(new_n779), .A3(new_n751), .A4(new_n966), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n967), .A2(new_n258), .A3(new_n772), .A4(new_n950), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n948), .B1(G900), .B2(G953), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n962), .A2(new_n964), .A3(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT126), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT125), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n970), .B(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n962), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n972), .B1(new_n975), .B2(new_n963), .ZN(new_n976));
  AOI211_X1 g790(.A(KEYINPUT126), .B(new_n964), .C1(new_n962), .C2(new_n974), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n971), .B1(new_n976), .B2(new_n977), .ZN(G72));
  NAND2_X1  g792(.A1(G472), .A2(G902), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT63), .Z(new_n980));
  NAND3_X1  g794(.A1(new_n967), .A2(new_n772), .A3(new_n950), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n980), .B1(new_n941), .B2(new_n981), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n306), .A2(new_n262), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT127), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n980), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n986), .B1(new_n961), .B2(new_n940), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n985), .B(new_n877), .C1(new_n987), .C2(new_n679), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n307), .A2(new_n309), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n986), .B1(new_n989), .B2(new_n632), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n988), .B1(new_n855), .B2(new_n990), .ZN(G57));
endmodule


