//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 0 0 1 1 1 1 1 1 0 1 1 0 1 0 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n809, new_n811, new_n813, new_n814, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n864, new_n865, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918;
  XNOR2_X1  g000(.A(G127gat), .B(G155gat), .ZN(new_n202));
  INV_X1    g001(.A(G211gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G15gat), .B(G22gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT93), .ZN(new_n206));
  INV_X1    g005(.A(G1gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT16), .ZN(new_n208));
  AOI22_X1  g007(.A1(new_n206), .A2(new_n207), .B1(new_n208), .B2(new_n205), .ZN(new_n209));
  NAND2_X1  g008(.A1(KEYINPUT94), .A2(G8gat), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n209), .B(new_n210), .C1(new_n207), .C2(new_n206), .ZN(new_n211));
  NOR2_X1   g010(.A1(KEYINPUT94), .A2(G8gat), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  OR2_X1    g012(.A1(KEYINPUT96), .A2(G57gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(KEYINPUT96), .A2(G57gat), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n214), .B(G64gat), .C1(KEYINPUT97), .C2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G57gat), .ZN(new_n217));
  OR3_X1    g016(.A1(new_n217), .A2(KEYINPUT97), .A3(G64gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n219), .B(KEYINPUT98), .ZN(new_n220));
  AND2_X1   g019(.A1(G71gat), .A2(G78gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(G71gat), .A2(G78gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n220), .B(new_n224), .C1(KEYINPUT9), .C2(new_n221), .ZN(new_n225));
  XNOR2_X1  g024(.A(G57gat), .B(G64gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT9), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n223), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT21), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n213), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G183gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n231), .B(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT99), .ZN(new_n234));
  OR2_X1    g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n234), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n235), .A2(new_n236), .A3(G231gat), .A4(G233gat), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  AOI22_X1  g037(.A1(new_n235), .A2(new_n236), .B1(G231gat), .B2(G233gat), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n204), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n239), .ZN(new_n241));
  INV_X1    g040(.A(new_n204), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n241), .A2(new_n237), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n229), .A2(new_n230), .ZN(new_n244));
  XOR2_X1   g043(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  AND3_X1   g045(.A1(new_n240), .A2(new_n243), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n246), .B1(new_n240), .B2(new_n243), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(G29gat), .ZN(new_n251));
  INV_X1    g050(.A(G36gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n251), .A2(new_n252), .A3(KEYINPUT14), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT14), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n254), .B1(G29gat), .B2(G36gat), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n253), .B(new_n255), .C1(new_n251), .C2(new_n252), .ZN(new_n256));
  XOR2_X1   g055(.A(KEYINPUT91), .B(G43gat), .Z(new_n257));
  INV_X1    g056(.A(G50gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n257), .A2(KEYINPUT92), .A3(new_n258), .ZN(new_n259));
  OR2_X1    g058(.A1(new_n258), .A2(G43gat), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT92), .ZN(new_n261));
  XNOR2_X1  g060(.A(KEYINPUT91), .B(G43gat), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n261), .B1(new_n262), .B2(G50gat), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n259), .A2(new_n260), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT15), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n256), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n258), .A2(G43gat), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n260), .A2(KEYINPUT15), .A3(new_n267), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n268), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n270), .A2(new_n256), .ZN(new_n271));
  OR2_X1    g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT17), .ZN(new_n273));
  NAND2_X1  g072(.A1(G99gat), .A2(G106gat), .ZN(new_n274));
  INV_X1    g073(.A(G85gat), .ZN(new_n275));
  INV_X1    g074(.A(G92gat), .ZN(new_n276));
  AOI22_X1  g075(.A1(KEYINPUT8), .A2(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(KEYINPUT101), .A2(KEYINPUT7), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n278), .B1(new_n275), .B2(new_n276), .ZN(new_n279));
  NAND4_X1  g078(.A1(KEYINPUT101), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n277), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  XOR2_X1   g080(.A(G99gat), .B(G106gat), .Z(new_n282));
  XOR2_X1   g081(.A(new_n281), .B(new_n282), .Z(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  OR3_X1    g083(.A1(new_n269), .A2(KEYINPUT17), .A3(new_n271), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n273), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  AND2_X1   g085(.A1(G232gat), .A2(G233gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT41), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n286), .B(new_n288), .C1(new_n284), .C2(new_n272), .ZN(new_n289));
  XNOR2_X1  g088(.A(G134gat), .B(G162gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n290), .B(KEYINPUT100), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n289), .B(new_n291), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n287), .A2(KEYINPUT41), .ZN(new_n293));
  XNOR2_X1  g092(.A(G190gat), .B(G218gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n292), .B(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n250), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT79), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT2), .ZN(new_n299));
  INV_X1    g098(.A(G155gat), .ZN(new_n300));
  INV_X1    g099(.A(G162gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G155gat), .A2(G162gat), .ZN(new_n303));
  INV_X1    g102(.A(G148gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G141gat), .ZN(new_n305));
  INV_X1    g104(.A(G141gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G148gat), .ZN(new_n307));
  AOI22_X1  g106(.A1(new_n302), .A2(new_n303), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n303), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n305), .A2(new_n307), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT78), .B(KEYINPUT2), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n300), .A2(new_n301), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n308), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT3), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n298), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT1), .ZN(new_n317));
  INV_X1    g116(.A(G113gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n318), .A2(G120gat), .ZN(new_n319));
  INV_X1    g118(.A(G120gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n320), .A2(G113gat), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n317), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(G127gat), .A2(G134gat), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  NOR2_X1   g123(.A1(KEYINPUT70), .A2(G127gat), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(KEYINPUT70), .A2(G127gat), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n326), .A2(G134gat), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n322), .A2(new_n324), .A3(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT71), .B1(new_n320), .B2(G113gat), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT71), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n331), .A2(new_n318), .A3(G120gat), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n330), .B(new_n332), .C1(new_n318), .C2(G120gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(G127gat), .A2(G134gat), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT1), .B1(new_n324), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n329), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n299), .A2(KEYINPUT78), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT78), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT2), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G141gat), .B(G148gat), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n303), .B(new_n313), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n302), .A2(new_n303), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n310), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n346), .A2(KEYINPUT79), .A3(KEYINPUT3), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n314), .A2(new_n315), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n316), .A2(new_n337), .A3(new_n347), .A4(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT4), .B1(new_n337), .B2(new_n346), .ZN(new_n350));
  AND2_X1   g149(.A1(KEYINPUT70), .A2(G127gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n351), .A2(new_n325), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n323), .B1(new_n352), .B2(G134gat), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n353), .A2(new_n322), .B1(new_n333), .B2(new_n335), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT4), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n354), .A2(new_n314), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n350), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n349), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(G225gat), .A2(G233gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n361), .A2(KEYINPUT5), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n350), .A2(new_n356), .A3(KEYINPUT80), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT80), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n364), .B(KEYINPUT4), .C1(new_n337), .C2(new_n346), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n349), .A2(new_n363), .A3(new_n360), .A4(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT5), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n337), .B(new_n346), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n367), .B1(new_n368), .B2(new_n361), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n359), .A2(new_n362), .B1(new_n366), .B2(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT0), .B(G57gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n371), .B(G85gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(G1gat), .B(G29gat), .ZN(new_n373));
  XOR2_X1   g172(.A(new_n372), .B(new_n373), .Z(new_n374));
  AOI21_X1  g173(.A(KEYINPUT6), .B1(new_n370), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT81), .B1(new_n370), .B2(new_n374), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n366), .A2(new_n369), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n349), .A2(new_n357), .A3(new_n362), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n374), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT81), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n375), .A2(new_n376), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT82), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT83), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n379), .A2(new_n385), .A3(KEYINPUT6), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n385), .B1(new_n379), .B2(KEYINPUT6), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n375), .A2(new_n376), .A3(new_n381), .A4(KEYINPUT82), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n384), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(G64gat), .B(G92gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n392), .B(G36gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n393), .B(KEYINPUT77), .ZN(new_n394));
  XOR2_X1   g193(.A(new_n394), .B(G8gat), .Z(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT29), .ZN(new_n397));
  NAND2_X1  g196(.A1(G226gat), .A2(G233gat), .ZN(new_n398));
  INV_X1    g197(.A(G169gat), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT65), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n400), .A2(G176gat), .ZN(new_n401));
  INV_X1    g200(.A(G176gat), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n402), .A2(KEYINPUT65), .ZN(new_n403));
  OAI211_X1 g202(.A(KEYINPUT23), .B(new_n399), .C1(new_n401), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n399), .A2(new_n402), .ZN(new_n405));
  NAND2_X1  g204(.A1(G169gat), .A2(G176gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g207(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n405), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(G190gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n232), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(G183gat), .A2(G190gat), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n412), .A2(KEYINPUT24), .A3(new_n413), .ZN(new_n414));
  OR2_X1    g213(.A1(new_n413), .A2(KEYINPUT24), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n404), .A2(new_n410), .A3(new_n414), .A4(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n417));
  AND3_X1   g216(.A1(new_n416), .A2(KEYINPUT67), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT67), .B1(new_n416), .B2(new_n417), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n414), .A2(new_n415), .ZN(new_n420));
  NOR2_X1   g219(.A1(G169gat), .A2(G176gat), .ZN(new_n421));
  AOI22_X1  g220(.A1(KEYINPUT66), .A2(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n422));
  INV_X1    g221(.A(new_n409), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n421), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT25), .ZN(new_n425));
  AND2_X1   g224(.A1(new_n421), .A2(KEYINPUT23), .ZN(new_n426));
  NOR4_X1   g225(.A1(new_n420), .A2(new_n424), .A3(new_n425), .A4(new_n426), .ZN(new_n427));
  NOR3_X1   g226(.A1(new_n418), .A2(new_n419), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT26), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n405), .A2(new_n429), .A3(new_n406), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n421), .A2(KEYINPUT26), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n430), .A2(new_n413), .A3(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(KEYINPUT69), .ZN(new_n433));
  XNOR2_X1  g232(.A(KEYINPUT27), .B(G183gat), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n434), .A2(new_n411), .ZN(new_n435));
  OR2_X1    g234(.A1(new_n435), .A2(KEYINPUT28), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT68), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n434), .B(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n438), .A2(KEYINPUT28), .A3(new_n411), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n433), .B1(new_n436), .B2(new_n439), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n397), .B(new_n398), .C1(new_n428), .C2(new_n440), .ZN(new_n441));
  XOR2_X1   g240(.A(KEYINPUT76), .B(KEYINPUT22), .Z(new_n442));
  NAND2_X1  g241(.A1(G211gat), .A2(G218gat), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OR2_X1    g243(.A1(G211gat), .A2(G218gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n443), .ZN(new_n446));
  XNOR2_X1  g245(.A(G197gat), .B(G204gat), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n444), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n447), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n443), .B(new_n445), .C1(new_n449), .C2(new_n442), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n416), .A2(new_n417), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT67), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n427), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n416), .A2(KEYINPUT67), .A3(new_n417), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n439), .A2(new_n436), .ZN(new_n459));
  XOR2_X1   g258(.A(new_n432), .B(KEYINPUT69), .Z(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n398), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n458), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  AND3_X1   g262(.A1(new_n441), .A2(new_n452), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n452), .B1(new_n441), .B2(new_n463), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n396), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n441), .A2(new_n463), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n451), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n441), .A2(new_n452), .A3(new_n463), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n468), .A2(new_n469), .A3(new_n395), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n466), .A2(new_n470), .A3(KEYINPUT30), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n464), .A2(new_n465), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT30), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(new_n473), .A3(new_n395), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n391), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n451), .B1(new_n348), .B2(new_n397), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(G228gat), .ZN(new_n479));
  INV_X1    g278(.A(G233gat), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT3), .B1(new_n451), .B2(new_n397), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n478), .B(new_n481), .C1(new_n314), .C2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n481), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n451), .A2(new_n397), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n314), .B1(new_n485), .B2(new_n315), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n484), .B1(new_n486), .B2(new_n477), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(G22gat), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n488), .A2(KEYINPUT84), .A3(new_n489), .ZN(new_n490));
  XOR2_X1   g289(.A(G78gat), .B(G106gat), .Z(new_n491));
  XNOR2_X1  g290(.A(new_n491), .B(KEYINPUT31), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n492), .B(new_n258), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n489), .A2(KEYINPUT84), .ZN(new_n495));
  OR2_X1    g294(.A1(new_n489), .A2(KEYINPUT84), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n483), .A2(new_n487), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n490), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  AND2_X1   g298(.A1(KEYINPUT85), .A2(G22gat), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n483), .A2(new_n487), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n501), .B1(new_n483), .B2(new_n487), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n493), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT86), .ZN(new_n506));
  NOR4_X1   g305(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT86), .A4(new_n494), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n499), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n476), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n337), .B1(new_n428), .B2(new_n440), .ZN(new_n511));
  NAND2_X1  g310(.A1(G227gat), .A2(G233gat), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n458), .A2(new_n461), .A3(new_n354), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n515), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n511), .A2(new_n512), .A3(new_n513), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G15gat), .B(G43gat), .ZN(new_n521));
  INV_X1    g320(.A(G71gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n521), .B(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(G99gat), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n512), .B1(new_n511), .B2(new_n513), .ZN(new_n525));
  XNOR2_X1  g324(.A(KEYINPUT72), .B(KEYINPUT33), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT32), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n524), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT73), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT73), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n532), .B(new_n524), .C1(new_n525), .C2(new_n529), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n524), .A2(new_n526), .ZN(new_n535));
  NOR3_X1   g334(.A1(new_n525), .A2(new_n527), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n520), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  AOI211_X1 g337(.A(new_n536), .B(new_n519), .C1(new_n531), .C2(new_n533), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT75), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT36), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g341(.A(KEYINPUT75), .B(KEYINPUT36), .C1(new_n538), .C2(new_n539), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n510), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT87), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n375), .B1(new_n374), .B2(new_n370), .ZN(new_n547));
  INV_X1    g346(.A(new_n388), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n547), .A2(new_n548), .A3(new_n386), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT89), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n468), .A2(new_n550), .A3(new_n469), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n551), .B(KEYINPUT37), .C1(new_n550), .C2(new_n469), .ZN(new_n552));
  XNOR2_X1  g351(.A(KEYINPUT90), .B(KEYINPUT37), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n395), .B1(new_n472), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(KEYINPUT38), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(KEYINPUT37), .B1(new_n464), .B2(new_n465), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n468), .A2(new_n469), .A3(new_n553), .ZN(new_n557));
  AND4_X1   g356(.A1(KEYINPUT38), .A2(new_n556), .A3(new_n557), .A4(new_n396), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n549), .B(new_n470), .C1(new_n555), .C2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT88), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n475), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n471), .A2(KEYINPUT88), .A3(new_n474), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n358), .A2(new_n361), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n563), .B(KEYINPUT39), .C1(new_n361), .C2(new_n368), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n564), .B(new_n374), .C1(KEYINPUT39), .C2(new_n563), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT40), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n379), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n565), .A2(new_n566), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n561), .A2(new_n562), .A3(new_n567), .A4(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT86), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n570), .B1(new_n504), .B2(new_n493), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n498), .B1(new_n571), .B2(new_n507), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n559), .A2(new_n569), .A3(new_n572), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n510), .A2(new_n542), .A3(KEYINPUT87), .A4(new_n543), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n546), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NOR3_X1   g374(.A1(new_n509), .A2(new_n538), .A3(new_n539), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n549), .B1(new_n561), .B2(new_n562), .ZN(new_n577));
  AOI21_X1  g376(.A(KEYINPUT35), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n534), .A2(new_n537), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(new_n519), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n534), .A2(new_n537), .A3(new_n520), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n580), .A2(KEYINPUT35), .A3(new_n572), .A4(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n582), .A2(new_n476), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n575), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n272), .A2(new_n213), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT95), .ZN(new_n587));
  NAND2_X1  g386(.A1(G229gat), .A2(G233gat), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n273), .A2(new_n213), .A3(new_n285), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT18), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n272), .A2(new_n213), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n587), .A2(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n588), .B(KEYINPUT13), .Z(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n587), .A2(KEYINPUT18), .A3(new_n588), .A4(new_n589), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n592), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(KEYINPUT11), .B(G169gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(G197gat), .ZN(new_n600));
  XOR2_X1   g399(.A(G113gat), .B(G141gat), .Z(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT12), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n598), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n592), .A2(new_n596), .A3(new_n603), .A4(new_n597), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n229), .A2(new_n284), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT10), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n225), .A2(new_n228), .A3(new_n283), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n611), .A2(new_n610), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(G230gat), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n615), .A2(new_n480), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n609), .A2(new_n611), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(new_n616), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G176gat), .B(G204gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT102), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(G120gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(new_n304), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n618), .A2(new_n620), .A3(new_n625), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n608), .A2(new_n629), .ZN(new_n630));
  AND3_X1   g429(.A1(new_n297), .A2(new_n585), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n391), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(G1gat), .ZN(G1324gat));
  INV_X1    g433(.A(new_n562), .ZN(new_n635));
  AOI21_X1  g434(.A(KEYINPUT88), .B1(new_n471), .B2(new_n474), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n631), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT103), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT42), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n639), .B1(new_n640), .B2(G8gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(KEYINPUT16), .B(G8gat), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n631), .A2(KEYINPUT42), .A3(new_n637), .A4(new_n643), .ZN(new_n644));
  OAI211_X1 g443(.A(new_n641), .B(new_n644), .C1(KEYINPUT42), .C2(new_n643), .ZN(G1325gat));
  NOR2_X1   g444(.A1(new_n538), .A2(new_n539), .ZN(new_n646));
  AOI21_X1  g445(.A(G15gat), .B1(new_n631), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n542), .A2(new_n543), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n631), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n647), .B1(G15gat), .B2(new_n649), .ZN(G1326gat));
  NAND2_X1  g449(.A1(new_n631), .A2(new_n509), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT43), .B(G22gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(G1327gat));
  INV_X1    g452(.A(KEYINPUT106), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n654), .B1(new_n578), .B2(new_n583), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n576), .A2(KEYINPUT35), .A3(new_n391), .A4(new_n475), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT35), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n389), .A2(new_n547), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n658), .B1(new_n635), .B2(new_n636), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n580), .A2(new_n572), .A3(new_n581), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n657), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n656), .A2(new_n661), .A3(KEYINPUT106), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n573), .A2(new_n510), .A3(new_n543), .A4(new_n542), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n655), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n665));
  AND3_X1   g464(.A1(new_n664), .A2(new_n665), .A3(new_n296), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT105), .ZN(new_n667));
  INV_X1    g466(.A(new_n296), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n668), .B1(new_n575), .B2(new_n584), .ZN(new_n669));
  OAI22_X1  g468(.A1(new_n666), .A2(new_n667), .B1(new_n669), .B2(new_n665), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n585), .A2(new_n296), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n671), .A2(KEYINPUT105), .A3(KEYINPUT44), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n250), .A2(new_n630), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(KEYINPUT107), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT107), .ZN(new_n677));
  AOI211_X1 g476(.A(new_n677), .B(new_n674), .C1(new_n670), .C2(new_n672), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(G29gat), .B1(new_n679), .B2(new_n391), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n671), .A2(new_n674), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n681), .A2(new_n251), .A3(new_n632), .ZN(new_n682));
  XOR2_X1   g481(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n680), .A2(new_n684), .ZN(G1328gat));
  INV_X1    g484(.A(new_n637), .ZN(new_n686));
  OAI21_X1  g485(.A(G36gat), .B1(new_n679), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n681), .A2(new_n252), .A3(new_n637), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT46), .Z(new_n689));
  NAND2_X1  g488(.A1(new_n687), .A2(new_n689), .ZN(G1329gat));
  NAND3_X1  g489(.A1(new_n664), .A2(new_n665), .A3(new_n296), .ZN(new_n691));
  AOI22_X1  g490(.A1(new_n671), .A2(KEYINPUT44), .B1(KEYINPUT105), .B2(new_n691), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n669), .A2(new_n667), .A3(new_n665), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n675), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n648), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n257), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n681), .A2(new_n262), .A3(new_n646), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n696), .A2(KEYINPUT47), .A3(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n697), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n648), .B1(new_n676), .B2(new_n678), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n699), .B1(new_n700), .B2(new_n257), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n698), .B1(new_n701), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n694), .A2(new_n677), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n673), .A2(KEYINPUT107), .A3(new_n675), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n572), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n703), .B1(new_n706), .B2(new_n258), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n681), .A2(new_n258), .A3(new_n509), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n509), .B1(new_n676), .B2(new_n678), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n709), .A2(KEYINPUT108), .A3(G50gat), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n707), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT48), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(G50gat), .B1(new_n694), .B2(new_n572), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n714), .A2(KEYINPUT48), .A3(new_n708), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(G1331gat));
  AND3_X1   g515(.A1(new_n297), .A2(new_n608), .A3(new_n664), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(new_n629), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n718), .A2(new_n391), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT109), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n214), .A2(new_n215), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(G1332gat));
  INV_X1    g521(.A(new_n718), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n686), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT110), .ZN(new_n726));
  NOR2_X1   g525(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n727));
  XOR2_X1   g526(.A(new_n726), .B(new_n727), .Z(G1333gat));
  NOR3_X1   g527(.A1(new_n718), .A2(new_n522), .A3(new_n695), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT111), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n723), .A2(new_n646), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n522), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g534(.A1(new_n723), .A2(new_n509), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g536(.A1(new_n249), .A2(new_n607), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n673), .A2(new_n629), .A3(new_n738), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n739), .A2(new_n275), .A3(new_n391), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n738), .A2(new_n296), .A3(new_n664), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT51), .ZN(new_n742));
  INV_X1    g541(.A(new_n629), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(G85gat), .B1(new_n744), .B2(new_n632), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n740), .A2(new_n745), .ZN(G1336gat));
  NAND2_X1  g545(.A1(new_n741), .A2(KEYINPUT112), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT51), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n686), .A2(G92gat), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n748), .A2(new_n629), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT113), .ZN(new_n751));
  INV_X1    g550(.A(new_n739), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n276), .B1(new_n752), .B2(new_n637), .ZN(new_n753));
  OAI21_X1  g552(.A(KEYINPUT52), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n744), .A2(new_n749), .ZN(new_n755));
  OR2_X1    g554(.A1(new_n755), .A2(KEYINPUT52), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n754), .B1(new_n753), .B2(new_n756), .ZN(G1337gat));
  XNOR2_X1  g556(.A(KEYINPUT114), .B(G99gat), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(new_n739), .B2(new_n695), .ZN(new_n759));
  INV_X1    g558(.A(new_n758), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n744), .A2(new_n646), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n761), .ZN(G1338gat));
  OAI21_X1  g561(.A(G106gat), .B1(new_n739), .B2(new_n572), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n572), .A2(G106gat), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT53), .B1(new_n744), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n748), .A2(new_n629), .A3(new_n764), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n766), .B1(new_n768), .B2(new_n769), .ZN(G1339gat));
  NOR2_X1   g569(.A1(new_n318), .A2(KEYINPUT118), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n594), .A2(new_n595), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n588), .B1(new_n587), .B2(new_n589), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n602), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n606), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n629), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT117), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n606), .A2(new_n774), .ZN(new_n778));
  OR3_X1    g577(.A1(new_n778), .A2(KEYINPUT117), .A3(new_n743), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n612), .A2(new_n613), .A3(new_n616), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n618), .A2(KEYINPUT54), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n614), .A2(new_n783), .A3(new_n617), .ZN(new_n784));
  AND3_X1   g583(.A1(new_n784), .A2(KEYINPUT115), .A3(new_n626), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT115), .B1(new_n784), .B2(new_n626), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n782), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI211_X1 g588(.A(KEYINPUT55), .B(new_n782), .C1(new_n785), .C2(new_n786), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n789), .A2(new_n628), .A3(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n608), .A2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n668), .B1(new_n780), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n296), .B1(new_n778), .B2(KEYINPUT116), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n778), .A2(KEYINPUT116), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n794), .A2(new_n795), .A3(new_n791), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n249), .B1(new_n793), .B2(new_n797), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n249), .A2(new_n668), .A3(new_n608), .A4(new_n743), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  OR2_X1    g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n801), .A2(new_n576), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n802), .A2(new_n632), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n686), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n771), .B1(new_n804), .B2(new_n608), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n803), .A2(new_n686), .ZN(new_n806));
  AOI22_X1  g605(.A1(new_n806), .A2(new_n607), .B1(KEYINPUT118), .B2(new_n318), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n805), .B1(new_n807), .B2(new_n771), .ZN(G1340gat));
  NOR2_X1   g607(.A1(new_n804), .A2(new_n743), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(new_n320), .ZN(G1341gat));
  NAND2_X1  g609(.A1(new_n806), .A2(new_n249), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(new_n352), .ZN(G1342gat));
  NAND3_X1  g611(.A1(new_n803), .A2(new_n296), .A3(new_n686), .ZN(new_n813));
  OR3_X1    g612(.A1(new_n813), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(G134gat), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT56), .B1(new_n813), .B2(G134gat), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(G1343gat));
  OAI21_X1  g616(.A(new_n509), .B1(new_n798), .B2(new_n800), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n648), .A2(new_n391), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n819), .A2(KEYINPUT121), .A3(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT121), .ZN(new_n822));
  INV_X1    g621(.A(new_n820), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n822), .B1(new_n818), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n637), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n608), .A2(G141gat), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT58), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT57), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n828), .B(new_n509), .C1(new_n798), .C2(new_n800), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n820), .A2(new_n686), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n791), .A2(KEYINPUT119), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n789), .A2(new_n833), .A3(new_n628), .A4(new_n790), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n832), .A2(new_n607), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n296), .B1(new_n835), .B2(new_n776), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n250), .B1(new_n836), .B2(new_n796), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n572), .B1(new_n837), .B2(new_n799), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n829), .B(new_n831), .C1(new_n828), .C2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(G141gat), .B1(new_n839), .B2(new_n608), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n827), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n819), .A2(new_n686), .A3(new_n820), .A4(new_n826), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n843), .A2(KEYINPUT120), .A3(KEYINPUT58), .ZN(new_n844));
  AOI21_X1  g643(.A(KEYINPUT120), .B1(new_n843), .B2(KEYINPUT58), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n841), .B1(new_n844), .B2(new_n845), .ZN(G1344gat));
  INV_X1    g645(.A(KEYINPUT122), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n791), .A2(KEYINPUT119), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n834), .A2(new_n607), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n776), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n796), .B1(new_n850), .B2(new_n668), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n847), .B(new_n799), .C1(new_n851), .C2(new_n249), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n847), .B1(new_n837), .B2(new_n799), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n828), .B(new_n509), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n818), .A2(KEYINPUT57), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n857), .A2(KEYINPUT59), .A3(new_n629), .A4(new_n831), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n859), .B1(new_n839), .B2(new_n743), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n304), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(G148gat), .B1(new_n825), .B2(new_n629), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n861), .B1(KEYINPUT59), .B2(new_n862), .ZN(G1345gat));
  NOR3_X1   g662(.A1(new_n839), .A2(new_n300), .A3(new_n250), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n825), .A2(new_n249), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n864), .B1(new_n865), .B2(new_n300), .ZN(G1346gat));
  NOR3_X1   g665(.A1(new_n839), .A2(new_n301), .A3(new_n668), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n825), .A2(new_n296), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n867), .B1(new_n868), .B2(new_n301), .ZN(G1347gat));
  NOR2_X1   g668(.A1(new_n686), .A2(new_n632), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n802), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n871), .A2(new_n608), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(new_n399), .ZN(G1348gat));
  NOR2_X1   g672(.A1(new_n871), .A2(new_n743), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n874), .B1(new_n401), .B2(new_n403), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n875), .B1(new_n402), .B2(new_n874), .ZN(G1349gat));
  OAI21_X1  g675(.A(G183gat), .B1(new_n871), .B2(new_n250), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT123), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n802), .A2(new_n249), .A3(new_n438), .A4(new_n870), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n880), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g680(.A1(new_n802), .A2(new_n296), .A3(new_n870), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n882), .A2(G190gat), .ZN(new_n883));
  XOR2_X1   g682(.A(KEYINPUT124), .B(KEYINPUT61), .Z(new_n884));
  OR2_X1    g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n882), .A2(G190gat), .A3(new_n884), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n885), .B(new_n886), .C1(G190gat), .C2(new_n882), .ZN(G1351gat));
  INV_X1    g686(.A(new_n870), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n818), .A2(new_n648), .A3(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(G197gat), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n889), .A2(new_n890), .A3(new_n607), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n888), .A2(new_n648), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n857), .A2(new_n892), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n893), .A2(new_n607), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n891), .B1(new_n894), .B2(new_n890), .ZN(G1352gat));
  INV_X1    g694(.A(G204gat), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n889), .A2(new_n896), .A3(new_n629), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT62), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n897), .B(new_n898), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n855), .A2(new_n629), .A3(new_n856), .A4(new_n892), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(G204gat), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT125), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n899), .A2(KEYINPUT125), .A3(new_n901), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(G1353gat));
  NAND3_X1  g705(.A1(new_n889), .A2(new_n203), .A3(new_n249), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n855), .A2(new_n249), .A3(new_n856), .A4(new_n892), .ZN(new_n908));
  AND3_X1   g707(.A1(new_n908), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n909));
  AOI21_X1  g708(.A(KEYINPUT63), .B1(new_n908), .B2(G211gat), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n907), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(KEYINPUT126), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT126), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n913), .B(new_n907), .C1(new_n909), .C2(new_n910), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n914), .ZN(G1354gat));
  AOI21_X1  g714(.A(G218gat), .B1(new_n889), .B2(new_n296), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n296), .A2(G218gat), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT127), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n916), .B1(new_n893), .B2(new_n918), .ZN(G1355gat));
endmodule


