//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 0 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 0 1 0 0 0 0 0 0 0 1 1 0 0 1 1 0 0 0 0 0 0 1 1 0 1 1 0 1 0 0 1 0 1 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n801, new_n802, new_n803, new_n804, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(G101), .ZN(new_n188));
  INV_X1    g002(.A(G107), .ZN(new_n189));
  AOI21_X1  g003(.A(KEYINPUT79), .B1(new_n189), .B2(G104), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n189), .A2(G104), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(KEYINPUT79), .A3(G104), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n188), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G104), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT3), .B1(new_n195), .B2(G107), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT3), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(new_n189), .A3(G104), .ZN(new_n198));
  AND2_X1   g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n188), .A2(KEYINPUT77), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT77), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G101), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n195), .A2(G107), .ZN(new_n203));
  AND3_X1   g017(.A1(new_n200), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT78), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n199), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n196), .A2(new_n198), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n200), .A2(new_n202), .A3(new_n203), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT78), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n194), .B1(new_n206), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G116), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(G119), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n214), .B1(new_n211), .B2(G119), .ZN(new_n215));
  INV_X1    g029(.A(G119), .ZN(new_n216));
  NOR3_X1   g030(.A1(new_n216), .A2(KEYINPUT66), .A3(G116), .ZN(new_n217));
  OAI211_X1 g031(.A(KEYINPUT5), .B(new_n213), .C1(new_n215), .C2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G113), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT5), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n219), .B1(new_n212), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT66), .B1(new_n216), .B2(G116), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n214), .A2(new_n211), .A3(G119), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n212), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n219), .A2(KEYINPUT2), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT2), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G113), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  AOI22_X1  g042(.A1(new_n218), .A2(new_n221), .B1(new_n224), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n210), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT4), .ZN(new_n231));
  AOI211_X1 g045(.A(new_n231), .B(new_n188), .C1(new_n199), .C2(new_n203), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n205), .B1(new_n199), .B2(new_n204), .ZN(new_n233));
  NOR3_X1   g047(.A1(new_n207), .A2(new_n208), .A3(KEYINPUT78), .ZN(new_n234));
  OAI21_X1  g048(.A(KEYINPUT4), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n188), .B1(new_n199), .B2(new_n203), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n232), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT67), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n222), .A2(new_n223), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n240), .A2(new_n213), .A3(new_n228), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n228), .B1(new_n240), .B2(new_n213), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n239), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n213), .B1(new_n215), .B2(new_n217), .ZN(new_n244));
  INV_X1    g058(.A(new_n228), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n224), .A2(new_n228), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n247), .A3(KEYINPUT67), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n243), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n230), .B1(new_n238), .B2(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(G110), .B(G122), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n230), .B(new_n251), .C1(new_n238), .C2(new_n249), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(KEYINPUT6), .A3(new_n254), .ZN(new_n255));
  AND2_X1   g069(.A1(KEYINPUT0), .A2(G128), .ZN(new_n256));
  NOR2_X1   g070(.A1(KEYINPUT0), .A2(G128), .ZN(new_n257));
  OR2_X1    g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G146), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT64), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(G143), .ZN(new_n261));
  INV_X1    g075(.A(G143), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n262), .A2(KEYINPUT64), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n259), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n259), .A2(G143), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n258), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n262), .A2(KEYINPUT64), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n260), .A2(G143), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n268), .A2(new_n269), .A3(G146), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n259), .A2(G143), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n270), .A2(new_n256), .A3(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(G125), .B1(new_n267), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT83), .ZN(new_n274));
  INV_X1    g088(.A(G128), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n275), .A2(KEYINPUT1), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n270), .A2(new_n271), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(G125), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n268), .A2(new_n269), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n265), .B1(new_n279), .B2(new_n259), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n275), .B1(new_n271), .B2(KEYINPUT1), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n277), .B(new_n278), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n273), .A2(new_n274), .A3(new_n282), .ZN(new_n283));
  OAI211_X1 g097(.A(KEYINPUT83), .B(G125), .C1(new_n267), .C2(new_n272), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G953), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(G224), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n285), .B(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT6), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n250), .A2(new_n289), .A3(new_n252), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n255), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n287), .A2(KEYINPUT7), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n283), .A2(new_n284), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT85), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT85), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n283), .A2(new_n295), .A3(new_n284), .A4(new_n292), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT86), .ZN(new_n298));
  XOR2_X1   g112(.A(new_n251), .B(KEYINPUT8), .Z(new_n299));
  NAND2_X1  g113(.A1(new_n206), .A2(new_n209), .ZN(new_n300));
  INV_X1    g114(.A(new_n194), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n229), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT84), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n299), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n303), .B1(new_n210), .B2(new_n229), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n301), .B1(new_n233), .B2(new_n234), .ZN(new_n306));
  INV_X1    g120(.A(new_n229), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n292), .ZN(new_n310));
  AOI22_X1  g124(.A1(new_n304), .A2(new_n309), .B1(new_n285), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n297), .A2(new_n298), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n254), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n298), .B1(new_n297), .B2(new_n311), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n187), .B(new_n291), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(G210), .B1(G237), .B2(G902), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(KEYINPUT87), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n297), .A2(new_n311), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT86), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(new_n254), .A3(new_n312), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n321), .A2(new_n187), .A3(new_n291), .A4(new_n316), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n318), .A2(KEYINPUT88), .A3(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT88), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n315), .A2(new_n324), .A3(new_n317), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(G214), .B1(G237), .B2(G902), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(KEYINPUT89), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT89), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n323), .A2(new_n330), .A3(new_n327), .A4(new_n325), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G217), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n333), .B1(G234), .B2(new_n187), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT25), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT22), .B(G137), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n286), .A2(G221), .A3(G234), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n337), .B(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT74), .ZN(new_n341));
  INV_X1    g155(.A(G140), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G125), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n278), .A2(G140), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(new_n344), .A3(KEYINPUT16), .ZN(new_n345));
  OR3_X1    g159(.A1(new_n278), .A2(KEYINPUT16), .A3(G140), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n341), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NOR3_X1   g161(.A1(new_n278), .A2(KEYINPUT16), .A3(G140), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n348), .A2(KEYINPUT74), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n259), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n349), .ZN(new_n351));
  XNOR2_X1  g165(.A(G125), .B(G140), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n348), .B1(new_n352), .B2(KEYINPUT16), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n351), .B(G146), .C1(new_n353), .C2(new_n341), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n350), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT23), .B1(new_n275), .B2(G119), .ZN(new_n356));
  AOI21_X1  g170(.A(KEYINPUT73), .B1(new_n275), .B2(G119), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n216), .A2(G128), .ZN(new_n358));
  OR2_X1    g172(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n359));
  AOI22_X1  g173(.A1(new_n356), .A2(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G110), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  XOR2_X1   g176(.A(G119), .B(G128), .Z(new_n363));
  XNOR2_X1  g177(.A(KEYINPUT24), .B(G110), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n355), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n360), .A2(new_n361), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n363), .A2(new_n364), .ZN(new_n369));
  AOI22_X1  g183(.A1(new_n368), .A2(new_n369), .B1(new_n259), .B2(new_n352), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n354), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n340), .B1(new_n367), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n367), .A2(new_n371), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT75), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT75), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n367), .A2(new_n375), .A3(new_n371), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n372), .B1(new_n377), .B2(new_n340), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n336), .B1(new_n378), .B2(G902), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n339), .B1(new_n374), .B2(new_n376), .ZN(new_n380));
  OAI211_X1 g194(.A(KEYINPUT25), .B(new_n187), .C1(new_n380), .C2(new_n372), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n335), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NOR3_X1   g196(.A1(new_n378), .A2(G902), .A3(new_n334), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NOR3_X1   g199(.A1(new_n241), .A2(new_n242), .A3(new_n239), .ZN(new_n386));
  AOI21_X1  g200(.A(KEYINPUT67), .B1(new_n246), .B2(new_n247), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n270), .A2(new_n256), .A3(new_n271), .ZN(new_n389));
  XNOR2_X1  g203(.A(KEYINPUT64), .B(G143), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n266), .B1(new_n390), .B2(G146), .ZN(new_n391));
  INV_X1    g205(.A(new_n258), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G131), .ZN(new_n394));
  INV_X1    g208(.A(G134), .ZN(new_n395));
  OAI21_X1  g209(.A(KEYINPUT65), .B1(new_n395), .B2(G137), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT11), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT11), .ZN(new_n398));
  OAI211_X1 g212(.A(KEYINPUT65), .B(new_n398), .C1(new_n395), .C2(G137), .ZN(new_n399));
  INV_X1    g213(.A(G137), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n400), .A2(G134), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  AND4_X1   g216(.A1(new_n394), .A2(new_n397), .A3(new_n399), .A4(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n401), .B1(new_n396), .B2(KEYINPUT11), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n394), .B1(new_n404), .B2(new_n399), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n389), .B(new_n393), .C1(new_n403), .C2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT30), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n404), .A2(new_n394), .A3(new_n399), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n395), .A2(G137), .ZN(new_n409));
  OAI21_X1  g223(.A(G131), .B1(new_n409), .B2(new_n401), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n281), .B1(new_n264), .B2(new_n266), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n270), .A2(new_n271), .A3(new_n276), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n408), .B(new_n410), .C1(new_n411), .C2(new_n412), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n406), .A2(new_n407), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n407), .B1(new_n406), .B2(new_n413), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n388), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n249), .A2(new_n406), .A3(new_n413), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT68), .ZN(new_n418));
  INV_X1    g232(.A(G237), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(KEYINPUT68), .A2(G237), .ZN(new_n421));
  AOI21_X1  g235(.A(G953), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(G210), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n423), .B(KEYINPUT27), .ZN(new_n424));
  XOR2_X1   g238(.A(KEYINPUT26), .B(G101), .Z(new_n425));
  XOR2_X1   g239(.A(new_n424), .B(new_n425), .Z(new_n426));
  NAND3_X1  g240(.A1(new_n416), .A2(new_n417), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT31), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n424), .B(new_n425), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT28), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n406), .A2(new_n413), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n388), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n430), .B1(new_n432), .B2(new_n417), .ZN(new_n433));
  INV_X1    g247(.A(new_n405), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n408), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n267), .A2(new_n272), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n408), .A2(new_n410), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n277), .B1(new_n280), .B2(new_n281), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n435), .A2(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(KEYINPUT28), .B1(new_n439), .B2(new_n249), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n429), .B1(new_n433), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n428), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n417), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n431), .A2(KEYINPUT30), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n406), .A2(new_n407), .A3(new_n413), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n443), .B1(new_n446), .B2(new_n388), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT69), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT31), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n447), .A2(new_n448), .A3(new_n449), .A4(new_n426), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n416), .A2(new_n449), .A3(new_n417), .A4(new_n426), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT69), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n442), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(G472), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n187), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT70), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT32), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n450), .A2(new_n452), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n432), .A2(new_n417), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT28), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n417), .A2(new_n430), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n462), .A2(new_n429), .B1(new_n427), .B2(KEYINPUT31), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n455), .B1(new_n458), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT70), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n456), .A2(new_n457), .A3(new_n466), .ZN(new_n467));
  NOR3_X1   g281(.A1(new_n433), .A2(new_n429), .A3(new_n440), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n426), .B1(new_n416), .B2(new_n417), .ZN(new_n469));
  NOR3_X1   g283(.A1(new_n468), .A2(new_n469), .A3(KEYINPUT29), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n440), .A2(KEYINPUT71), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT71), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n461), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT29), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n429), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n460), .A2(new_n471), .A3(new_n473), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n187), .ZN(new_n477));
  OAI21_X1  g291(.A(G472), .B1(new_n470), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(KEYINPUT72), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT72), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n480), .B(G472), .C1(new_n470), .C2(new_n477), .ZN(new_n481));
  AOI22_X1  g295(.A1(new_n479), .A2(new_n481), .B1(KEYINPUT32), .B2(new_n464), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n385), .B1(new_n467), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n438), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT80), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n306), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(KEYINPUT80), .B1(new_n210), .B2(new_n438), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n264), .A2(KEYINPUT1), .ZN(new_n488));
  AOI22_X1  g302(.A1(new_n488), .A2(G128), .B1(new_n271), .B2(new_n270), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n210), .B1(new_n489), .B2(new_n412), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n486), .A2(new_n487), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n435), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT12), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n493), .A2(KEYINPUT81), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(KEYINPUT81), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n492), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT10), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n484), .A2(new_n498), .ZN(new_n499));
  AOI22_X1  g313(.A1(new_n490), .A2(new_n498), .B1(new_n499), .B2(new_n210), .ZN(new_n500));
  INV_X1    g314(.A(new_n435), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n236), .A2(KEYINPUT4), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n231), .B1(new_n206), .B2(new_n209), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n502), .B1(new_n503), .B2(new_n236), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n436), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n500), .A2(new_n501), .A3(new_n505), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n491), .A2(KEYINPUT81), .A3(new_n493), .A4(new_n435), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n497), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(G110), .B(G140), .ZN(new_n509));
  INV_X1    g323(.A(G227), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n510), .A2(G953), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n509), .B(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n506), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n490), .A2(new_n498), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n499), .A2(new_n210), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n505), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n435), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n508), .A2(new_n512), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(G469), .B1(new_n519), .B2(G902), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT82), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI211_X1 g336(.A(KEYINPUT82), .B(G469), .C1(new_n519), .C2(G902), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n497), .A2(new_n506), .A3(new_n507), .A4(new_n513), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n517), .A2(new_n435), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n501), .B1(new_n500), .B2(new_n505), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n512), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AOI211_X1 g341(.A(G469), .B(G902), .C1(new_n524), .C2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n522), .A2(new_n523), .A3(new_n529), .ZN(new_n530));
  XNOR2_X1  g344(.A(KEYINPUT9), .B(G234), .ZN(new_n531));
  OAI21_X1  g345(.A(G221), .B1(new_n531), .B2(G902), .ZN(new_n532));
  XOR2_X1   g346(.A(new_n532), .B(KEYINPUT76), .Z(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT20), .ZN(new_n536));
  NOR2_X1   g350(.A1(G475), .A2(G902), .ZN(new_n537));
  XNOR2_X1  g351(.A(G113), .B(G122), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(new_n195), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n422), .A2(G143), .A3(G214), .ZN(new_n541));
  INV_X1    g355(.A(new_n421), .ZN(new_n542));
  NOR2_X1   g356(.A1(KEYINPUT68), .A2(G237), .ZN(new_n543));
  OAI211_X1 g357(.A(G214), .B(new_n286), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n390), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n394), .B1(new_n541), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT18), .ZN(new_n547));
  NAND2_X1  g361(.A1(KEYINPUT18), .A2(G131), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n541), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n352), .B(new_n259), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n355), .B1(KEYINPUT17), .B2(new_n546), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n541), .A2(new_n545), .A3(new_n394), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT91), .ZN(new_n554));
  INV_X1    g368(.A(new_n546), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT17), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT91), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n541), .A2(new_n545), .A3(new_n557), .A4(new_n394), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n554), .A2(new_n555), .A3(new_n556), .A4(new_n558), .ZN(new_n559));
  AOI221_X4 g373(.A(new_n540), .B1(new_n547), .B2(new_n551), .C1(new_n552), .C2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n554), .A2(new_n555), .A3(new_n558), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n352), .B(KEYINPUT19), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n259), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n561), .A2(new_n354), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n551), .A2(new_n547), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n539), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n536), .B(new_n537), .C1(new_n560), .C2(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n537), .B1(new_n560), .B2(new_n566), .ZN(new_n568));
  XNOR2_X1  g382(.A(KEYINPUT90), .B(KEYINPUT20), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n567), .A2(KEYINPUT92), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n566), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n552), .A2(new_n559), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(new_n539), .A3(new_n565), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT92), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n575), .A2(new_n576), .A3(new_n536), .A4(new_n537), .ZN(new_n577));
  INV_X1    g391(.A(G475), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n539), .B1(new_n573), .B2(new_n565), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n187), .B1(new_n560), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n578), .B1(new_n580), .B2(KEYINPUT93), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT93), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n582), .B(new_n187), .C1(new_n560), .C2(new_n579), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n571), .A2(new_n577), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(G234), .A2(G237), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n585), .A2(G952), .A3(new_n286), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n585), .A2(G902), .A3(G953), .ZN(new_n587));
  XNOR2_X1  g401(.A(KEYINPUT21), .B(G898), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT96), .ZN(new_n591));
  XNOR2_X1  g405(.A(KEYINPUT94), .B(G122), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(G116), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT95), .ZN(new_n594));
  INV_X1    g408(.A(G122), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n594), .B1(new_n595), .B2(G116), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n211), .A2(KEYINPUT95), .A3(G122), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n593), .A2(new_n189), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n268), .A2(new_n269), .A3(G128), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n275), .A2(G143), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n600), .A2(new_n395), .A3(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n395), .B1(new_n600), .B2(new_n601), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n599), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g419(.A1(new_n598), .A2(KEYINPUT14), .B1(new_n592), .B2(G116), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT14), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n596), .A2(new_n607), .A3(new_n597), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n189), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n591), .B1(new_n605), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n598), .A2(KEYINPUT14), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n611), .A2(new_n608), .A3(new_n593), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(G107), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n600), .A2(new_n601), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(G134), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n602), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n613), .A2(new_n616), .A3(KEYINPUT96), .A4(new_n599), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n600), .A2(KEYINPUT13), .A3(new_n601), .ZN(new_n618));
  OAI211_X1 g432(.A(new_n618), .B(G134), .C1(KEYINPUT13), .C2(new_n600), .ZN(new_n619));
  INV_X1    g433(.A(new_n599), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n189), .B1(new_n593), .B2(new_n598), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n619), .B(new_n602), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n610), .A2(new_n617), .A3(new_n622), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n531), .A2(new_n333), .A3(G953), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n610), .A2(new_n617), .A3(new_n622), .A4(new_n624), .ZN(new_n627));
  AOI21_X1  g441(.A(G902), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(G478), .ZN(new_n629));
  OR2_X1    g443(.A1(new_n629), .A2(KEYINPUT15), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n628), .B(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n584), .A2(new_n590), .A3(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n535), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n332), .A2(new_n483), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n200), .A2(new_n202), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G3));
  INV_X1    g451(.A(new_n316), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n315), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n328), .B1(new_n639), .B2(new_n322), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n640), .A2(KEYINPUT98), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT98), .ZN(new_n642));
  AOI211_X1 g456(.A(new_n642), .B(new_n328), .C1(new_n639), .C2(new_n322), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n567), .A2(KEYINPUT92), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n568), .A2(new_n570), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n577), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n580), .A2(KEYINPUT93), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n647), .A2(G475), .A3(new_n583), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n626), .A2(new_n627), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(KEYINPUT33), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT33), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n626), .A2(new_n652), .A3(new_n627), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n651), .A2(G478), .A3(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT99), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n629), .A2(new_n187), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n656), .B1(new_n628), .B2(new_n629), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n654), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n655), .B1(new_n654), .B2(new_n657), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n649), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NOR4_X1   g474(.A1(new_n641), .A2(new_n643), .A3(new_n589), .A4(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n458), .A2(new_n463), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n187), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT97), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n663), .A2(new_n664), .A3(G472), .ZN(new_n665));
  AOI21_X1  g479(.A(G902), .B1(new_n458), .B2(new_n463), .ZN(new_n666));
  OAI21_X1  g480(.A(KEYINPUT97), .B1(new_n666), .B2(new_n454), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n464), .B(KEYINPUT70), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n668), .A2(new_n669), .A3(new_n384), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(new_n535), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n661), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT34), .B(G104), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G6));
  INV_X1    g488(.A(KEYINPUT102), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n641), .A2(new_n643), .A3(new_n589), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n575), .A2(new_n537), .A3(new_n569), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n645), .A2(new_n677), .A3(KEYINPUT100), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT100), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n575), .A2(new_n679), .A3(new_n537), .A4(new_n569), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n678), .A2(new_n631), .A3(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT101), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n648), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(KEYINPUT101), .B1(new_n581), .B2(new_n583), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n681), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n675), .B1(new_n676), .B2(new_n685), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n291), .A2(new_n187), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n316), .B1(new_n687), .B2(new_n321), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n315), .A2(new_n638), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n327), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n642), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n640), .A2(KEYINPUT98), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n691), .A2(new_n590), .A3(new_n692), .A4(new_n685), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n693), .A2(KEYINPUT102), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n671), .B1(new_n686), .B2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT103), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT35), .B(G107), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G9));
  NAND2_X1  g512(.A1(new_n668), .A2(new_n669), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n379), .A2(new_n381), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n334), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n340), .A2(KEYINPUT36), .ZN(new_n702));
  XOR2_X1   g516(.A(new_n377), .B(new_n702), .Z(new_n703));
  NAND3_X1  g517(.A1(new_n703), .A2(new_n187), .A3(new_n335), .ZN(new_n704));
  AND2_X1   g518(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n699), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n332), .A2(new_n634), .A3(new_n706), .ZN(new_n707));
  XOR2_X1   g521(.A(KEYINPUT37), .B(G110), .Z(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G12));
  NOR2_X1   g523(.A1(new_n641), .A2(new_n643), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n528), .B1(new_n520), .B2(new_n521), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n533), .B1(new_n711), .B2(new_n523), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n705), .B1(new_n467), .B2(new_n482), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n648), .B(new_n682), .ZN(new_n714));
  INV_X1    g528(.A(G900), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n587), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n586), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n714), .A2(new_n681), .A3(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n710), .A2(new_n712), .A3(new_n713), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G128), .ZN(G30));
  XNOR2_X1  g536(.A(new_n718), .B(KEYINPUT39), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n712), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(KEYINPUT40), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT106), .ZN(new_n726));
  OR2_X1    g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n725), .A2(new_n726), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n464), .A2(KEYINPUT32), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n447), .A2(new_n429), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n187), .B1(new_n459), .B2(new_n426), .ZN(new_n731));
  OAI21_X1  g545(.A(G472), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n467), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n649), .A2(new_n631), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n701), .A2(new_n704), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n735), .A2(new_n736), .A3(new_n328), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n734), .B1(new_n737), .B2(KEYINPUT105), .ZN(new_n738));
  XOR2_X1   g552(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n739));
  XNOR2_X1  g553(.A(new_n326), .B(new_n739), .ZN(new_n740));
  AOI211_X1 g554(.A(new_n738), .B(new_n740), .C1(KEYINPUT105), .C2(new_n737), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n727), .A2(new_n728), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(new_n279), .ZN(G45));
  NOR2_X1   g557(.A1(new_n658), .A2(new_n659), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n744), .A2(new_n584), .A3(new_n719), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n710), .A2(new_n712), .A3(new_n713), .A4(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G146), .ZN(G48));
  INV_X1    g561(.A(KEYINPUT108), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n467), .A2(new_n482), .ZN(new_n749));
  AOI21_X1  g563(.A(G902), .B1(new_n524), .B2(new_n527), .ZN(new_n750));
  INV_X1    g564(.A(G469), .ZN(new_n751));
  AOI21_X1  g565(.A(KEYINPUT107), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n513), .B1(new_n518), .B2(new_n506), .ZN(new_n753));
  INV_X1    g567(.A(new_n496), .ZN(new_n754));
  AOI211_X1 g568(.A(new_n494), .B(new_n754), .C1(new_n491), .C2(new_n435), .ZN(new_n755));
  INV_X1    g569(.A(new_n507), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n753), .B1(new_n757), .B2(new_n514), .ZN(new_n758));
  OAI21_X1  g572(.A(G469), .B1(new_n758), .B2(G902), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n752), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT107), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n750), .A2(new_n761), .A3(new_n751), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n533), .B1(new_n760), .B2(new_n763), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n749), .A2(new_n384), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n748), .B1(new_n661), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n744), .A2(new_n584), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n691), .A2(new_n590), .A3(new_n767), .A4(new_n692), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n749), .A2(new_n384), .A3(new_n764), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n768), .A2(new_n769), .A3(KEYINPUT108), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  XOR2_X1   g585(.A(KEYINPUT41), .B(G113), .Z(new_n772));
  XNOR2_X1  g586(.A(new_n771), .B(new_n772), .ZN(G15));
  OAI21_X1  g587(.A(new_n765), .B1(new_n686), .B2(new_n694), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT109), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT109), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n776), .B(new_n765), .C1(new_n686), .C2(new_n694), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  XOR2_X1   g592(.A(KEYINPUT110), .B(G116), .Z(new_n779));
  XNOR2_X1  g593(.A(new_n778), .B(new_n779), .ZN(G18));
  NOR2_X1   g594(.A1(new_n750), .A2(new_n751), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n781), .A2(new_n528), .A3(KEYINPUT107), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n534), .B1(new_n782), .B2(new_n762), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n783), .A2(new_n641), .A3(new_n643), .ZN(new_n784));
  AOI211_X1 g598(.A(new_n705), .B(new_n633), .C1(new_n467), .C2(new_n482), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G119), .ZN(G21));
  NOR3_X1   g601(.A1(new_n641), .A2(new_n643), .A3(new_n735), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n460), .A2(new_n471), .A3(new_n473), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT111), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n429), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n789), .A2(new_n790), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n458), .B(new_n428), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n794), .A2(new_n454), .A3(new_n187), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n663), .A2(G472), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n795), .A2(new_n796), .A3(new_n384), .A4(new_n590), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n783), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n788), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G122), .ZN(G24));
  INV_X1    g614(.A(new_n745), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n795), .A2(new_n796), .A3(new_n736), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n784), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G125), .ZN(G27));
  AOI21_X1  g619(.A(new_n328), .B1(new_n323), .B2(new_n325), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n533), .B1(new_n529), .B2(new_n520), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n806), .A2(new_n745), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n479), .A2(new_n481), .ZN(new_n809));
  OAI211_X1 g623(.A(KEYINPUT112), .B(new_n457), .C1(new_n453), .C2(new_n455), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT112), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n811), .B1(new_n464), .B2(KEYINPUT32), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n809), .A2(new_n810), .A3(new_n729), .A4(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT113), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n813), .A2(new_n814), .A3(new_n384), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n814), .B1(new_n813), .B2(new_n384), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n808), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT42), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n483), .A2(new_n806), .A3(new_n807), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT42), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n819), .A2(new_n820), .A3(new_n745), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(new_n394), .ZN(G33));
  NAND2_X1  g637(.A1(new_n819), .A2(new_n720), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(G134), .ZN(G36));
  INV_X1    g639(.A(new_n744), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n584), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT43), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n829), .A2(new_n699), .A3(new_n736), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT44), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n519), .A2(KEYINPUT45), .ZN(new_n833));
  OAI21_X1  g647(.A(G469), .B1(new_n519), .B2(KEYINPUT45), .ZN(new_n834));
  OAI22_X1  g648(.A1(new_n833), .A2(new_n834), .B1(new_n751), .B2(new_n187), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT46), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n528), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n837), .B1(new_n836), .B2(new_n835), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n838), .A2(new_n534), .A3(new_n723), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n832), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n830), .A2(new_n831), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(new_n806), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT114), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n842), .A2(KEYINPUT114), .A3(new_n806), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n841), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(new_n400), .ZN(G39));
  AND3_X1   g662(.A1(new_n838), .A2(KEYINPUT47), .A3(new_n534), .ZN(new_n849));
  AOI21_X1  g663(.A(KEYINPUT47), .B1(new_n838), .B2(new_n534), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n806), .ZN(new_n853));
  NOR4_X1   g667(.A1(new_n853), .A2(new_n801), .A3(new_n749), .A4(new_n384), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT115), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n855), .B(new_n856), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(G140), .ZN(G42));
  NOR4_X1   g672(.A1(new_n827), .A2(new_n385), .A3(new_n328), .A4(new_n533), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT49), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n760), .A2(new_n763), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(KEYINPUT116), .ZN(new_n863));
  INV_X1    g677(.A(new_n734), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n861), .A2(new_n860), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT117), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n863), .A2(new_n864), .A3(new_n740), .A4(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n736), .A2(new_n719), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n788), .A2(new_n734), .A3(new_n807), .A4(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n869), .A2(new_n804), .A3(new_n721), .A4(new_n746), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT52), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n784), .A2(new_n785), .B1(new_n788), .B2(new_n798), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n649), .A2(new_n632), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n767), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n874), .A2(new_n589), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n332), .A2(new_n671), .A3(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n872), .A2(new_n707), .A3(new_n635), .A4(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n877), .A2(new_n771), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n678), .A2(new_n632), .A3(new_n680), .A4(new_n718), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n714), .A2(new_n879), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n712), .A2(new_n880), .A3(new_n806), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n806), .A2(new_n807), .ZN(new_n882));
  AOI22_X1  g696(.A1(new_n881), .A2(new_n713), .B1(new_n803), .B2(new_n882), .ZN(new_n883));
  AND4_X1   g697(.A1(new_n818), .A2(new_n821), .A3(new_n824), .A4(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n778), .A2(new_n878), .A3(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT118), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n871), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n778), .A2(new_n878), .A3(new_n884), .A4(KEYINPUT118), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n887), .A2(KEYINPUT53), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT53), .B1(new_n887), .B2(new_n888), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n889), .B1(new_n890), .B2(KEYINPUT119), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT119), .ZN(new_n892));
  AOI211_X1 g706(.A(new_n892), .B(KEYINPUT53), .C1(new_n887), .C2(new_n888), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT54), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n890), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT54), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT53), .ZN(new_n897));
  OR2_X1    g711(.A1(new_n871), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n898), .A2(new_n885), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n895), .A2(new_n896), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n894), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n829), .A2(new_n586), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n795), .A2(new_n796), .A3(new_n384), .ZN(new_n904));
  OR2_X1    g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n740), .A2(new_n328), .A3(new_n764), .ZN(new_n906));
  OAI21_X1  g720(.A(KEYINPUT120), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT50), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n907), .A2(new_n908), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n806), .A2(new_n764), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n903), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n802), .ZN(new_n913));
  NOR4_X1   g727(.A1(new_n911), .A2(new_n734), .A3(new_n385), .A4(new_n717), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n826), .A2(new_n649), .ZN(new_n915));
  AOI22_X1  g729(.A1(new_n912), .A2(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n909), .A2(new_n910), .A3(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT51), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n861), .A2(new_n533), .ZN(new_n919));
  AOI211_X1 g733(.A(new_n853), .B(new_n905), .C1(new_n851), .C2(new_n919), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n917), .A2(new_n918), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n918), .B1(new_n917), .B2(new_n920), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n912), .B1(new_n815), .B2(new_n816), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT48), .Z(new_n924));
  INV_X1    g738(.A(G952), .ZN(new_n925));
  AOI211_X1 g739(.A(new_n925), .B(G953), .C1(new_n914), .C2(new_n767), .ZN(new_n926));
  INV_X1    g740(.A(new_n784), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n926), .B1(new_n905), .B2(new_n927), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n928), .A2(KEYINPUT121), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n928), .A2(KEYINPUT121), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n924), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n922), .A2(new_n931), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n902), .A2(new_n921), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n925), .A2(new_n286), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT122), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n867), .B1(new_n933), .B2(new_n935), .ZN(G75));
  NOR2_X1   g750(.A1(new_n286), .A2(G952), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n255), .A2(new_n290), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT123), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT55), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(new_n288), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n890), .A2(new_n899), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n942), .A2(new_n187), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(G210), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT56), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n941), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n943), .A2(new_n317), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n941), .A2(new_n945), .ZN(new_n948));
  AOI211_X1 g762(.A(new_n937), .B(new_n946), .C1(new_n947), .C2(new_n948), .ZN(G51));
  INV_X1    g763(.A(new_n758), .ZN(new_n950));
  OAI21_X1  g764(.A(KEYINPUT54), .B1(new_n890), .B2(new_n899), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n901), .A2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n751), .A2(new_n187), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT57), .Z(new_n955));
  OAI21_X1  g769(.A(new_n950), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n833), .A2(new_n834), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n943), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n937), .B1(new_n956), .B2(new_n958), .ZN(G54));
  NAND3_X1  g773(.A1(new_n943), .A2(KEYINPUT58), .A3(G475), .ZN(new_n960));
  INV_X1    g774(.A(new_n575), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n960), .A2(new_n961), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n962), .A2(new_n963), .A3(new_n937), .ZN(G60));
  XNOR2_X1  g778(.A(new_n656), .B(KEYINPUT59), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n965), .B1(new_n651), .B2(new_n653), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n937), .B1(new_n952), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n965), .B1(new_n894), .B2(new_n901), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n651), .A2(new_n653), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT124), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI211_X1 g786(.A(KEYINPUT124), .B(new_n967), .C1(new_n968), .C2(new_n969), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(G63));
  NAND2_X1  g788(.A1(G217), .A2(G902), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT60), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n942), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n703), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n378), .B1(new_n942), .B2(new_n976), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n978), .B(new_n979), .C1(G952), .C2(new_n286), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT61), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n980), .B(new_n981), .ZN(G66));
  INV_X1    g796(.A(G224), .ZN(new_n983));
  OAI21_X1  g797(.A(G953), .B1(new_n588), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n778), .A2(new_n878), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n984), .B1(new_n986), .B2(G953), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n939), .B1(G898), .B2(new_n286), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(G69));
  NAND2_X1  g803(.A1(new_n845), .A2(new_n846), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n840), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n804), .A2(new_n721), .A3(new_n746), .ZN(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n991), .A2(KEYINPUT126), .A3(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT126), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n995), .B1(new_n847), .B2(new_n992), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n822), .B1(new_n720), .B2(new_n819), .ZN(new_n998));
  INV_X1    g812(.A(new_n839), .ZN(new_n999));
  OAI211_X1 g813(.A(new_n999), .B(new_n788), .C1(new_n815), .C2(new_n816), .ZN(new_n1000));
  AND3_X1   g814(.A1(new_n857), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n997), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(new_n286), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n286), .A2(G900), .ZN(new_n1004));
  INV_X1    g818(.A(new_n1004), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1003), .A2(KEYINPUT127), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT127), .ZN(new_n1007));
  AOI21_X1  g821(.A(G953), .B1(new_n997), .B2(new_n1001), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1007), .B1(new_n1008), .B2(new_n1004), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  XOR2_X1   g824(.A(new_n562), .B(KEYINPUT125), .Z(new_n1011));
  XNOR2_X1  g825(.A(new_n446), .B(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  OAI211_X1 g827(.A(new_n483), .B(new_n806), .C1(new_n767), .C2(new_n873), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n1014), .A2(new_n724), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n847), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n742), .A2(new_n993), .ZN(new_n1017));
  OR2_X1    g831(.A1(new_n1017), .A2(KEYINPUT62), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1017), .A2(KEYINPUT62), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n1016), .A2(new_n1018), .A3(new_n857), .A4(new_n1019), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n1012), .A2(G953), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g836(.A(G953), .B1(new_n510), .B2(new_n715), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1023), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1013), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(new_n1012), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1026), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1027));
  INV_X1    g841(.A(new_n1022), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1023), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1025), .A2(new_n1029), .ZN(G72));
  NAND2_X1  g844(.A1(G472), .A2(G902), .ZN(new_n1031));
  XOR2_X1   g845(.A(new_n1031), .B(KEYINPUT63), .Z(new_n1032));
  OAI21_X1  g846(.A(new_n1032), .B1(new_n1002), .B2(new_n985), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n1033), .A2(new_n447), .A3(new_n429), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1032), .B1(new_n1020), .B2(new_n985), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n937), .B1(new_n1035), .B2(new_n730), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  OR2_X1    g851(.A1(new_n891), .A2(new_n893), .ZN(new_n1038));
  INV_X1    g852(.A(new_n1032), .ZN(new_n1039));
  OR2_X1    g853(.A1(new_n447), .A2(new_n426), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n1039), .B1(new_n1040), .B2(new_n427), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n1037), .B1(new_n1038), .B2(new_n1041), .ZN(G57));
endmodule


