//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 0 0 1 0 1 1 0 1 0 0 0 0 0 1 1 0 0 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 0 0 0 1 0 0 1 0 0 1 1 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010;
  INV_X1    g000(.A(G104), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT3), .B1(new_n187), .B2(G107), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G104), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n187), .A2(G107), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n188), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT77), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT77), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n188), .A2(new_n191), .A3(new_n195), .A4(new_n192), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(G101), .A3(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G101), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n188), .A2(new_n191), .A3(new_n198), .A4(new_n192), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n197), .A2(KEYINPUT4), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT64), .ZN(new_n201));
  XNOR2_X1  g015(.A(G143), .B(G146), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT0), .B(G128), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n201), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  AND2_X1   g018(.A1(KEYINPUT0), .A2(G128), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n202), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G143), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(KEYINPUT0), .A2(G128), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n205), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n211), .A2(new_n213), .A3(KEYINPUT64), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n204), .A2(new_n206), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT78), .B(KEYINPUT4), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n194), .A2(G101), .A3(new_n196), .A4(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n200), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n190), .A2(G104), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n187), .A2(G107), .ZN(new_n221));
  OAI21_X1  g035(.A(G101), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n199), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n224), .B(KEYINPUT1), .C1(new_n209), .C2(G146), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G128), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n224), .B1(new_n208), .B2(KEYINPUT1), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n211), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT1), .ZN(new_n229));
  AND4_X1   g043(.A1(new_n229), .A2(new_n208), .A3(new_n210), .A4(G128), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n223), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT1), .B1(new_n209), .B2(G146), .ZN(new_n233));
  AOI22_X1  g047(.A1(new_n233), .A2(G128), .B1(new_n208), .B2(new_n210), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n199), .B(new_n222), .C1(new_n230), .C2(new_n234), .ZN(new_n235));
  XOR2_X1   g049(.A(KEYINPUT79), .B(KEYINPUT10), .Z(new_n236));
  AOI22_X1  g050(.A1(new_n232), .A2(KEYINPUT10), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT11), .ZN(new_n238));
  INV_X1    g052(.A(G134), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n238), .B1(new_n239), .B2(G137), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(G137), .ZN(new_n241));
  INV_X1    g055(.A(G137), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(KEYINPUT11), .A3(G134), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n240), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G131), .ZN(new_n245));
  INV_X1    g059(.A(G131), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n240), .A2(new_n243), .A3(new_n246), .A4(new_n241), .ZN(new_n247));
  AND2_X1   g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n219), .A2(new_n237), .A3(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(G110), .B(G140), .ZN(new_n250));
  INV_X1    g064(.A(G953), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n251), .A2(G227), .ZN(new_n252));
  XOR2_X1   g066(.A(new_n250), .B(new_n252), .Z(new_n253));
  AND2_X1   g067(.A1(new_n249), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n219), .A2(new_n237), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n245), .A2(new_n247), .ZN(new_n256));
  AOI21_X1  g070(.A(KEYINPUT80), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT80), .ZN(new_n258));
  AOI211_X1 g072(.A(new_n258), .B(new_n248), .C1(new_n219), .C2(new_n237), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n254), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n253), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n228), .A2(new_n231), .ZN(new_n262));
  INV_X1    g076(.A(new_n223), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n235), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  AND3_X1   g078(.A1(new_n264), .A2(KEYINPUT12), .A3(new_n256), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT12), .B1(new_n264), .B2(new_n256), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n249), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n261), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n260), .A2(KEYINPUT81), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT81), .B1(new_n260), .B2(new_n269), .ZN(new_n271));
  OAI21_X1  g085(.A(G469), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G469), .ZN(new_n273));
  INV_X1    g087(.A(G902), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n248), .B1(new_n219), .B2(new_n237), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n275), .B(KEYINPUT80), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n253), .B1(new_n276), .B2(new_n249), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n249), .A2(new_n253), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n278), .A2(new_n267), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n273), .B(new_n274), .C1(new_n277), .C2(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n273), .A2(new_n274), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n272), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(G214), .B1(G237), .B2(G902), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(G210), .B1(G237), .B2(G902), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n215), .A2(G125), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n288), .B1(G125), .B2(new_n262), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n251), .A2(G224), .ZN(new_n290));
  XOR2_X1   g104(.A(new_n289), .B(new_n290), .Z(new_n291));
  XOR2_X1   g105(.A(G110), .B(G122), .Z(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  XNOR2_X1  g107(.A(KEYINPUT2), .B(G113), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G119), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n296), .A2(G116), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT68), .B(G119), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n297), .B1(new_n298), .B2(G116), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT67), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n295), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  AND2_X1   g115(.A1(KEYINPUT68), .A2(G119), .ZN(new_n302));
  NOR2_X1   g116(.A1(KEYINPUT68), .A2(G119), .ZN(new_n303));
  OAI21_X1  g117(.A(G116), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n297), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n306), .A2(KEYINPUT67), .A3(new_n294), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n301), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n200), .A2(new_n308), .A3(new_n218), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT5), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n298), .A2(new_n310), .A3(G116), .ZN(new_n311));
  OAI211_X1 g125(.A(G113), .B(new_n311), .C1(new_n306), .C2(new_n310), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n299), .A2(new_n295), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(new_n263), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n293), .B1(new_n309), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n309), .A2(new_n314), .A3(new_n293), .ZN(new_n316));
  NAND2_X1  g130(.A1(KEYINPUT82), .A2(KEYINPUT6), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n315), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  AOI211_X1 g133(.A(new_n293), .B(new_n317), .C1(new_n309), .C2(new_n314), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n291), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n274), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n290), .A2(KEYINPUT7), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n289), .B(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n312), .A2(new_n313), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT83), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT83), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n312), .A2(new_n328), .A3(new_n313), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n263), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT84), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n223), .B1(new_n327), .B2(new_n329), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n326), .A2(new_n223), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(KEYINPUT84), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n333), .A2(new_n337), .A3(new_n316), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n292), .B(KEYINPUT8), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n316), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n325), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n287), .B1(new_n322), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n332), .B1(new_n331), .B2(new_n335), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n316), .B1(new_n334), .B2(KEYINPUT84), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n340), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n324), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n346), .A2(new_n274), .A3(new_n286), .A4(new_n321), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n285), .B1(new_n342), .B2(new_n347), .ZN(new_n348));
  XOR2_X1   g162(.A(KEYINPUT9), .B(G234), .Z(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(G221), .B1(new_n350), .B2(G902), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n283), .A2(new_n348), .A3(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(G128), .B(G143), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n239), .B1(new_n353), .B2(KEYINPUT13), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n209), .A2(G128), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n354), .B1(KEYINPUT13), .B2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n356), .B(KEYINPUT91), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n353), .A2(new_n239), .ZN(new_n358));
  AND2_X1   g172(.A1(KEYINPUT89), .A2(G122), .ZN(new_n359));
  NOR2_X1   g173(.A1(KEYINPUT89), .A2(G122), .ZN(new_n360));
  OAI21_X1  g174(.A(G116), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT90), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT90), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n363), .B(G116), .C1(new_n359), .C2(new_n360), .ZN(new_n364));
  INV_X1    g178(.A(G116), .ZN(new_n365));
  AOI22_X1  g179(.A1(new_n362), .A2(new_n364), .B1(new_n365), .B2(G122), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n366), .A2(new_n190), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n366), .A2(new_n190), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n357), .B(new_n358), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G217), .ZN(new_n370));
  NOR3_X1   g184(.A1(new_n350), .A2(new_n370), .A3(G953), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n362), .A2(new_n364), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n365), .A2(G122), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n373), .B(KEYINPUT14), .ZN(new_n374));
  OAI21_X1  g188(.A(G107), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT92), .ZN(new_n376));
  OR2_X1    g190(.A1(new_n353), .A2(new_n239), .ZN(new_n377));
  AOI22_X1  g191(.A1(new_n366), .A2(new_n190), .B1(new_n358), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT92), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n379), .B(G107), .C1(new_n372), .C2(new_n374), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n376), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n369), .A2(new_n371), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n371), .B1(new_n369), .B2(new_n381), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n274), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT15), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n385), .A3(G478), .ZN(new_n386));
  INV_X1    g200(.A(G478), .ZN(new_n387));
  OAI221_X1 g201(.A(new_n274), .B1(KEYINPUT15), .B2(new_n387), .C1(new_n382), .C2(new_n383), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT20), .ZN(new_n391));
  OR2_X1    g205(.A1(G475), .A2(G902), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT16), .ZN(new_n393));
  INV_X1    g207(.A(G125), .ZN(new_n394));
  INV_X1    g208(.A(G140), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(G125), .A2(G140), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n393), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n393), .A2(new_n395), .A3(G125), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n207), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n397), .ZN(new_n402));
  NOR2_X1   g216(.A1(G125), .A2(G140), .ZN(new_n403));
  OAI21_X1  g217(.A(KEYINPUT16), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(G146), .A3(new_n399), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n401), .A2(KEYINPUT75), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT75), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n404), .A2(new_n407), .A3(G146), .A4(new_n399), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT17), .ZN(new_n410));
  INV_X1    g224(.A(G237), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(new_n251), .A3(G214), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT85), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n412), .A2(new_n413), .A3(new_n209), .ZN(new_n414));
  NOR2_X1   g228(.A1(G237), .A2(G953), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n415), .B(G214), .C1(KEYINPUT85), .C2(G143), .ZN(new_n416));
  AOI211_X1 g230(.A(new_n410), .B(new_n246), .C1(new_n414), .C2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n409), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT87), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n414), .A2(new_n416), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n246), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n422), .A2(G131), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(new_n410), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n409), .A2(KEYINPUT87), .A3(new_n418), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n421), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(G113), .B(G122), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n429), .B(new_n187), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT18), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n423), .B1(new_n431), .B2(new_n246), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n396), .A2(new_n397), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n433), .B(new_n207), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n425), .A2(new_n431), .ZN(new_n436));
  OR2_X1    g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n428), .A2(new_n430), .A3(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT19), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n433), .B(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n405), .B1(new_n440), .B2(G146), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT86), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n424), .A2(new_n425), .ZN(new_n444));
  OAI211_X1 g258(.A(KEYINPUT86), .B(new_n405), .C1(new_n440), .C2(G146), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n437), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n430), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n392), .B1(new_n438), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n391), .B1(new_n450), .B2(KEYINPUT88), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT88), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n430), .B1(new_n437), .B2(new_n446), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n435), .A2(new_n436), .ZN(new_n454));
  AOI211_X1 g268(.A(new_n420), .B(new_n417), .C1(new_n408), .C2(new_n406), .ZN(new_n455));
  AOI21_X1  g269(.A(KEYINPUT87), .B1(new_n409), .B2(new_n418), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n454), .B1(new_n457), .B2(new_n426), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n453), .B1(new_n458), .B2(new_n430), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n452), .B1(new_n459), .B2(new_n392), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n451), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n428), .A2(new_n437), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(new_n430), .ZN(new_n463));
  OAI21_X1  g277(.A(G475), .B1(new_n463), .B2(G902), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n452), .B(new_n391), .C1(new_n459), .C2(new_n392), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n390), .A2(new_n461), .A3(new_n464), .A4(new_n465), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n251), .A2(G952), .ZN(new_n467));
  NAND2_X1  g281(.A1(G234), .A2(G237), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  XOR2_X1   g284(.A(KEYINPUT21), .B(G898), .Z(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n468), .A2(G902), .A3(G953), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n470), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(KEYINPUT93), .B1(new_n466), .B2(new_n475), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n461), .A2(new_n464), .A3(new_n465), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT93), .ZN(new_n478));
  INV_X1    g292(.A(new_n475), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n477), .A2(new_n478), .A3(new_n479), .A4(new_n390), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n352), .B1(new_n476), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n433), .A2(new_n207), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n296), .A2(G128), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n483), .B1(new_n298), .B2(G128), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT23), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n298), .A2(G128), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n487), .A2(KEYINPUT23), .ZN(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT76), .B(G110), .ZN(new_n489));
  NOR3_X1   g303(.A1(new_n486), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT24), .B(G110), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(KEYINPUT74), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n492), .A2(new_n484), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n405), .B(new_n482), .C1(new_n490), .C2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(G110), .B1(new_n486), .B2(new_n488), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n492), .A2(new_n484), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n495), .A2(new_n496), .A3(new_n408), .A4(new_n406), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n251), .A2(G221), .A3(G234), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n499), .B(KEYINPUT22), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n500), .B(G137), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n494), .A2(new_n497), .A3(new_n501), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n274), .ZN(new_n506));
  INV_X1    g320(.A(G234), .ZN(new_n507));
  OAI21_X1  g321(.A(G217), .B1(new_n507), .B2(G902), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(KEYINPUT73), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT25), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n506), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n503), .A2(new_n504), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n514), .A2(new_n512), .A3(G902), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n511), .B1(new_n517), .B2(new_n510), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n520), .B(G101), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n415), .A2(G210), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n521), .B(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT28), .ZN(new_n525));
  NOR3_X1   g339(.A1(new_n299), .A2(new_n300), .A3(new_n295), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n294), .B1(new_n306), .B2(KEYINPUT67), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT70), .ZN(new_n528));
  NOR3_X1   g342(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(KEYINPUT70), .B1(new_n301), .B2(new_n307), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n247), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n532), .B1(new_n228), .B2(new_n231), .ZN(new_n533));
  OR3_X1    g347(.A1(new_n239), .A2(KEYINPUT65), .A3(G137), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT65), .B1(new_n239), .B2(G137), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n241), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(G131), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n256), .A2(new_n206), .A3(new_n204), .A4(new_n214), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n525), .B1(new_n531), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT71), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI22_X1  g357(.A1(new_n256), .A2(new_n216), .B1(new_n533), .B2(new_n537), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n528), .B1(new_n526), .B2(new_n527), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n301), .A2(KEYINPUT70), .A3(new_n307), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n548), .A2(KEYINPUT71), .A3(new_n525), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n543), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n216), .A2(KEYINPUT69), .A3(new_n256), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT69), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n552), .B1(new_n248), .B2(new_n215), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n554), .A2(new_n538), .A3(new_n547), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n540), .A2(new_n308), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n525), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n524), .B1(new_n550), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT30), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n538), .A2(new_n559), .A3(new_n539), .ZN(new_n560));
  AOI21_X1  g374(.A(KEYINPUT69), .B1(new_n216), .B2(new_n256), .ZN(new_n561));
  NOR3_X1   g375(.A1(new_n248), .A2(new_n215), .A3(new_n552), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n538), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n560), .B1(new_n563), .B2(KEYINPUT30), .ZN(new_n564));
  INV_X1    g378(.A(new_n308), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n555), .B(new_n523), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT31), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n554), .A2(new_n538), .A3(new_n547), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n544), .A2(new_n559), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n551), .A2(new_n553), .B1(new_n537), .B2(new_n533), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n569), .B1(new_n570), .B2(new_n559), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n568), .B1(new_n571), .B2(new_n308), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT31), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n572), .A2(new_n573), .A3(new_n523), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n558), .A2(new_n567), .A3(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(G472), .A2(G902), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n575), .A2(KEYINPUT32), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(KEYINPUT32), .B1(new_n575), .B2(new_n576), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n563), .A2(new_n531), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n525), .B1(new_n580), .B2(new_n555), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n550), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT72), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n582), .A2(new_n583), .A3(KEYINPUT29), .A4(new_n523), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n555), .B1(new_n564), .B2(new_n565), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n524), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n555), .A2(new_n556), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT28), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n588), .A2(new_n543), .A3(new_n549), .A4(new_n523), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT29), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n586), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(KEYINPUT71), .B1(new_n548), .B2(new_n525), .ZN(new_n592));
  AOI211_X1 g406(.A(new_n542), .B(KEYINPUT28), .C1(new_n544), .C2(new_n547), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n547), .B1(new_n554), .B2(new_n538), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT28), .B1(new_n568), .B2(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n594), .A2(KEYINPUT29), .A3(new_n596), .A4(new_n523), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(KEYINPUT72), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n584), .A2(new_n591), .A3(new_n598), .A4(new_n274), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(G472), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n519), .B1(new_n579), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n481), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(G101), .ZN(G3));
  NAND3_X1  g417(.A1(new_n283), .A2(new_n518), .A3(new_n351), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n575), .A2(new_n274), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(G472), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n575), .A2(new_n576), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n348), .A2(new_n479), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n461), .A2(new_n464), .A3(new_n465), .ZN(new_n611));
  INV_X1    g425(.A(new_n383), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT33), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n369), .A2(new_n371), .A3(new_n381), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(KEYINPUT33), .B1(new_n382), .B2(new_n383), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n615), .A2(new_n616), .A3(G478), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n387), .B(new_n274), .C1(new_n382), .C2(new_n383), .ZN(new_n618));
  NAND2_X1  g432(.A1(G478), .A2(G902), .ZN(new_n619));
  AND3_X1   g433(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n611), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n610), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n609), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT34), .B(G104), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G6));
  NAND4_X1  g439(.A1(new_n461), .A2(new_n464), .A3(new_n389), .A4(new_n465), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n610), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n609), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT35), .B(G107), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G9));
  NOR2_X1   g444(.A1(new_n514), .A2(G902), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n631), .A2(KEYINPUT25), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n510), .B1(new_n632), .B2(new_n515), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n498), .A2(KEYINPUT94), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n498), .A2(KEYINPUT94), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n502), .A2(KEYINPUT36), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n637), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n634), .A2(new_n635), .A3(new_n639), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n274), .B(new_n509), .C1(new_n638), .C2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n633), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n606), .A2(new_n607), .A3(new_n642), .ZN(new_n643));
  AOI211_X1 g457(.A(new_n643), .B(new_n352), .C1(new_n476), .C2(new_n480), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT37), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G110), .ZN(G12));
  INV_X1    g460(.A(new_n348), .ZN(new_n647));
  INV_X1    g461(.A(G900), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n470), .B1(new_n474), .B2(new_n648), .ZN(new_n649));
  NOR4_X1   g463(.A1(new_n647), .A2(new_n626), .A3(KEYINPUT95), .A4(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT95), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n626), .A2(new_n649), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n651), .B1(new_n652), .B2(new_n348), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n578), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n575), .A2(KEYINPUT32), .A3(new_n576), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n600), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n283), .A2(new_n351), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n657), .A2(new_n658), .A3(new_n642), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G128), .ZN(G30));
  XOR2_X1   g475(.A(new_n649), .B(KEYINPUT39), .Z(new_n662));
  NAND2_X1  g476(.A1(new_n658), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(new_n663), .B(KEYINPUT40), .Z(new_n664));
  NAND2_X1  g478(.A1(new_n342), .A2(new_n347), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  OR2_X1    g480(.A1(new_n666), .A2(KEYINPUT38), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(KEYINPUT38), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n611), .A2(new_n389), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n572), .A2(new_n524), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n580), .A2(new_n555), .A3(new_n524), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n274), .ZN(new_n675));
  OAI21_X1  g489(.A(G472), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n642), .B1(new_n579), .B2(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n664), .A2(new_n672), .A3(new_n284), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G143), .ZN(G45));
  AND2_X1   g493(.A1(new_n611), .A2(new_n620), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT96), .ZN(new_n681));
  INV_X1    g495(.A(new_n649), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n680), .A2(new_n681), .A3(new_n348), .A4(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n642), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n684), .B1(new_n579), .B2(new_n600), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n348), .A2(new_n611), .A3(new_n620), .A4(new_n682), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(KEYINPUT96), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n683), .A2(new_n685), .A3(new_n658), .A4(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(KEYINPUT97), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT97), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n659), .A2(new_n690), .A3(new_n687), .A4(new_n683), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G146), .ZN(G48));
  OAI21_X1  g507(.A(new_n249), .B1(new_n257), .B2(new_n259), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n279), .B1(new_n694), .B2(new_n261), .ZN(new_n695));
  OAI21_X1  g509(.A(G469), .B1(new_n695), .B2(G902), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n280), .A2(new_n696), .A3(new_n351), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(KEYINPUT98), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT98), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n280), .A2(new_n696), .A3(new_n699), .A4(new_n351), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n698), .A2(KEYINPUT99), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(KEYINPUT99), .B1(new_n698), .B2(new_n700), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n601), .B(new_n622), .C1(new_n701), .C2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT41), .B(G113), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G15));
  OAI211_X1 g519(.A(new_n601), .B(new_n627), .C1(new_n701), .C2(new_n702), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G116), .ZN(G18));
  NAND3_X1  g521(.A1(new_n698), .A2(new_n348), .A3(new_n700), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(KEYINPUT100), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT100), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n698), .A2(new_n710), .A3(new_n348), .A4(new_n700), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n476), .A2(new_n480), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n712), .A2(new_n713), .A3(new_n685), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G119), .ZN(G21));
  OAI211_X1 g529(.A(new_n567), .B(new_n574), .C1(new_n582), .C2(new_n523), .ZN(new_n716));
  XOR2_X1   g530(.A(new_n576), .B(KEYINPUT101), .Z(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n606), .A2(new_n518), .A3(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n671), .ZN(new_n720));
  INV_X1    g534(.A(new_n610), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n720), .B(new_n721), .C1(new_n701), .C2(new_n702), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G122), .ZN(G24));
  NAND3_X1  g537(.A1(new_n611), .A2(new_n620), .A3(new_n682), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n606), .A2(new_n642), .A3(new_n718), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT102), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n606), .A2(new_n642), .A3(KEYINPUT102), .A4(new_n718), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n724), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n712), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G125), .ZN(G27));
  AND2_X1   g545(.A1(new_n260), .A2(new_n269), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(G469), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n280), .A2(new_n282), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(KEYINPUT103), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT103), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n280), .A2(new_n736), .A3(new_n282), .A4(new_n733), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n735), .A2(new_n351), .A3(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(KEYINPUT104), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n665), .A2(new_n285), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT104), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n742), .B1(new_n738), .B2(new_n743), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n740), .A2(new_n744), .A3(new_n601), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n724), .A2(KEYINPUT42), .ZN(new_n746));
  INV_X1    g560(.A(new_n724), .ZN(new_n747));
  AOI22_X1  g561(.A1(new_n655), .A2(KEYINPUT105), .B1(new_n599), .B2(G472), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT105), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n749), .B1(new_n577), .B2(new_n578), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n519), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n740), .A2(new_n744), .A3(new_n747), .A4(new_n751), .ZN(new_n752));
  AOI22_X1  g566(.A1(new_n745), .A2(new_n746), .B1(new_n752), .B2(KEYINPUT42), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G131), .ZN(G33));
  NAND4_X1  g568(.A1(new_n740), .A2(new_n744), .A3(new_n601), .A4(new_n652), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G134), .ZN(G36));
  INV_X1    g570(.A(KEYINPUT108), .ZN(new_n757));
  AOI22_X1  g571(.A1(new_n477), .A2(new_n620), .B1(new_n757), .B2(KEYINPUT43), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n477), .A2(new_n620), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  XOR2_X1   g574(.A(KEYINPUT108), .B(KEYINPUT43), .Z(new_n761));
  AOI21_X1  g575(.A(new_n758), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n762), .A2(KEYINPUT109), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n763), .A2(new_n684), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n762), .A2(KEYINPUT109), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n764), .A2(new_n608), .A3(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT44), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n742), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n270), .A2(new_n271), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT106), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n273), .B1(new_n732), .B2(KEYINPUT45), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n772), .B1(new_n771), .B2(new_n773), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n776), .A2(new_n281), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n777), .A2(KEYINPUT46), .ZN(new_n778));
  OAI211_X1 g592(.A(KEYINPUT46), .B(new_n282), .C1(new_n774), .C2(new_n775), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n280), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT107), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT107), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n779), .A2(new_n782), .A3(new_n280), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n778), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n351), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n764), .A2(KEYINPUT44), .A3(new_n608), .A4(new_n765), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n768), .A2(new_n662), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G137), .ZN(G39));
  INV_X1    g603(.A(KEYINPUT47), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n785), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n784), .A2(KEYINPUT47), .A3(new_n351), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n657), .A2(new_n742), .A3(new_n518), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n793), .A2(new_n747), .A3(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G140), .ZN(G42));
  NAND2_X1  g610(.A1(new_n280), .A2(new_n696), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT110), .ZN(new_n798));
  INV_X1    g612(.A(new_n351), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n791), .A2(new_n792), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n762), .A2(new_n469), .ZN(new_n802));
  INV_X1    g616(.A(new_n719), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(new_n803), .A3(new_n741), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT117), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT51), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n698), .A2(new_n700), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n808), .A2(new_n741), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n579), .A2(new_n676), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n810), .A2(new_n469), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n809), .A2(new_n518), .A3(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n813), .A2(new_n611), .A3(new_n620), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n802), .A2(new_n809), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n815), .B1(new_n727), .B2(new_n728), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n807), .B1(new_n817), .B2(KEYINPUT118), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n669), .A2(new_n284), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n802), .A2(new_n819), .A3(new_n808), .A4(new_n803), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(KEYINPUT50), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT118), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n823), .B1(new_n814), .B2(new_n816), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n806), .A2(new_n818), .A3(new_n822), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n467), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n821), .B1(new_n801), .B2(new_n805), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT51), .B1(new_n827), .B2(new_n817), .ZN(new_n828));
  INV_X1    g642(.A(new_n751), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n815), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(KEYINPUT48), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n802), .A2(new_n803), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n832), .B1(new_n711), .B2(new_n709), .ZN(new_n833));
  NOR4_X1   g647(.A1(new_n826), .A2(new_n828), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n812), .A2(new_n680), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n622), .A2(KEYINPUT111), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT111), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n837), .B1(new_n610), .B2(new_n621), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n836), .A2(new_n609), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n602), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n609), .A2(new_n627), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n644), .A2(new_n842), .A3(KEYINPUT112), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT112), .ZN(new_n844));
  INV_X1    g658(.A(new_n643), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n481), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n844), .B1(new_n846), .B2(new_n628), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n841), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n740), .A2(new_n729), .A3(new_n744), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n466), .A2(new_n649), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n659), .A2(new_n741), .A3(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n755), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n714), .A2(new_n703), .A3(new_n706), .A4(new_n722), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n848), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n854), .A2(new_n753), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT114), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n659), .A2(new_n654), .B1(new_n712), .B2(new_n729), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n671), .A2(new_n647), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n739), .A2(new_n677), .A3(new_n682), .A4(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n692), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(KEYINPUT52), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT52), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n692), .A2(new_n857), .A3(new_n862), .A4(new_n859), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n855), .A2(new_n856), .A3(new_n865), .A4(KEYINPUT53), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n854), .A2(new_n753), .A3(new_n861), .A4(new_n863), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT114), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT113), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n864), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n861), .A2(KEYINPUT113), .A3(new_n863), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT53), .B1(new_n874), .B2(new_n855), .ZN(new_n875));
  OAI21_X1  g689(.A(KEYINPUT54), .B1(new_n870), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n868), .B1(new_n853), .B2(KEYINPUT116), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n706), .A2(new_n722), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT116), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n878), .A2(new_n879), .A3(new_n703), .A4(new_n714), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n877), .A2(new_n753), .A3(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(KEYINPUT115), .B1(new_n848), .B2(new_n852), .ZN(new_n882));
  OAI21_X1  g696(.A(KEYINPUT112), .B1(new_n644), .B2(new_n842), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n846), .A2(new_n844), .A3(new_n628), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n840), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n852), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT115), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n881), .B1(new_n882), .B2(new_n888), .ZN(new_n889));
  AOI22_X1  g703(.A1(new_n874), .A2(new_n889), .B1(new_n868), .B2(new_n867), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT54), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n834), .A2(new_n835), .A3(new_n876), .A4(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n893), .B1(G952), .B2(G953), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n798), .B(KEYINPUT49), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n895), .A2(new_n518), .A3(new_n284), .A4(new_n670), .ZN(new_n896));
  OR4_X1    g710(.A1(new_n799), .A2(new_n896), .A3(new_n810), .A4(new_n759), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n894), .A2(new_n897), .ZN(G75));
  INV_X1    g712(.A(KEYINPUT56), .ZN(new_n899));
  INV_X1    g713(.A(new_n881), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n882), .A2(new_n888), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n861), .A2(KEYINPUT113), .A3(new_n863), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT113), .B1(new_n861), .B2(new_n863), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n900), .B(new_n901), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n867), .A2(new_n868), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(G902), .ZN(new_n907));
  INV_X1    g721(.A(G210), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n899), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OR2_X1    g723(.A1(new_n319), .A2(new_n320), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(new_n291), .Z(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT55), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT119), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n912), .B1(new_n913), .B2(new_n899), .ZN(new_n914));
  OR2_X1    g728(.A1(new_n909), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n251), .A2(G952), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT120), .Z(new_n917));
  NAND2_X1  g731(.A1(new_n909), .A2(new_n914), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n915), .A2(new_n917), .A3(new_n918), .ZN(G51));
  NAND2_X1  g733(.A1(new_n906), .A2(KEYINPUT54), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n892), .A2(new_n920), .A3(KEYINPUT121), .ZN(new_n921));
  OR3_X1    g735(.A1(new_n890), .A2(KEYINPUT121), .A3(new_n891), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n281), .B(KEYINPUT57), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n924), .B1(new_n277), .B2(new_n279), .ZN(new_n925));
  INV_X1    g739(.A(new_n907), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n776), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n916), .B1(new_n925), .B2(new_n927), .ZN(G54));
  NAND3_X1  g742(.A1(new_n926), .A2(KEYINPUT58), .A3(G475), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n929), .A2(new_n459), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n929), .A2(new_n459), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n930), .A2(new_n931), .A3(new_n916), .ZN(G60));
  XOR2_X1   g746(.A(new_n619), .B(KEYINPUT59), .Z(new_n933));
  AOI21_X1  g747(.A(new_n933), .B1(new_n876), .B2(new_n892), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n615), .A2(new_n616), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT122), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n917), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(new_n933), .ZN(new_n938));
  AND4_X1   g752(.A1(new_n922), .A2(new_n921), .A3(new_n938), .A4(new_n936), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n937), .A2(new_n939), .ZN(G63));
  XNOR2_X1  g754(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n370), .A2(new_n274), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n941), .B(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n904), .B2(new_n905), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n917), .B1(new_n945), .B2(new_n505), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n638), .A2(new_n640), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n890), .A2(new_n947), .A3(new_n944), .ZN(new_n948));
  OAI21_X1  g762(.A(KEYINPUT124), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n514), .B1(new_n890), .B2(new_n944), .ZN(new_n950));
  INV_X1    g764(.A(new_n947), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n945), .A2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT124), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n950), .A2(new_n952), .A3(new_n953), .A4(new_n917), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n949), .A2(KEYINPUT61), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(KEYINPUT61), .B1(new_n949), .B2(new_n954), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n955), .A2(new_n956), .ZN(G66));
  INV_X1    g771(.A(G224), .ZN(new_n958));
  OAI21_X1  g772(.A(G953), .B1(new_n472), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n848), .A2(new_n853), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n959), .B1(new_n960), .B2(G953), .ZN(new_n961));
  INV_X1    g775(.A(G898), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n910), .B1(new_n962), .B2(G953), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n961), .B(new_n963), .Z(G69));
  AOI21_X1  g778(.A(new_n251), .B1(G227), .B2(G900), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n795), .A2(new_n755), .A3(new_n788), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT126), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n786), .A2(new_n662), .A3(new_n858), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n692), .B(new_n857), .C1(new_n968), .C2(new_n829), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n966), .A2(new_n967), .A3(new_n970), .A4(new_n753), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n795), .A2(new_n753), .A3(new_n755), .A4(new_n788), .ZN(new_n972));
  OAI21_X1  g786(.A(KEYINPUT126), .B1(new_n972), .B2(new_n969), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n971), .A2(new_n251), .A3(new_n973), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n571), .B(new_n440), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n975), .B1(G900), .B2(G953), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n795), .A2(new_n788), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n621), .A2(new_n626), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n601), .A2(new_n979), .ZN(new_n980));
  NOR3_X1   g794(.A1(new_n980), .A2(new_n663), .A3(new_n742), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n678), .A2(new_n692), .A3(new_n857), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT62), .ZN(new_n983));
  OR2_X1    g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n982), .A2(new_n983), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n981), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n978), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n251), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n988), .A2(KEYINPUT125), .A3(new_n975), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT125), .ZN(new_n990));
  AOI21_X1  g804(.A(G953), .B1(new_n978), .B2(new_n986), .ZN(new_n991));
  INV_X1    g805(.A(new_n975), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n989), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n965), .B1(new_n977), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n974), .A2(new_n976), .ZN(new_n996));
  INV_X1    g810(.A(new_n965), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n996), .A2(new_n997), .A3(new_n993), .A4(new_n989), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n995), .A2(new_n998), .ZN(G72));
  XNOR2_X1  g813(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1000));
  NAND2_X1  g814(.A1(G472), .A2(G902), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(new_n960), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n1002), .B1(new_n987), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n916), .B1(new_n1004), .B2(new_n673), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n586), .A2(new_n566), .ZN(new_n1006));
  OAI211_X1 g820(.A(new_n1002), .B(new_n1006), .C1(new_n870), .C2(new_n875), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n971), .A2(new_n960), .A3(new_n973), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n523), .B1(new_n1009), .B2(new_n1002), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1008), .B1(new_n572), .B2(new_n1010), .ZN(G57));
endmodule


