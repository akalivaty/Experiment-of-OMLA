//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 0 0 1 1 1 1 1 1 1 1 1 0 1 1 0 0 0 1 0 0 1 1 0 0 0 0 1 0 1 1 1 0 0 0 1 1 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n565, new_n566,
    new_n567, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n618,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1205, new_n1206, new_n1207, new_n1208;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT65), .Z(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n466));
  AND3_X1   g041(.A1(new_n463), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n466), .B1(new_n463), .B2(new_n465), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  INV_X1    g045(.A(G113), .ZN(new_n471));
  OAI22_X1  g046(.A1(new_n469), .A2(new_n470), .B1(new_n471), .B2(new_n464), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT67), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n473), .B1(new_n462), .B2(G2104), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n464), .A2(KEYINPUT67), .A3(KEYINPUT3), .ZN(new_n475));
  INV_X1    g050(.A(G137), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NAND4_X1  g052(.A1(new_n474), .A2(new_n475), .A3(new_n477), .A4(new_n463), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n464), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G101), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT68), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n478), .A2(KEYINPUT68), .A3(new_n480), .ZN(new_n484));
  AOI22_X1  g059(.A1(new_n472), .A2(G2105), .B1(new_n483), .B2(new_n484), .ZN(G160));
  NAND3_X1  g060(.A1(new_n474), .A2(new_n463), .A3(new_n475), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n486), .B(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G136), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n488), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G124), .ZN(new_n495));
  OR2_X1    g070(.A1(G100), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G112), .C2(new_n489), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n492), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G162));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  NOR3_X1   g075(.A1(new_n500), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n501), .B1(new_n467), .B2(new_n468), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n500), .A2(G2105), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n474), .A2(new_n475), .A3(new_n503), .A4(new_n463), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  AND2_X1   g081(.A1(new_n475), .A2(new_n463), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n508));
  AND2_X1   g083(.A1(G126), .A2(G2105), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n507), .A2(new_n508), .A3(new_n474), .A4(new_n509), .ZN(new_n510));
  NAND4_X1  g085(.A1(new_n474), .A2(new_n475), .A3(new_n463), .A4(new_n509), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT70), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g088(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n514));
  INV_X1    g089(.A(G114), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n514), .B1(new_n515), .B2(G2105), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n506), .A2(new_n513), .A3(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(G164));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(G75), .A2(G543), .ZN(new_n521));
  XOR2_X1   g096(.A(new_n521), .B(KEYINPUT71), .Z(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT5), .B(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G62), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n520), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G543), .ZN(new_n526));
  OR2_X1    g101(.A1(KEYINPUT6), .A2(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G50), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n527), .A2(new_n528), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(new_n523), .ZN(new_n532));
  INV_X1    g107(.A(G88), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n525), .A2(new_n534), .ZN(G303));
  INV_X1    g110(.A(G303), .ZN(G166));
  XNOR2_X1  g111(.A(KEYINPUT72), .B(KEYINPUT7), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n537), .B(new_n538), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n531), .A2(new_n523), .ZN(new_n540));
  XNOR2_X1  g115(.A(KEYINPUT73), .B(G89), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(KEYINPUT74), .ZN(new_n543));
  AND2_X1   g118(.A1(G63), .A2(G651), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n529), .A2(G51), .B1(new_n523), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n542), .A2(KEYINPUT74), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n546), .A2(new_n547), .ZN(G168));
  NAND2_X1  g123(.A1(new_n529), .A2(G52), .ZN(new_n549));
  INV_X1    g124(.A(G90), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n532), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(new_n520), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n551), .A2(new_n553), .ZN(G301));
  INV_X1    g129(.A(G301), .ZN(G171));
  NAND2_X1  g130(.A1(new_n529), .A2(G43), .ZN(new_n556));
  INV_X1    g131(.A(G81), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n532), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n523), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n559), .A2(new_n520), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT75), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g139(.A(KEYINPUT76), .B(KEYINPUT8), .Z(new_n565));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n565), .B(new_n566), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  AOI22_X1  g143(.A1(new_n523), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n569));
  INV_X1    g144(.A(G91), .ZN(new_n570));
  OAI22_X1  g145(.A1(new_n569), .A2(new_n520), .B1(new_n532), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT9), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n573), .B1(new_n529), .B2(G53), .ZN(new_n574));
  AND2_X1   g149(.A1(KEYINPUT6), .A2(G651), .ZN(new_n575));
  NOR2_X1   g150(.A1(KEYINPUT6), .A2(G651), .ZN(new_n576));
  OAI211_X1 g151(.A(G53), .B(G543), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n577), .A2(KEYINPUT9), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n572), .B1(new_n574), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n529), .A2(new_n573), .A3(G53), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n577), .A2(KEYINPUT9), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n580), .A2(new_n581), .A3(KEYINPUT77), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n571), .B1(new_n579), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G299));
  INV_X1    g159(.A(G168), .ZN(G286));
  OR2_X1    g160(.A1(new_n523), .A2(G74), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n586), .A2(G651), .B1(G49), .B2(new_n529), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT78), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n588), .B1(new_n540), .B2(G87), .ZN(new_n589));
  INV_X1    g164(.A(G87), .ZN(new_n590));
  NOR3_X1   g165(.A1(new_n532), .A2(KEYINPUT78), .A3(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n587), .B1(new_n589), .B2(new_n591), .ZN(G288));
  AOI22_X1  g167(.A1(new_n540), .A2(G86), .B1(G48), .B2(new_n529), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n523), .A2(G61), .ZN(new_n594));
  NAND2_X1  g169(.A1(G73), .A2(G543), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n520), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n593), .A2(new_n597), .ZN(G305));
  XNOR2_X1  g173(.A(KEYINPUT79), .B(G47), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n540), .A2(G85), .B1(new_n529), .B2(new_n599), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT80), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n520), .B2(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n540), .A2(G92), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT10), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n606), .B1(G54), .B2(new_n529), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n523), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n520), .B1(new_n608), .B2(KEYINPUT81), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(KEYINPUT81), .B2(new_n608), .ZN(new_n610));
  AND2_X1   g185(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n604), .B1(new_n611), .B2(G868), .ZN(G284));
  OAI21_X1  g187(.A(new_n604), .B1(new_n611), .B2(G868), .ZN(G321));
  INV_X1    g188(.A(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(G299), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G168), .B2(new_n614), .ZN(G297));
  OAI21_X1  g191(.A(new_n615), .B1(G168), .B2(new_n614), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n611), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND2_X1  g194(.A1(new_n611), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G868), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(G868), .B2(new_n561), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n463), .A2(new_n465), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(KEYINPUT66), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n463), .A2(new_n465), .A3(new_n466), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(new_n479), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2100), .ZN(new_n631));
  OR2_X1    g206(.A1(G99), .A2(G2105), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n632), .B(G2104), .C1(G111), .C2(new_n489), .ZN(new_n633));
  INV_X1    g208(.A(G135), .ZN(new_n634));
  INV_X1    g209(.A(G123), .ZN(new_n635));
  OAI221_X1 g210(.A(new_n633), .B1(new_n490), .B2(new_n634), .C1(new_n635), .C2(new_n493), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n636), .A2(G2096), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(G2096), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n631), .A2(new_n637), .A3(new_n638), .ZN(G156));
  XOR2_X1   g214(.A(KEYINPUT15), .B(G2435), .Z(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT83), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2427), .B(G2430), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT82), .B(KEYINPUT14), .Z(new_n646));
  NAND2_X1  g221(.A1(new_n642), .A2(new_n644), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n648), .B(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(G14), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n656), .B2(new_n654), .ZN(G401));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  XOR2_X1   g234(.A(G2072), .B(G2078), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT84), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT85), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n659), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n663), .B1(new_n662), .B2(new_n661), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2084), .B(G2090), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n661), .B(KEYINPUT17), .Z(new_n666));
  INV_X1    g241(.A(new_n659), .ZN(new_n667));
  OAI211_X1 g242(.A(new_n664), .B(new_n665), .C1(new_n666), .C2(new_n667), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(new_n665), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n661), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT18), .Z(new_n671));
  NOR2_X1   g246(.A1(new_n659), .A2(new_n665), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n668), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2096), .B(G2100), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(G227));
  XOR2_X1   g252(.A(G1971), .B(G1976), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  XOR2_X1   g255(.A(G1961), .B(G1966), .Z(new_n681));
  AND2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT20), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n680), .A2(new_n681), .ZN(new_n685));
  NOR3_X1   g260(.A1(new_n679), .A2(new_n682), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(new_n679), .B2(new_n685), .ZN(new_n687));
  AND2_X1   g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G1991), .B(G1996), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1981), .B(G1986), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(G229));
  NAND2_X1  g270(.A1(new_n491), .A2(G141), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n494), .A2(G129), .ZN(new_n697));
  NAND3_X1  g272(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT26), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  AOI22_X1  g276(.A1(new_n700), .A2(new_n701), .B1(G105), .B2(new_n479), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n696), .A2(new_n697), .A3(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G29), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n705), .A2(KEYINPUT94), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n705), .B(KEYINPUT94), .C1(G29), .C2(G32), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT27), .B(G1996), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(G164), .A2(G29), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G27), .B2(G29), .ZN(new_n713));
  INV_X1    g288(.A(G2078), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n491), .A2(G139), .ZN(new_n716));
  AOI22_X1  g291(.A1(new_n627), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n717), .A2(new_n489), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n489), .A2(G103), .A3(G2104), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT25), .Z(new_n720));
  NAND3_X1  g295(.A1(new_n716), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G29), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n723), .B2(G33), .ZN(new_n725));
  INV_X1    g300(.A(G2072), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n715), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(G160), .A2(G29), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT93), .B(KEYINPUT24), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(G34), .Z(new_n730));
  OAI21_X1  g305(.A(new_n728), .B1(G29), .B2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G2084), .ZN(new_n732));
  OAI22_X1  g307(.A1(new_n713), .A2(new_n714), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NOR3_X1   g308(.A1(new_n711), .A2(new_n727), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n725), .A2(KEYINPUT92), .A3(new_n726), .ZN(new_n735));
  AOI21_X1  g310(.A(KEYINPUT92), .B1(new_n725), .B2(new_n726), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n636), .A2(new_n723), .ZN(new_n737));
  INV_X1    g312(.A(G16), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G21), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G168), .B2(new_n738), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n737), .B1(new_n740), .B2(G1966), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT31), .B(G11), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT30), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n743), .A2(G28), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n723), .B1(new_n743), .B2(G28), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n738), .A2(G5), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G301), .B2(G16), .ZN(new_n747));
  INV_X1    g322(.A(G1961), .ZN(new_n748));
  OAI221_X1 g323(.A(new_n742), .B1(new_n744), .B2(new_n745), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n741), .B(new_n750), .C1(G1966), .C2(new_n740), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n736), .A2(new_n751), .ZN(new_n752));
  AND3_X1   g327(.A1(new_n734), .A2(new_n735), .A3(new_n752), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n708), .A2(new_n710), .B1(new_n748), .B2(new_n747), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n731), .A2(new_n732), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT95), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(KEYINPUT96), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n757), .A2(KEYINPUT96), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n753), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n760), .A2(KEYINPUT97), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT97), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n753), .A2(new_n759), .A3(new_n762), .A4(new_n758), .ZN(new_n763));
  NOR2_X1   g338(.A1(G29), .A2(G35), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G162), .B2(G29), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT98), .B(KEYINPUT29), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(G2090), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n738), .A2(G20), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT23), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n583), .B2(new_n738), .ZN(new_n772));
  INV_X1    g347(.A(G1956), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(G4), .A2(G16), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n611), .B2(G16), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n776), .A2(G1348), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n776), .A2(G1348), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n738), .A2(G19), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n561), .B2(new_n738), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1341), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n769), .A2(new_n774), .A3(new_n777), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n723), .A2(G26), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT28), .Z(new_n785));
  OR2_X1    g360(.A1(G104), .A2(G2105), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n786), .B(G2104), .C1(G116), .C2(new_n489), .ZN(new_n787));
  INV_X1    g362(.A(G140), .ZN(new_n788));
  INV_X1    g363(.A(G128), .ZN(new_n789));
  OAI221_X1 g364(.A(new_n787), .B1(new_n490), .B2(new_n788), .C1(new_n789), .C2(new_n493), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT91), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n785), .B1(new_n791), .B2(G29), .ZN(new_n792));
  INV_X1    g367(.A(G2067), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n767), .A2(new_n768), .ZN(new_n795));
  NOR3_X1   g370(.A1(new_n783), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n761), .A2(new_n763), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n738), .A2(G22), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G166), .B2(new_n738), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT88), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n800), .A2(G1971), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(G1971), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n738), .A2(G23), .ZN(new_n803));
  INV_X1    g378(.A(G288), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(new_n738), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT33), .B(G1976), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  MUX2_X1   g382(.A(G6), .B(G305), .S(G16), .Z(new_n808));
  XOR2_X1   g383(.A(KEYINPUT32), .B(G1981), .Z(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT87), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n808), .B(new_n810), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n801), .A2(new_n802), .A3(new_n807), .A4(new_n811), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n812), .A2(KEYINPUT34), .ZN(new_n813));
  OR2_X1    g388(.A1(G25), .A2(G29), .ZN(new_n814));
  OAI21_X1  g389(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n815));
  INV_X1    g390(.A(G107), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n815), .B1(new_n816), .B2(G2105), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(new_n491), .B2(G131), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT86), .ZN(new_n819));
  AND3_X1   g394(.A1(new_n494), .A2(new_n819), .A3(G119), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n819), .B1(new_n494), .B2(G119), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n818), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n814), .B1(new_n822), .B2(new_n723), .ZN(new_n823));
  XOR2_X1   g398(.A(KEYINPUT35), .B(G1991), .Z(new_n824));
  AOI22_X1  g399(.A1(new_n812), .A2(KEYINPUT34), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  MUX2_X1   g400(.A(G24), .B(G290), .S(G16), .Z(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(G1986), .Z(new_n827));
  OR2_X1    g402(.A1(new_n823), .A2(new_n824), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n813), .A2(new_n825), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n829), .A2(KEYINPUT36), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT90), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n829), .A2(KEYINPUT36), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT89), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n797), .B1(new_n832), .B2(new_n834), .ZN(G311));
  NAND2_X1  g410(.A1(new_n832), .A2(new_n834), .ZN(new_n836));
  AND3_X1   g411(.A1(new_n761), .A2(new_n763), .A3(new_n796), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(G150));
  NAND2_X1  g413(.A1(new_n611), .A2(G559), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT38), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n529), .A2(G55), .ZN(new_n841));
  INV_X1    g416(.A(G93), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n841), .B1(new_n532), .B2(new_n842), .ZN(new_n843));
  AOI22_X1  g418(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n844), .A2(new_n520), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n561), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n561), .A2(new_n846), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n840), .B(new_n850), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n851), .A2(KEYINPUT39), .ZN(new_n852));
  INV_X1    g427(.A(G860), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(KEYINPUT39), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n846), .A2(new_n853), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT37), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(G145));
  XNOR2_X1  g433(.A(new_n498), .B(G160), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(new_n636), .Z(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT99), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n791), .A2(new_n703), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n790), .A2(KEYINPUT91), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n790), .A2(KEYINPUT91), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n864), .A2(new_n704), .A3(new_n865), .ZN(new_n866));
  AND3_X1   g441(.A1(new_n863), .A2(G164), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(G164), .B1(new_n863), .B2(new_n866), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n862), .B(new_n722), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n863), .A2(new_n866), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(new_n518), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n722), .A2(new_n862), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n721), .A2(KEYINPUT99), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n863), .A2(G164), .A3(new_n866), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n871), .A2(new_n872), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n822), .B(new_n629), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n491), .A2(G142), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n494), .A2(G130), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n489), .A2(G118), .ZN(new_n879));
  OAI21_X1  g454(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n877), .B(new_n878), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n876), .B(new_n881), .Z(new_n882));
  AND3_X1   g457(.A1(new_n869), .A2(new_n875), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n882), .B1(new_n869), .B2(new_n875), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n861), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n869), .A2(new_n875), .ZN(new_n886));
  INV_X1    g461(.A(new_n882), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n869), .A2(new_n875), .A3(new_n882), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n888), .A2(new_n860), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(G37), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n885), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  XOR2_X1   g467(.A(KEYINPUT100), .B(KEYINPUT40), .Z(new_n893));
  XNOR2_X1  g468(.A(new_n892), .B(new_n893), .ZN(G395));
  XOR2_X1   g469(.A(G288), .B(KEYINPUT101), .Z(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(G305), .ZN(new_n896));
  XNOR2_X1  g471(.A(G290), .B(G166), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n896), .B(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n899));
  NOR3_X1   g474(.A1(new_n898), .A2(KEYINPUT102), .A3(new_n899), .ZN(new_n900));
  XOR2_X1   g475(.A(new_n896), .B(new_n897), .Z(new_n901));
  NOR2_X1   g476(.A1(new_n899), .A2(KEYINPUT102), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n899), .A2(KEYINPUT102), .ZN(new_n903));
  NOR3_X1   g478(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n607), .A2(new_n610), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(G299), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n905), .A2(G299), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT41), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n910), .B1(new_n907), .B2(new_n908), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n611), .A2(new_n583), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n912), .A2(KEYINPUT41), .A3(new_n906), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n620), .B(new_n850), .ZN(new_n916));
  MUX2_X1   g491(.A(new_n909), .B(new_n915), .S(new_n916), .Z(new_n917));
  AOI211_X1 g492(.A(new_n900), .B(new_n904), .C1(new_n917), .C2(KEYINPUT103), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n917), .A2(KEYINPUT103), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR4_X1   g495(.A1(new_n917), .A2(new_n904), .A3(KEYINPUT103), .A4(new_n900), .ZN(new_n921));
  OAI21_X1  g496(.A(G868), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n614), .B1(new_n843), .B2(new_n845), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(G295));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n923), .ZN(G331));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n926));
  XNOR2_X1  g501(.A(G301), .B(KEYINPUT104), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(new_n849), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n927), .A2(new_n849), .ZN(new_n930));
  OAI21_X1  g505(.A(G286), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n930), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n932), .A2(new_n928), .A3(G168), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n909), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n933), .A2(new_n931), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n934), .B1(new_n914), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n901), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n898), .B(new_n934), .C1(new_n914), .C2(new_n935), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n937), .A2(new_n938), .A3(new_n891), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT105), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n926), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT43), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n937), .A2(new_n938), .A3(new_n943), .A4(new_n891), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n940), .A2(new_n944), .ZN(new_n945));
  XOR2_X1   g520(.A(new_n942), .B(new_n945), .Z(G397));
  NAND2_X1  g521(.A1(new_n791), .A2(G2067), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n864), .A2(new_n793), .A3(new_n865), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n947), .A2(new_n704), .A3(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(G1384), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n518), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT45), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n470), .B1(new_n625), .B2(new_n626), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n471), .A2(new_n464), .ZN(new_n955));
  OAI21_X1  g530(.A(G2105), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n483), .A2(new_n484), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n956), .A2(new_n957), .A3(G40), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n953), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n949), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G1996), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n962), .B(KEYINPUT46), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT125), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT125), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n960), .A2(new_n966), .A3(new_n963), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT47), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n965), .A2(KEYINPUT47), .A3(new_n967), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n703), .B(new_n961), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n947), .A2(new_n948), .A3(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n824), .ZN(new_n974));
  OR2_X1    g549(.A1(new_n822), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n948), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n822), .B(new_n974), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n959), .B1(new_n973), .B2(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(G290), .A2(G1986), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(new_n959), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n980), .B(KEYINPUT48), .ZN(new_n981));
  AOI22_X1  g556(.A1(new_n959), .A2(new_n976), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n970), .A2(new_n971), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT126), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT126), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n970), .A2(new_n982), .A3(new_n985), .A4(new_n971), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT50), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(new_n518), .B2(new_n950), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n516), .B1(new_n510), .B2(new_n512), .ZN(new_n991));
  AOI21_X1  g566(.A(G1384), .B1(new_n991), .B2(new_n506), .ZN(new_n992));
  XNOR2_X1  g567(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n993));
  AOI22_X1  g568(.A1(new_n989), .A2(new_n990), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n956), .A2(new_n957), .A3(G40), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT109), .B1(new_n992), .B2(new_n988), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n994), .A2(new_n732), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1966), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n995), .B1(KEYINPUT45), .B2(new_n992), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n952), .A2(G1384), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n511), .A2(KEYINPUT70), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n511), .A2(KEYINPUT70), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n517), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n627), .A2(new_n501), .B1(KEYINPUT4), .B2(new_n504), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1000), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n998), .B1(new_n999), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n997), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(G8), .ZN(new_n1009));
  INV_X1    g584(.A(G8), .ZN(new_n1010));
  NOR2_X1   g585(.A1(G168), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1009), .A2(KEYINPUT51), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT51), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1014), .B(G8), .C1(new_n1008), .C2(G286), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT120), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n1008), .A2(KEYINPUT120), .A3(new_n1011), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1013), .B(new_n1015), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT62), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT107), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1005), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n518), .A2(KEYINPUT107), .A3(new_n1000), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n958), .B1(new_n951), .B2(new_n952), .ZN(new_n1024));
  AOI21_X1  g599(.A(G1971), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OAI211_X1 g600(.A(G160), .B(G40), .C1(new_n992), .C2(new_n993), .ZN(new_n1026));
  AOI211_X1 g601(.A(KEYINPUT50), .B(G1384), .C1(new_n991), .C2(new_n506), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n1026), .A2(G2090), .A3(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(G8), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(G303), .A2(G8), .ZN(new_n1030));
  XNOR2_X1  g605(.A(KEYINPUT110), .B(KEYINPUT55), .ZN(new_n1031));
  XNOR2_X1  g606(.A(new_n1030), .B(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1032), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n951), .A2(new_n990), .A3(KEYINPUT50), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n992), .A2(new_n993), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n958), .A2(G2090), .ZN(new_n1037));
  AND4_X1   g612(.A1(new_n996), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1034), .B(G8), .C1(new_n1038), .C2(new_n1025), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n587), .B(G1976), .C1(new_n589), .C2(new_n591), .ZN(new_n1040));
  OAI211_X1 g615(.A(G8), .B(new_n1040), .C1(new_n951), .C2(new_n958), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT52), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n995), .A2(new_n992), .ZN(new_n1043));
  INV_X1    g618(.A(G1981), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n593), .A2(new_n597), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n529), .A2(G48), .ZN(new_n1046));
  INV_X1    g621(.A(G86), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1046), .B1(new_n532), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(G1981), .B1(new_n1048), .B2(new_n596), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT112), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1045), .B(new_n1049), .C1(new_n1050), .C2(KEYINPUT49), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1050), .A2(KEYINPUT49), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1044), .B1(new_n593), .B2(new_n597), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n1048), .A2(new_n596), .A3(G1981), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1052), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1043), .A2(G8), .A3(new_n1051), .A4(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1042), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT111), .ZN(new_n1058));
  INV_X1    g633(.A(G1976), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT52), .B1(G288), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1058), .B1(new_n1041), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1010), .B1(new_n995), .B2(new_n992), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1063), .A2(KEYINPUT111), .A3(new_n1040), .A4(new_n1060), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1057), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1033), .A2(new_n1039), .A3(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1024), .A2(new_n714), .A3(new_n1005), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT122), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1024), .A2(KEYINPUT122), .A3(new_n714), .A4(new_n1005), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(KEYINPUT53), .A3(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1023), .A2(new_n714), .A3(new_n1024), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1035), .A2(new_n996), .A3(new_n995), .A4(new_n1036), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1072), .A2(new_n1073), .B1(new_n1074), .B2(new_n748), .ZN(new_n1075));
  AOI21_X1  g650(.A(G301), .B1(new_n1071), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1019), .A2(new_n1066), .A3(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1018), .A2(KEYINPUT62), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(G8), .B1(new_n1038), .B2(new_n1025), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1034), .B1(new_n1080), .B2(KEYINPUT116), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(KEYINPUT116), .B2(new_n1080), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1057), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT113), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1083), .A2(new_n1084), .A3(KEYINPUT113), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AOI211_X1 g664(.A(new_n1010), .B(G286), .C1(new_n997), .C2(new_n1007), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1039), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT63), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1082), .A2(new_n1089), .A3(new_n1090), .A4(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1090), .A2(new_n1033), .A3(new_n1039), .A4(new_n1065), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1095), .A2(KEYINPUT115), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1092), .B1(new_n1095), .B2(KEYINPUT115), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1094), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT114), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1039), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1056), .A2(new_n1059), .A3(new_n804), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n1045), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n1063), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1099), .B1(new_n1100), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1088), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT113), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1091), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1108), .A2(KEYINPUT114), .A3(new_n1103), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1105), .A2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT56), .B(G2072), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1023), .A2(new_n1024), .A3(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n773), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n571), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT57), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n580), .A2(new_n581), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1115), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1118), .B1(new_n583), .B2(new_n1116), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(KEYINPUT117), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT117), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1118), .B(new_n1121), .C1(new_n583), .C2(new_n1116), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1114), .A2(new_n1124), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n951), .A2(new_n958), .A3(G2067), .ZN(new_n1126));
  INV_X1    g701(.A(G1348), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1126), .B1(new_n1074), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1125), .B1(new_n905), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1112), .A2(new_n1123), .A3(new_n1113), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT118), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT118), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1112), .A2(new_n1123), .A3(new_n1113), .A4(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1129), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1125), .A2(KEYINPUT61), .A3(new_n1130), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT60), .ZN(new_n1138));
  AOI211_X1 g713(.A(new_n1138), .B(new_n1126), .C1(new_n1074), .C2(new_n1127), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(new_n905), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT59), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1023), .A2(new_n961), .A3(new_n1024), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT119), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1023), .A2(KEYINPUT119), .A3(new_n1024), .A4(new_n961), .ZN(new_n1146));
  XOR2_X1   g721(.A(KEYINPUT58), .B(G1341), .Z(new_n1147));
  NAND2_X1  g722(.A1(new_n1043), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1145), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1142), .B1(new_n1149), .B2(new_n561), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1149), .A2(new_n1142), .A3(new_n561), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1141), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1128), .A2(KEYINPUT60), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n1154), .A2(new_n1139), .A3(new_n905), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1134), .A2(new_n1125), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1155), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1136), .B1(new_n1153), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1074), .A2(new_n748), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1023), .A2(KEYINPUT53), .A3(new_n1024), .A4(new_n714), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(KEYINPUT123), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT123), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1075), .A2(new_n1165), .A3(new_n1162), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1164), .A2(G171), .A3(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1071), .A2(G301), .A3(new_n1075), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1167), .A2(KEYINPUT54), .A3(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g744(.A(KEYINPUT121), .B(KEYINPUT54), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1163), .A2(G171), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1170), .B1(new_n1171), .B2(new_n1076), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1169), .A2(new_n1018), .A3(new_n1066), .A4(new_n1172), .ZN(new_n1173));
  OAI211_X1 g748(.A(new_n1098), .B(new_n1110), .C1(new_n1159), .C2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT124), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT115), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1066), .A2(new_n1177), .A3(new_n1090), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1095), .A2(KEYINPUT115), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1178), .A2(new_n1092), .A3(new_n1179), .ZN(new_n1180));
  AOI22_X1  g755(.A1(new_n1180), .A2(new_n1094), .B1(new_n1105), .B2(new_n1109), .ZN(new_n1181));
  AND3_X1   g756(.A1(new_n1149), .A2(new_n1142), .A3(new_n561), .ZN(new_n1182));
  OAI211_X1 g757(.A(new_n1137), .B(new_n1140), .C1(new_n1182), .C2(new_n1150), .ZN(new_n1183));
  AOI22_X1  g758(.A1(new_n1131), .A2(new_n1133), .B1(new_n1124), .B2(new_n1114), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1128), .A2(KEYINPUT60), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1185), .A2(new_n611), .ZN(new_n1186));
  OAI22_X1  g761(.A1(new_n1184), .A2(KEYINPUT61), .B1(new_n1154), .B2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1135), .B1(new_n1183), .B2(new_n1187), .ZN(new_n1188));
  AND3_X1   g763(.A1(new_n1018), .A2(new_n1066), .A3(new_n1172), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1188), .A2(new_n1189), .A3(new_n1169), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1181), .A2(new_n1190), .A3(KEYINPUT124), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1079), .B1(new_n1176), .B2(new_n1191), .ZN(new_n1192));
  AND2_X1   g767(.A1(G290), .A2(G1986), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n959), .B1(new_n1193), .B2(new_n979), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n978), .A2(new_n1194), .ZN(new_n1195));
  XOR2_X1   g770(.A(new_n1195), .B(KEYINPUT106), .Z(new_n1196));
  OAI21_X1  g771(.A(new_n987), .B1(new_n1192), .B2(new_n1196), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g772(.A1(G401), .A2(G227), .A3(new_n460), .ZN(new_n1199));
  NAND2_X1  g773(.A1(new_n694), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g774(.A(new_n1200), .B1(new_n940), .B2(new_n944), .ZN(new_n1201));
  AND3_X1   g775(.A1(new_n892), .A2(KEYINPUT127), .A3(new_n1201), .ZN(new_n1202));
  AOI21_X1  g776(.A(KEYINPUT127), .B1(new_n892), .B2(new_n1201), .ZN(new_n1203));
  NOR2_X1   g777(.A1(new_n1202), .A2(new_n1203), .ZN(G308));
  NAND2_X1  g778(.A1(new_n892), .A2(new_n1201), .ZN(new_n1205));
  INV_X1    g779(.A(KEYINPUT127), .ZN(new_n1206));
  NAND2_X1  g780(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g781(.A1(new_n892), .A2(KEYINPUT127), .A3(new_n1201), .ZN(new_n1208));
  NAND2_X1  g782(.A1(new_n1207), .A2(new_n1208), .ZN(G225));
endmodule


