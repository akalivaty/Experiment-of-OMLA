//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 1 1 0 1 0 1 0 0 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 1 0 1 1 0 0 1 0 1 0 0 0 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1246, new_n1247, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT0), .Z(new_n206));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n207));
  INV_X1    g0007(.A(G87), .ZN(new_n208));
  INV_X1    g0008(.A(G250), .ZN(new_n209));
  INV_X1    g0009(.A(G97), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(KEYINPUT64), .ZN(new_n213));
  OR2_X1    g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(new_n212), .A2(new_n213), .B1(G77), .B2(G244), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G116), .A2(G270), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G68), .A2(G238), .ZN(new_n217));
  NAND4_X1  g0017(.A1(new_n214), .A2(new_n215), .A3(new_n216), .A4(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G50), .ZN(new_n219));
  INV_X1    g0019(.A(G226), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n203), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n222), .B(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(G58), .A2(G68), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G50), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n206), .B(new_n224), .C1(new_n227), .C2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(KEYINPUT66), .B(G250), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT67), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XOR2_X1   g0043(.A(G50), .B(G58), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G351));
  OAI21_X1  g0049(.A(G20), .B1(new_n229), .B2(G50), .ZN(new_n250));
  INV_X1    g0050(.A(G150), .ZN(new_n251));
  NOR2_X1   g0051(.A1(G20), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT8), .ZN(new_n254));
  INV_X1    g0054(.A(G58), .ZN(new_n255));
  OR3_X1    g0055(.A1(new_n254), .A2(new_n255), .A3(KEYINPUT69), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n254), .B1(new_n255), .B2(KEYINPUT69), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(G20), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  OAI221_X1 g0061(.A(new_n250), .B1(new_n251), .B2(new_n253), .C1(new_n258), .C2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n225), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G13), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(new_n226), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n262), .A2(new_n264), .B1(new_n219), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n265), .A2(G20), .ZN(new_n269));
  XNOR2_X1  g0069(.A(new_n269), .B(KEYINPUT71), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G50), .ZN(new_n271));
  XOR2_X1   g0071(.A(new_n271), .B(KEYINPUT72), .Z(new_n272));
  INV_X1    g0072(.A(new_n264), .ZN(new_n273));
  INV_X1    g0073(.A(G13), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(G1), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G20), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT70), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n273), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(KEYINPUT70), .B1(new_n267), .B2(new_n264), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n268), .B1(new_n272), .B2(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(new_n281), .B(KEYINPUT9), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT3), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n287), .A2(G222), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT68), .ZN(new_n290));
  OR2_X1    g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n286), .A2(G77), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n287), .A2(G223), .A3(G1698), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n289), .A2(new_n290), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n291), .A2(new_n292), .A3(new_n293), .A4(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n225), .B1(G33), .B2(G41), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n265), .B1(G41), .B2(G45), .ZN(new_n298));
  INV_X1    g0098(.A(G274), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n296), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n302), .A2(new_n298), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G226), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n297), .A2(new_n301), .A3(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G190), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n282), .A2(KEYINPUT75), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT10), .ZN(new_n310));
  INV_X1    g0110(.A(G200), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n309), .A2(new_n310), .A3(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(KEYINPUT10), .B1(new_n308), .B2(new_n312), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G179), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n306), .A2(new_n317), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n318), .B(new_n281), .C1(G169), .C2(new_n306), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n278), .A2(new_n279), .A3(new_n270), .ZN(new_n321));
  INV_X1    g0121(.A(new_n258), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n258), .A2(new_n276), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT79), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT79), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n323), .A2(new_n327), .A3(new_n324), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n284), .A2(G33), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT77), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(new_n259), .B2(KEYINPUT3), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n284), .A2(KEYINPUT77), .A3(G33), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n330), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n220), .A2(G1698), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(G223), .A2(G1698), .ZN(new_n337));
  OAI22_X1  g0137(.A1(new_n336), .A2(new_n337), .B1(new_n259), .B2(new_n208), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n296), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n303), .A2(G232), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n339), .A2(new_n301), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(G200), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT16), .ZN(new_n343));
  INV_X1    g0143(.A(G68), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT7), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(new_n287), .B2(G20), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n286), .A2(KEYINPUT7), .A3(new_n226), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n344), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n255), .A2(new_n344), .ZN(new_n349));
  OAI21_X1  g0149(.A(G20), .B1(new_n349), .B2(new_n228), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT78), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n252), .A2(G159), .ZN(new_n353));
  OAI211_X1 g0153(.A(KEYINPUT78), .B(G20), .C1(new_n349), .C2(new_n228), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n343), .B1(new_n348), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n332), .A2(new_n333), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n283), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n358), .A2(new_n345), .A3(new_n226), .ZN(new_n359));
  OAI21_X1  g0159(.A(KEYINPUT7), .B1(new_n334), .B2(G20), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n359), .A2(G68), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n355), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n361), .A2(new_n362), .A3(KEYINPUT16), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n356), .A2(new_n363), .A3(new_n264), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n339), .A2(G190), .A3(new_n301), .A4(new_n340), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n329), .A2(new_n342), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n366), .A2(KEYINPUT17), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n334), .A2(G20), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n344), .B1(new_n368), .B2(new_n345), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n355), .B1(new_n369), .B2(new_n360), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n273), .B1(new_n370), .B2(KEYINPUT16), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n371), .A2(new_n356), .B1(new_n326), .B2(new_n328), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n372), .A2(KEYINPUT80), .A3(new_n342), .A4(new_n365), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT80), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n366), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n367), .B1(new_n376), .B2(KEYINPUT17), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n341), .A2(G169), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(new_n317), .B2(new_n341), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n329), .A2(new_n364), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g0181(.A(new_n381), .B(KEYINPUT18), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n287), .A2(G232), .A3(new_n288), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n287), .A2(G238), .A3(G1698), .ZN(new_n385));
  INV_X1    g0185(.A(G107), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n384), .B(new_n385), .C1(new_n386), .C2(new_n287), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n296), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n303), .A2(G244), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(new_n301), .A3(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n390), .A2(G179), .ZN(new_n391));
  INV_X1    g0191(.A(G169), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n391), .B1(new_n392), .B2(new_n390), .ZN(new_n393));
  INV_X1    g0193(.A(G77), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n267), .A2(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n267), .A2(new_n264), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n270), .A2(new_n396), .A3(G77), .ZN(new_n397));
  XOR2_X1   g0197(.A(KEYINPUT8), .B(G58), .Z(new_n398));
  AOI22_X1  g0198(.A1(new_n398), .A2(new_n252), .B1(G20), .B2(G77), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT73), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  XOR2_X1   g0202(.A(KEYINPUT15), .B(G87), .Z(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n404), .A2(new_n261), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n399), .A2(new_n400), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n402), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  AND3_X1   g0208(.A1(new_n408), .A2(KEYINPUT74), .A3(new_n264), .ZN(new_n409));
  AOI21_X1  g0209(.A(KEYINPUT74), .B1(new_n408), .B2(new_n264), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n395), .B(new_n397), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n393), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(G190), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n390), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n300), .B1(new_n387), .B2(new_n296), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n311), .B1(new_n415), .B2(new_n389), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n408), .A2(new_n264), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT74), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n408), .A2(KEYINPUT74), .A3(new_n264), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n417), .A2(new_n422), .A3(new_n395), .A4(new_n397), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n383), .A2(new_n412), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT14), .ZN(new_n425));
  NAND2_X1  g0225(.A1(G33), .A2(G97), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n220), .A2(new_n288), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(G232), .B2(new_n288), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n426), .B1(new_n428), .B2(new_n286), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n296), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT76), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n303), .A2(G238), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n431), .B1(new_n432), .B2(new_n301), .ZN(new_n433));
  AOI211_X1 g0233(.A(KEYINPUT76), .B(new_n300), .C1(new_n303), .C2(G238), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n430), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT13), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT13), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n437), .B(new_n430), .C1(new_n433), .C2(new_n434), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n425), .B1(new_n439), .B2(G169), .ZN(new_n440));
  AOI211_X1 g0240(.A(KEYINPUT14), .B(new_n392), .C1(new_n436), .C2(new_n438), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n439), .A2(new_n317), .ZN(new_n442));
  OR3_X1    g0242(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n260), .A2(G77), .B1(G20), .B2(new_n344), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(new_n219), .B2(new_n253), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n445), .A2(KEYINPUT11), .A3(new_n264), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n445), .A2(new_n264), .ZN(new_n447));
  OR2_X1    g0247(.A1(new_n447), .A2(KEYINPUT11), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n275), .A2(G20), .A3(new_n344), .ZN(new_n449));
  XNOR2_X1  g0249(.A(new_n449), .B(KEYINPUT12), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n270), .A2(new_n396), .A3(G68), .ZN(new_n451));
  AND4_X1   g0251(.A1(new_n446), .A2(new_n448), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n443), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n452), .B1(new_n439), .B2(new_n413), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n311), .B1(new_n436), .B2(new_n438), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  NOR3_X1   g0259(.A1(new_n320), .A2(new_n424), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT88), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n226), .A2(G87), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n461), .B1(new_n358), .B2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n334), .A2(KEYINPUT88), .A3(new_n226), .A4(G87), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(KEYINPUT22), .A3(new_n464), .ZN(new_n465));
  OR3_X1    g0265(.A1(new_n286), .A2(KEYINPUT22), .A3(new_n462), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n386), .A2(G20), .ZN(new_n468));
  XOR2_X1   g0268(.A(new_n468), .B(KEYINPUT23), .Z(new_n469));
  NAND3_X1  g0269(.A1(new_n226), .A2(G33), .A3(G116), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n467), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT24), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n467), .A2(KEYINPUT24), .A3(new_n469), .A4(new_n470), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n473), .A2(new_n264), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(G41), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(KEYINPUT5), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n265), .A2(G45), .ZN(new_n478));
  OAI21_X1  g0278(.A(KEYINPUT83), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n476), .A2(KEYINPUT5), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT5), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G41), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT83), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n482), .A2(new_n483), .A3(new_n265), .A4(G45), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n479), .A2(new_n480), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n485), .A2(G264), .A3(new_n302), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n209), .A2(new_n288), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n211), .A2(G1698), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n334), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(G33), .A2(G294), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n302), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n479), .A2(new_n484), .A3(G274), .A4(new_n480), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n493), .A2(new_n296), .ZN(new_n494));
  NOR3_X1   g0294(.A1(new_n487), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G190), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n396), .B1(G1), .B2(new_n259), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G107), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n266), .A2(new_n468), .ZN(new_n500));
  XNOR2_X1  g0300(.A(new_n500), .B(KEYINPUT25), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n475), .A2(new_n496), .A3(new_n499), .A4(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n495), .A2(new_n311), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT84), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n485), .A2(G257), .A3(new_n302), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n506), .A2(new_n494), .ZN(new_n507));
  XNOR2_X1  g0307(.A(KEYINPUT82), .B(KEYINPUT4), .ZN(new_n508));
  INV_X1    g0308(.A(G244), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n509), .A2(G1698), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n508), .B1(new_n334), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G33), .A2(G283), .ZN(new_n512));
  AND2_X1   g0312(.A1(G250), .A2(G1698), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n513), .B1(new_n510), .B2(KEYINPUT4), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n512), .B1(new_n514), .B2(new_n286), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n296), .B1(new_n511), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n505), .B1(new_n507), .B2(new_n516), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n479), .A2(new_n484), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n518), .A2(G274), .A3(new_n302), .A4(new_n480), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n485), .A2(G257), .A3(new_n302), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n516), .A2(new_n519), .A3(new_n505), .A4(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n392), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n507), .A2(new_n317), .A3(new_n516), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n497), .A2(new_n210), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n252), .A2(G77), .ZN(new_n527));
  AND2_X1   g0327(.A1(KEYINPUT81), .A2(G97), .ZN(new_n528));
  NOR2_X1   g0328(.A1(KEYINPUT81), .A2(G97), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n530), .A2(KEYINPUT6), .A3(new_n386), .ZN(new_n531));
  XOR2_X1   g0331(.A(G97), .B(G107), .Z(new_n532));
  OAI21_X1  g0332(.A(new_n531), .B1(KEYINPUT6), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(G20), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n346), .A2(new_n347), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n527), .B(new_n534), .C1(new_n535), .C2(new_n386), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n526), .B1(new_n536), .B2(new_n264), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(G97), .B2(new_n276), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n524), .A2(new_n525), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n478), .A2(new_n209), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n302), .B(new_n540), .C1(G274), .C2(new_n478), .ZN(new_n541));
  NOR2_X1   g0341(.A1(G238), .A2(G1698), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n542), .B1(new_n509), .B2(G1698), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n334), .A2(new_n543), .B1(G33), .B2(G116), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n541), .B1(new_n544), .B2(new_n302), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n317), .ZN(new_n547));
  AOI21_X1  g0347(.A(KEYINPUT19), .B1(new_n530), .B2(new_n260), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT19), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n226), .B1(new_n426), .B2(new_n549), .ZN(new_n550));
  XNOR2_X1  g0350(.A(KEYINPUT81), .B(G97), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n551), .A2(new_n208), .A3(new_n386), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n548), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n334), .A2(new_n226), .A3(G68), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT85), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n334), .A2(KEYINPUT85), .A3(new_n226), .A4(G68), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n553), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n558), .A2(new_n264), .B1(new_n267), .B2(new_n404), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n498), .A2(new_n403), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n559), .A2(new_n560), .B1(new_n392), .B2(new_n545), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n498), .A2(G87), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  MUX2_X1   g0363(.A(new_n413), .B(new_n311), .S(new_n545), .Z(new_n564));
  AOI22_X1  g0364(.A1(new_n547), .A2(new_n561), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n276), .A2(G97), .ZN(new_n566));
  AOI211_X1 g0366(.A(new_n566), .B(new_n526), .C1(new_n536), .C2(new_n264), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n516), .A2(new_n519), .A3(new_n520), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(G200), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n567), .B(new_n569), .C1(new_n523), .C2(new_n413), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n539), .A2(new_n565), .A3(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n504), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(G116), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n263), .A2(new_n225), .B1(G20), .B2(new_n573), .ZN(new_n574));
  NOR3_X1   g0374(.A1(new_n528), .A2(new_n529), .A3(G33), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n512), .A2(new_n226), .ZN(new_n576));
  OAI211_X1 g0376(.A(KEYINPUT20), .B(new_n574), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(KEYINPUT86), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT20), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n575), .A2(new_n576), .ZN(new_n580));
  INV_X1    g0380(.A(new_n574), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n226), .B(new_n512), .C1(new_n551), .C2(G33), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT86), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n583), .A2(new_n584), .A3(KEYINPUT20), .A4(new_n574), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n578), .A2(new_n582), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n275), .A2(G20), .A3(new_n573), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n498), .A2(G116), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT87), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n586), .A2(KEYINPUT87), .A3(new_n588), .A4(new_n587), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n485), .A2(new_n302), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n494), .B1(new_n594), .B2(G270), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n211), .A2(new_n288), .ZN(new_n596));
  OR2_X1    g0396(.A1(new_n288), .A2(G264), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n357), .A2(new_n283), .A3(new_n596), .A4(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n286), .A2(G303), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n296), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n595), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n593), .A2(G169), .A3(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT21), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n485), .A2(G270), .A3(new_n302), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n601), .A2(new_n519), .A3(G179), .A4(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n593), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n392), .B1(new_n591), .B2(new_n592), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n610), .A2(KEYINPUT21), .A3(new_n602), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n605), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n475), .A2(new_n499), .A3(new_n501), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n495), .A2(G169), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n614), .B1(new_n317), .B2(new_n495), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n602), .A2(G200), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n595), .A2(G190), .A3(new_n601), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n618), .A2(new_n591), .A3(new_n592), .A4(new_n619), .ZN(new_n620));
  AND4_X1   g0420(.A1(new_n460), .A2(new_n572), .A3(new_n617), .A4(new_n620), .ZN(G372));
  INV_X1    g0421(.A(new_n319), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT18), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT90), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n379), .A2(new_n380), .A3(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n624), .B1(new_n379), .B2(new_n380), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n623), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n381), .A2(KEYINPUT90), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n629), .A2(KEYINPUT18), .A3(new_n625), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n412), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n443), .A2(new_n453), .B1(new_n458), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n631), .B1(new_n633), .B2(new_n377), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n622), .B1(new_n634), .B2(new_n316), .ZN(new_n635));
  INV_X1    g0435(.A(new_n460), .ZN(new_n636));
  OAI21_X1  g0436(.A(KEYINPUT89), .B1(new_n612), .B2(new_n616), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n610), .A2(KEYINPUT21), .A3(new_n602), .ZN(new_n638));
  AOI21_X1  g0438(.A(KEYINPUT21), .B1(new_n610), .B2(new_n602), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT89), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n613), .A2(new_n615), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n640), .A2(new_n641), .A3(new_n609), .A4(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n637), .A2(new_n643), .A3(new_n572), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n561), .A2(new_n547), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n563), .A2(new_n564), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT26), .ZN(new_n648));
  OR3_X1    g0448(.A1(new_n539), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n648), .B1(new_n539), .B2(new_n647), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n649), .A2(new_n650), .B1(new_n547), .B2(new_n561), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n644), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n635), .B1(new_n636), .B2(new_n653), .ZN(G369));
  OR3_X1    g0454(.A1(new_n266), .A2(KEYINPUT27), .A3(G20), .ZN(new_n655));
  OAI21_X1  g0455(.A(KEYINPUT27), .B1(new_n266), .B2(G20), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(G213), .A3(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(G343), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n593), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g0460(.A(new_n612), .B(new_n660), .Z(new_n661));
  NAND3_X1  g0461(.A1(new_n661), .A2(G330), .A3(new_n620), .ZN(new_n662));
  INV_X1    g0462(.A(new_n659), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n616), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n504), .B1(new_n613), .B2(new_n659), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n664), .B1(new_n665), .B2(new_n616), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n665), .A2(new_n612), .A3(new_n642), .A4(new_n663), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n664), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n667), .A2(new_n669), .ZN(G399));
  OR2_X1    g0470(.A1(new_n552), .A2(G116), .ZN(new_n671));
  XOR2_X1   g0471(.A(new_n671), .B(KEYINPUT91), .Z(new_n672));
  INV_X1    g0472(.A(new_n204), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(G41), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n672), .A2(G1), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(new_n230), .B2(new_n675), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT28), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT30), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n544), .A2(new_n302), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n490), .A2(new_n491), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n296), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n680), .A2(new_n682), .A3(new_n541), .A4(new_n486), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n517), .B2(new_n522), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT92), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n595), .A2(new_n686), .A3(G179), .A4(new_n601), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n607), .A2(KEYINPUT92), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n679), .B1(new_n685), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n568), .A2(KEYINPUT84), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n683), .B1(new_n691), .B2(new_n521), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n692), .A2(KEYINPUT30), .A3(new_n688), .A4(new_n687), .ZN(new_n693));
  INV_X1    g0493(.A(new_n495), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n546), .A2(G179), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n694), .A2(new_n568), .A3(new_n602), .A4(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n690), .A2(new_n693), .A3(new_n696), .ZN(new_n697));
  AND3_X1   g0497(.A1(new_n697), .A2(KEYINPUT31), .A3(new_n659), .ZN(new_n698));
  AOI21_X1  g0498(.A(KEYINPUT31), .B1(new_n697), .B2(new_n659), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT93), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n699), .A2(new_n700), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(KEYINPUT94), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT94), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n697), .A2(new_n659), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT31), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n697), .A2(KEYINPUT31), .A3(new_n659), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n705), .B(new_n702), .C1(new_n710), .C2(new_n700), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n617), .A2(new_n572), .A3(new_n620), .A4(new_n663), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n704), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  AND3_X1   g0513(.A1(new_n713), .A2(KEYINPUT95), .A3(G330), .ZN(new_n714));
  AOI21_X1  g0514(.A(KEYINPUT95), .B1(new_n713), .B2(G330), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT29), .ZN(new_n717));
  INV_X1    g0517(.A(new_n572), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n651), .B1(new_n718), .B2(new_n617), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n717), .B1(new_n719), .B2(new_n663), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n653), .A2(new_n659), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n720), .B1(new_n721), .B2(new_n717), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n716), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n678), .B1(new_n724), .B2(G1), .ZN(G364));
  AOI21_X1  g0525(.A(new_n225), .B1(G20), .B2(new_n392), .ZN(new_n726));
  NOR2_X1   g0526(.A1(G13), .A2(G33), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(G20), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n334), .A2(new_n673), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(G45), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n731), .B1(new_n732), .B2(new_n231), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n245), .A2(G45), .ZN(new_n734));
  AOI22_X1  g0534(.A1(new_n733), .A2(new_n734), .B1(new_n573), .B2(new_n673), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n287), .A2(G355), .A3(new_n204), .ZN(new_n736));
  AOI211_X1 g0536(.A(new_n726), .B(new_n729), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n274), .A2(G20), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n265), .B1(new_n738), .B2(G45), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n674), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n661), .A2(new_n620), .ZN(new_n743));
  AOI211_X1 g0543(.A(new_n737), .B(new_n742), .C1(new_n743), .C2(new_n729), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G179), .A2(G200), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n226), .B1(new_n745), .B2(G190), .ZN(new_n746));
  INV_X1    g0546(.A(G294), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n226), .A2(new_n413), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n750), .A2(new_n317), .A3(G200), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n317), .A2(new_n311), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n226), .A2(G190), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  XNOR2_X1  g0555(.A(KEYINPUT33), .B(G317), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n751), .A2(G322), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  XOR2_X1   g0557(.A(new_n757), .B(KEYINPUT98), .Z(new_n758));
  NOR2_X1   g0558(.A1(new_n311), .A2(G179), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n749), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G303), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n749), .A2(new_n752), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n287), .B1(new_n764), .B2(G326), .ZN(new_n765));
  INV_X1    g0565(.A(new_n753), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n766), .A2(new_n317), .A3(G200), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n753), .A2(new_n745), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n767), .A2(G311), .B1(G329), .B2(new_n769), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n758), .A2(new_n762), .A3(new_n765), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n759), .A2(new_n753), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n748), .B(new_n771), .C1(G283), .C2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n767), .ZN(new_n775));
  OR2_X1    g0575(.A1(new_n775), .A2(KEYINPUT96), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(KEYINPUT96), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G77), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n773), .A2(G107), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n746), .A2(KEYINPUT97), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n746), .A2(KEYINPUT97), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G97), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n760), .A2(new_n208), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n780), .A2(new_n781), .A3(new_n787), .A4(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G159), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n768), .A2(KEYINPUT32), .A3(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n754), .A2(new_n344), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n286), .B1(new_n751), .B2(G58), .ZN(new_n794));
  OAI21_X1  g0594(.A(KEYINPUT32), .B1(new_n768), .B2(new_n791), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n794), .B(new_n795), .C1(new_n219), .C2(new_n763), .ZN(new_n796));
  NOR4_X1   g0596(.A1(new_n790), .A2(new_n792), .A3(new_n793), .A4(new_n796), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n726), .B1(new_n774), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n744), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G330), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n743), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n801), .A2(new_n662), .A3(new_n742), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n799), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(G396));
  NAND2_X1  g0604(.A1(new_n411), .A2(new_n659), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n412), .A2(new_n423), .A3(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT100), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n412), .A2(new_n423), .A3(new_n805), .A4(KEYINPUT100), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n652), .A2(new_n663), .A3(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n808), .A2(new_n809), .B1(new_n632), .B2(new_n659), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n812), .B1(new_n721), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n742), .B1(new_n716), .B2(new_n815), .ZN(new_n816));
  OR2_X1    g0616(.A1(new_n816), .A2(KEYINPUT101), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n716), .A2(new_n815), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n816), .A2(KEYINPUT101), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(G132), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n334), .B1(new_n821), .B2(new_n768), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n751), .A2(G143), .B1(G150), .B2(new_n755), .ZN(new_n823));
  INV_X1    g0623(.A(G137), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n823), .B1(new_n824), .B2(new_n763), .C1(new_n778), .C2(new_n791), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT34), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n825), .A2(new_n826), .B1(new_n344), .B2(new_n772), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n822), .B(new_n827), .C1(new_n826), .C2(new_n825), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n828), .B1(new_n219), .B2(new_n760), .C1(new_n255), .C2(new_n746), .ZN(new_n829));
  INV_X1    g0629(.A(new_n751), .ZN(new_n830));
  INV_X1    g0630(.A(G283), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n830), .A2(new_n747), .B1(new_n754), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n779), .A2(G116), .ZN(new_n833));
  AOI22_X1  g0633(.A1(G107), .A2(new_n761), .B1(new_n773), .B2(G87), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n833), .A2(new_n286), .A3(new_n787), .A4(new_n834), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n832), .B(new_n835), .C1(G303), .C2(new_n764), .ZN(new_n836));
  INV_X1    g0636(.A(G311), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n836), .B1(new_n837), .B2(new_n768), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n829), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT99), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n742), .B1(new_n840), .B2(new_n726), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n726), .A2(new_n727), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n841), .B1(G77), .B2(new_n843), .C1(new_n728), .C2(new_n814), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n820), .A2(new_n844), .ZN(G384));
  INV_X1    g0645(.A(KEYINPUT40), .ZN(new_n846));
  INV_X1    g0646(.A(new_n657), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n370), .A2(KEYINPUT16), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n363), .A2(new_n264), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n328), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n327), .B1(new_n323), .B2(new_n324), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(KEYINPUT102), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT102), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n329), .B(new_n855), .C1(new_n849), .C2(new_n848), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n847), .B(new_n857), .C1(new_n377), .C2(new_n382), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n373), .A2(new_n375), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n378), .B(new_n657), .C1(new_n317), .C2(new_n341), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n854), .A2(new_n856), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(KEYINPUT37), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT37), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n380), .A2(new_n847), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n376), .A2(new_n863), .A3(new_n381), .A4(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  AND3_X1   g0666(.A1(new_n858), .A2(KEYINPUT38), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT38), .B1(new_n858), .B2(new_n866), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n698), .A2(new_n699), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n712), .A2(new_n870), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n453), .B(new_n659), .C1(new_n443), .C2(new_n457), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n452), .A2(new_n663), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  NOR3_X1   g0674(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n458), .B(new_n874), .C1(new_n875), .C2(new_n452), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n871), .A2(new_n814), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n846), .B1(new_n869), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT104), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n813), .B1(new_n712), .B2(new_n870), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n882), .B(new_n877), .C1(new_n867), .C2(new_n868), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n883), .A2(KEYINPUT104), .A3(new_n846), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT38), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n366), .B(new_n864), .C1(new_n626), .C2(new_n627), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT37), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n865), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n377), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n864), .B1(new_n891), .B2(new_n631), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n886), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n858), .A2(new_n866), .A3(KEYINPUT38), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n895), .A2(KEYINPUT40), .A3(new_n877), .A4(new_n882), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n885), .A2(new_n896), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n460), .A2(new_n871), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n897), .B(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(G330), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT105), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n635), .B1(new_n722), .B2(new_n636), .ZN(new_n902));
  XOR2_X1   g0702(.A(new_n901), .B(new_n902), .Z(new_n903));
  NAND2_X1  g0703(.A1(new_n858), .A2(new_n866), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n886), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n894), .ZN(new_n906));
  AOI211_X1 g0706(.A(new_n659), .B(new_n810), .C1(new_n644), .C2(new_n651), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n412), .A2(new_n659), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n906), .B(new_n877), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n628), .A2(new_n630), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n657), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT103), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n909), .A2(KEYINPUT103), .A3(new_n911), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT39), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n380), .B(new_n847), .C1(new_n910), .C2(new_n377), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT38), .B1(new_n917), .B2(new_n889), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n916), .B1(new_n918), .B2(new_n867), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n869), .A2(KEYINPUT39), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n454), .A2(new_n659), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n914), .A2(new_n915), .A3(new_n922), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n903), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n903), .A2(new_n923), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n924), .B(new_n925), .C1(new_n265), .C2(new_n738), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n573), .B1(new_n533), .B2(KEYINPUT35), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n927), .B(new_n227), .C1(KEYINPUT35), .C2(new_n533), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT36), .ZN(new_n929));
  OAI21_X1  g0729(.A(G77), .B1(new_n255), .B2(new_n344), .ZN(new_n930));
  OAI22_X1  g0730(.A1(new_n230), .A2(new_n930), .B1(G50), .B2(new_n344), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n931), .A2(G1), .A3(new_n274), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n926), .A2(new_n929), .A3(new_n932), .ZN(G367));
  OR2_X1    g0733(.A1(new_n539), .A2(new_n663), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n539), .B(new_n570), .C1(new_n567), .C2(new_n663), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  OR3_X1    g0737(.A1(new_n668), .A2(new_n937), .A3(KEYINPUT42), .ZN(new_n938));
  OAI21_X1  g0738(.A(KEYINPUT42), .B1(new_n668), .B2(new_n937), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n616), .A2(new_n570), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n940), .A2(new_n539), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n938), .B(new_n939), .C1(new_n659), .C2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n667), .A2(new_n936), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n563), .A2(new_n663), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n944), .A2(new_n547), .A3(new_n561), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n647), .B2(new_n944), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(KEYINPUT43), .ZN(new_n947));
  AND3_X1   g0747(.A1(new_n942), .A2(new_n943), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n943), .B1(new_n942), .B2(new_n947), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n946), .A2(KEYINPUT43), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  OR3_X1    g0751(.A1(new_n948), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n951), .B1(new_n948), .B2(new_n949), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n674), .B(KEYINPUT41), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n662), .A2(new_n668), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n612), .A2(new_n663), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n666), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(KEYINPUT107), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n958), .B(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n716), .A2(new_n722), .A3(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n669), .A2(new_n937), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT45), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n964), .B(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n667), .A2(KEYINPUT106), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n669), .ZN(new_n969));
  OAI21_X1  g0769(.A(KEYINPUT44), .B1(new_n969), .B2(new_n936), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT44), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n669), .A2(new_n971), .A3(new_n937), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NOR3_X1   g0773(.A1(new_n966), .A2(new_n968), .A3(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n963), .A2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n973), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n964), .B(KEYINPUT45), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n967), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n975), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n957), .B1(new_n980), .B2(new_n724), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n955), .B1(new_n981), .B2(new_n740), .ZN(new_n982));
  INV_X1    g0782(.A(G317), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n772), .A2(new_n551), .B1(new_n768), .B2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n746), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n984), .B1(G107), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n747), .B2(new_n754), .ZN(new_n987));
  INV_X1    g0787(.A(G303), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n830), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n763), .A2(new_n837), .ZN(new_n990));
  NOR4_X1   g0790(.A1(new_n987), .A2(new_n334), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n761), .A2(G116), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT46), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n991), .B(new_n993), .C1(new_n831), .C2(new_n778), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT109), .Z(new_n995));
  NAND2_X1  g0795(.A1(new_n786), .A2(G68), .ZN(new_n996));
  XOR2_X1   g0796(.A(KEYINPUT110), .B(G137), .Z(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n996), .B1(new_n251), .B2(new_n830), .C1(new_n768), .C2(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(G159), .B2(new_n755), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n773), .A2(G77), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n764), .A2(G143), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n761), .A2(G58), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n287), .B1(new_n778), .B2(new_n219), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n995), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT47), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n726), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n945), .B(new_n729), .C1(new_n647), .C2(new_n944), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n729), .A2(new_n726), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1010), .B1(new_n204), .B2(new_n404), .C1(new_n236), .C2(new_n731), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n741), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT108), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1008), .A2(new_n1009), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n982), .A2(new_n1014), .ZN(G387));
  NAND2_X1  g0815(.A1(new_n962), .A2(new_n740), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n287), .A2(new_n204), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n672), .A2(new_n1017), .B1(G107), .B2(new_n204), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT111), .Z(new_n1019));
  NAND2_X1  g0819(.A1(new_n241), .A2(G45), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n672), .B(new_n732), .C1(new_n344), .C2(new_n394), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT112), .Z(new_n1022));
  NAND2_X1  g0822(.A1(new_n398), .A2(new_n219), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT50), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1020), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1019), .B1(new_n1025), .B2(new_n731), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n742), .B1(new_n1026), .B2(new_n1010), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT113), .Z(new_n1028));
  NOR2_X1   g0828(.A1(new_n785), .A2(new_n404), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(G68), .B2(new_n767), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n219), .B2(new_n830), .C1(new_n210), .C2(new_n772), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(G159), .B2(new_n764), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n761), .A2(G77), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(KEYINPUT114), .B(G150), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n769), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n358), .B1(new_n322), .B2(new_n755), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1032), .A2(new_n1033), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n751), .A2(G317), .B1(G311), .B2(new_n755), .ZN(new_n1038));
  INV_X1    g0838(.A(G322), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1038), .B1(new_n1039), .B2(new_n763), .C1(new_n778), .C2(new_n988), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT48), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(new_n831), .B2(new_n746), .C1(new_n747), .C2(new_n760), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT49), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n769), .A2(G326), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n773), .A2(G116), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1044), .A2(new_n358), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1037), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n1049), .A2(new_n726), .B1(new_n666), .B2(new_n729), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1028), .A2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n724), .A2(new_n962), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n674), .B(KEYINPUT115), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n963), .A2(new_n1054), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1016), .B(new_n1051), .C1(new_n1052), .C2(new_n1055), .ZN(G393));
  OAI211_X1 g0856(.A(new_n977), .B(new_n976), .C1(new_n662), .C2(new_n666), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n667), .B1(new_n966), .B2(new_n973), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n963), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n980), .A2(new_n1060), .A3(new_n1054), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1057), .A2(new_n740), .A3(new_n1058), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n742), .B1(new_n937), .B2(new_n729), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1010), .B1(new_n204), .B2(new_n551), .C1(new_n248), .C2(new_n731), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n358), .B1(new_n779), .B2(new_n398), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n769), .A2(G143), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n751), .A2(G159), .B1(new_n764), .B2(G150), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1065), .B(new_n1066), .C1(KEYINPUT51), .C2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n754), .A2(new_n219), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n760), .A2(new_n344), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n785), .A2(new_n394), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(KEYINPUT51), .B2(new_n1067), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n208), .B2(new_n772), .ZN(new_n1073));
  NOR4_X1   g0873(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .A4(new_n1073), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n751), .A2(G311), .B1(new_n764), .B2(G317), .ZN(new_n1075));
  XOR2_X1   g0875(.A(new_n1075), .B(KEYINPUT52), .Z(new_n1076));
  NAND2_X1  g0876(.A1(new_n985), .A2(G116), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n760), .A2(new_n831), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n754), .A2(new_n988), .B1(new_n768), .B2(new_n1039), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1078), .B(new_n1079), .C1(G294), .C2(new_n767), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1076), .A2(new_n286), .A3(new_n1077), .A4(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(G107), .B2(new_n773), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n726), .B1(new_n1074), .B2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1063), .A2(new_n1064), .A3(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1061), .A2(new_n1062), .A3(new_n1084), .ZN(G390));
  NAND2_X1  g0885(.A1(new_n919), .A2(new_n920), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n877), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n908), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1087), .B1(new_n812), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1086), .B1(new_n921), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n921), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n895), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n719), .A2(new_n663), .A3(new_n811), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1087), .B1(new_n1093), .B2(new_n1088), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1090), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n882), .A2(G330), .A3(new_n877), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n814), .B(new_n877), .C1(new_n714), .C2(new_n715), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1099), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n740), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1086), .A2(new_n727), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n726), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n287), .B1(new_n998), .B2(new_n754), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n761), .A2(new_n1034), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT53), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1106), .A2(new_n1107), .B1(G50), .B2(new_n773), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n1107), .B2(new_n1106), .ZN(new_n1109));
  XOR2_X1   g0909(.A(KEYINPUT54), .B(G143), .Z(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT116), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1109), .B1(new_n779), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n791), .B2(new_n785), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n1105), .B(new_n1113), .C1(G125), .C2(new_n769), .ZN(new_n1114));
  INV_X1    g0914(.A(G128), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1114), .B1(new_n1115), .B2(new_n763), .C1(new_n821), .C2(new_n830), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n778), .A2(new_n551), .B1(new_n344), .B2(new_n772), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n1071), .B(new_n1117), .C1(G107), .C2(new_n755), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n751), .A2(G116), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n764), .A2(G283), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n287), .B(new_n788), .C1(G294), .C2(new_n769), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .A4(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1104), .B1(new_n1116), .B2(new_n1122), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n742), .B(new_n1123), .C1(new_n258), .C2(new_n842), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1103), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n877), .B1(new_n882), .B2(G330), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n1093), .A2(new_n1088), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1100), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1098), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n814), .B1(new_n714), .B2(new_n715), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1130), .B1(new_n1131), .B2(new_n1087), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n812), .A2(new_n1088), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1129), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n898), .A2(G330), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n902), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1140), .A2(new_n1101), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1130), .B1(new_n1090), .B2(new_n1096), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1097), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1100), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1142), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1054), .B1(new_n1139), .B2(new_n1145), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1102), .B(new_n1125), .C1(new_n1141), .C2(new_n1146), .ZN(G378));
  INV_X1    g0947(.A(KEYINPUT57), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n883), .A2(KEYINPUT104), .A3(new_n846), .ZN(new_n1149));
  AOI21_X1  g0949(.A(KEYINPUT104), .B1(new_n883), .B2(new_n846), .ZN(new_n1150));
  OAI211_X1 g0950(.A(G330), .B(new_n896), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1151));
  XOR2_X1   g0951(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n320), .B(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n281), .A2(new_n847), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1154), .B(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1151), .A2(new_n1157), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n885), .A2(G330), .A3(new_n1156), .A4(new_n896), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT119), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n923), .A2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1160), .B(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1138), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(new_n1101), .B2(new_n1135), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1148), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1160), .B(new_n923), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n713), .A2(G330), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT95), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n713), .A2(KEYINPUT95), .A3(G330), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n813), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1098), .B1(new_n1172), .B2(new_n877), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1126), .B1(new_n1172), .B2(new_n877), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n1133), .A2(new_n1173), .B1(new_n1174), .B2(new_n1128), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1138), .B1(new_n1175), .B2(new_n1145), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1167), .A2(KEYINPUT57), .A3(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1166), .A2(new_n1054), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n357), .A2(G33), .ZN(new_n1179));
  AOI21_X1  g0979(.A(G50), .B1(new_n1179), .B2(new_n476), .ZN(new_n1180));
  AOI21_X1  g0980(.A(G41), .B1(new_n751), .B2(G107), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n772), .A2(new_n255), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1182), .A2(new_n334), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1181), .A2(new_n1033), .A3(new_n1183), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n996), .B1(new_n210), .B2(new_n754), .C1(new_n831), .C2(new_n768), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n1184), .B(new_n1185), .C1(new_n403), .C2(new_n767), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n573), .B2(new_n763), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT117), .Z(new_n1188));
  INV_X1    g0988(.A(KEYINPUT58), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1180), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n1190), .B(KEYINPUT118), .Z(new_n1191));
  OAI22_X1  g0991(.A1(new_n830), .A2(new_n1115), .B1(new_n754), .B2(new_n821), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n764), .A2(G125), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n785), .B2(new_n251), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1192), .B(new_n1194), .C1(new_n761), .C2(new_n1111), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n824), .B2(new_n775), .ZN(new_n1196));
  OR2_X1    g0996(.A1(new_n1196), .A2(KEYINPUT59), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n773), .A2(G159), .ZN(new_n1198));
  AOI21_X1  g0998(.A(G41), .B1(new_n769), .B2(G124), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1197), .A2(new_n259), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1200));
  AND2_X1   g1000(.A1(new_n1196), .A2(KEYINPUT59), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n1188), .A2(new_n1189), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n726), .B1(new_n1191), .B2(new_n1202), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1203), .B(new_n741), .C1(G50), .C2(new_n843), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(new_n1157), .B2(new_n727), .ZN(new_n1205));
  AND3_X1   g1005(.A1(new_n909), .A2(KEYINPUT103), .A3(new_n911), .ZN(new_n1206));
  AOI21_X1  g1006(.A(KEYINPUT103), .B1(new_n909), .B2(new_n911), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(KEYINPUT119), .B1(new_n1208), .B2(new_n922), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n1160), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1162), .A2(new_n1159), .A3(new_n1158), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1205), .B1(new_n1212), .B2(new_n740), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1178), .A2(new_n1213), .ZN(G375));
  NAND2_X1  g1014(.A1(new_n1087), .A2(new_n727), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n843), .A2(G68), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n785), .A2(new_n404), .B1(new_n830), .B2(new_n831), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n754), .A2(new_n573), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n286), .B1(new_n760), .B2(new_n210), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1001), .B1(new_n747), .B2(new_n763), .ZN(new_n1220));
  NOR4_X1   g1020(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .A4(new_n1220), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n1221), .B1(new_n386), .B2(new_n778), .C1(new_n988), .C2(new_n768), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n785), .A2(new_n219), .B1(new_n251), .B2(new_n775), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT120), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1182), .B(new_n1224), .C1(new_n751), .C2(new_n997), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1111), .A2(new_n755), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n358), .B1(G159), .B2(new_n761), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n769), .A2(G128), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n763), .A2(new_n821), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1222), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n742), .B(new_n1216), .C1(new_n1231), .C2(new_n726), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1135), .A2(new_n740), .B1(new_n1215), .B2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n956), .B1(new_n1135), .B2(new_n1138), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1233), .B1(new_n1140), .B2(new_n1234), .ZN(new_n1235));
  XOR2_X1   g1035(.A(new_n1235), .B(KEYINPUT121), .Z(G381));
  XNOR2_X1  g1036(.A(G375), .B(KEYINPUT122), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1237), .A2(G378), .ZN(new_n1238));
  INV_X1    g1038(.A(G384), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1055), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n724), .B2(new_n962), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1241), .A2(new_n803), .A3(new_n1016), .A4(new_n1051), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(G387), .A2(new_n1242), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(G381), .A2(G390), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1238), .A2(new_n1239), .A3(new_n1243), .A4(new_n1244), .ZN(G407));
  INV_X1    g1045(.A(G213), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(new_n1238), .B2(new_n658), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(G407), .ZN(G409));
  NAND3_X1  g1048(.A1(new_n982), .A2(new_n1014), .A3(G390), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(G393), .A2(G396), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1242), .A2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(G390), .B1(new_n982), .B2(new_n1014), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT126), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1242), .A2(new_n1251), .A3(new_n1254), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n1250), .A2(new_n1252), .B1(new_n1253), .B2(new_n1255), .ZN(new_n1256));
  AND3_X1   g1056(.A1(new_n1061), .A2(new_n1062), .A3(new_n1084), .ZN(new_n1257));
  NOR3_X1   g1057(.A1(new_n963), .A2(new_n978), .A3(new_n974), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n956), .B1(new_n1258), .B2(new_n723), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n954), .B1(new_n1259), .B2(new_n739), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1014), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1257), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1255), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1262), .A2(new_n1263), .A3(new_n1249), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1256), .A2(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1246), .A2(G343), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT60), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1267), .B1(new_n1135), .B2(new_n1138), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1173), .A2(new_n1133), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1269), .A2(KEYINPUT60), .A3(new_n1164), .A4(new_n1129), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1268), .A2(new_n1054), .A3(new_n1270), .A4(new_n1139), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1233), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n1239), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1271), .A2(G384), .A3(new_n1233), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1176), .A2(new_n956), .A3(new_n1212), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(KEYINPUT123), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1205), .B1(new_n1167), .B2(new_n740), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT123), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1176), .A2(new_n1212), .A3(new_n1279), .A4(new_n956), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1277), .A2(new_n1278), .A3(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(G378), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1178), .A2(G378), .A3(new_n1213), .ZN(new_n1284));
  AOI211_X1 g1084(.A(new_n1266), .B(new_n1275), .C1(new_n1283), .C2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT62), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1266), .ZN(new_n1287));
  INV_X1    g1087(.A(G2897), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1271), .A2(G384), .A3(new_n1233), .ZN(new_n1290));
  AOI21_X1  g1090(.A(G384), .B1(new_n1271), .B2(new_n1233), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1287), .A2(KEYINPUT125), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1289), .B1(new_n1292), .B2(new_n1294), .ZN(new_n1295));
  AND4_X1   g1095(.A1(new_n1273), .A2(new_n1274), .A3(new_n1289), .A4(new_n1294), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1266), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1298));
  OAI22_X1  g1098(.A1(new_n1285), .A2(new_n1286), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1300), .A2(new_n1286), .A3(new_n1287), .A4(new_n1292), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT61), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1265), .B1(new_n1299), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1300), .A2(new_n1287), .ZN(new_n1305));
  OAI22_X1  g1105(.A1(new_n1275), .A2(new_n1293), .B1(new_n1288), .B2(new_n1287), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1292), .A2(new_n1289), .A3(new_n1294), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1253), .A2(new_n1255), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1252), .A2(new_n982), .A3(new_n1014), .A4(G390), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1264), .A2(new_n1302), .A3(new_n1309), .A4(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(KEYINPUT127), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT127), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1256), .A2(new_n1313), .A3(new_n1302), .A4(new_n1264), .ZN(new_n1314));
  AOI22_X1  g1114(.A1(new_n1305), .A2(new_n1308), .B1(new_n1312), .B2(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(KEYINPUT63), .B1(new_n1285), .B2(KEYINPUT124), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT124), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT63), .ZN(new_n1318));
  OAI211_X1 g1118(.A(new_n1317), .B(new_n1318), .C1(new_n1305), .C2(new_n1275), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1315), .A2(new_n1316), .A3(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1304), .A2(new_n1320), .ZN(G405));
  XNOR2_X1  g1121(.A(G375), .B(G378), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n1275), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1323), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1322), .A2(new_n1275), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1265), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  OR2_X1    g1126(.A1(new_n1322), .A2(new_n1275), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1327), .A2(new_n1256), .A3(new_n1264), .A4(new_n1323), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1326), .A2(new_n1328), .ZN(G402));
endmodule


