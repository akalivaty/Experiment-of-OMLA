//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 1 0 0 0 0 1 1 0 1 0 1 0 0 0 1 0 1 1 0 0 1 0 0 1 0 0 0 1 0 0 0 1 0 0 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n842,
    new_n843, new_n844, new_n845, new_n847, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955;
  INV_X1    g000(.A(KEYINPUT74), .ZN(new_n202));
  AND3_X1   g001(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT24), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT64), .ZN(new_n209));
  AOI21_X1  g008(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT64), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n205), .A2(new_n209), .A3(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n214));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n215), .B1(new_n216), .B2(KEYINPUT23), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n218));
  NOR3_X1   g017(.A1(new_n218), .A2(G169gat), .A3(G176gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n214), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G169gat), .ZN(new_n221));
  INV_X1    g020(.A(G176gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n221), .A2(new_n222), .A3(KEYINPUT23), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n218), .B1(G169gat), .B2(G176gat), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT65), .A4(new_n215), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n213), .A2(new_n220), .A3(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT25), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n217), .A2(new_n219), .ZN(new_n229));
  NAND3_X1  g028(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n208), .B(new_n230), .C1(G183gat), .C2(G190gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n229), .A2(new_n231), .A3(new_n232), .A4(KEYINPUT25), .ZN(new_n233));
  NOR3_X1   g032(.A1(new_n203), .A2(new_n210), .A3(new_n204), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT25), .A4(new_n215), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT66), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n228), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G120gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G113gat), .ZN(new_n240));
  INV_X1    g039(.A(G113gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G120gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G127gat), .B(G134gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(G127gat), .ZN(new_n247));
  INV_X1    g046(.A(G134gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT68), .B(G127gat), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n249), .B1(new_n250), .B2(new_n248), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT1), .B1(new_n240), .B2(new_n242), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n246), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT70), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT70), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n255), .B(new_n246), .C1(new_n251), .C2(new_n252), .ZN(new_n256));
  AND2_X1   g055(.A1(G169gat), .A2(G176gat), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT26), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n257), .B1(new_n258), .B2(new_n216), .ZN(new_n259));
  OAI21_X1  g058(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n260));
  AND2_X1   g059(.A1(new_n260), .A2(KEYINPUT67), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(KEYINPUT67), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n259), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n206), .ZN(new_n264));
  INV_X1    g063(.A(G183gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT27), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT27), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(G183gat), .ZN(new_n268));
  INV_X1    g067(.A(G190gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n266), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n264), .B1(new_n270), .B2(KEYINPUT28), .ZN(new_n271));
  XNOR2_X1  g070(.A(KEYINPUT27), .B(G183gat), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT28), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n272), .A2(new_n273), .A3(new_n269), .ZN(new_n274));
  AND3_X1   g073(.A1(new_n263), .A2(new_n271), .A3(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n238), .A2(new_n254), .A3(new_n256), .A4(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n254), .A2(new_n256), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n227), .A2(new_n226), .B1(new_n233), .B2(new_n236), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n278), .B1(new_n279), .B2(new_n275), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT34), .ZN(new_n281));
  NAND2_X1  g080(.A1(G227gat), .A2(G233gat), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n277), .A2(new_n280), .A3(new_n281), .A4(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(KEYINPUT73), .ZN(new_n284));
  INV_X1    g083(.A(new_n282), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n277), .A2(new_n280), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n277), .A2(new_n280), .A3(KEYINPUT71), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n281), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n284), .B1(new_n290), .B2(KEYINPUT72), .ZN(new_n291));
  AND3_X1   g090(.A1(new_n277), .A2(new_n280), .A3(KEYINPUT71), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT71), .B1(new_n277), .B2(new_n280), .ZN(new_n293));
  NOR3_X1   g092(.A1(new_n292), .A2(new_n293), .A3(new_n285), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT72), .ZN(new_n295));
  NOR3_X1   g094(.A1(new_n294), .A2(new_n295), .A3(new_n281), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n202), .B1(new_n291), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n295), .B1(new_n294), .B2(new_n281), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n288), .A2(new_n289), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n299), .A2(KEYINPUT72), .A3(KEYINPUT34), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n298), .A2(KEYINPUT74), .A3(new_n300), .A4(new_n284), .ZN(new_n301));
  XOR2_X1   g100(.A(G15gat), .B(G43gat), .Z(new_n302));
  XNOR2_X1  g101(.A(G71gat), .B(G99gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n282), .B1(new_n277), .B2(new_n280), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n304), .B1(new_n305), .B2(KEYINPUT33), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT32), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  AOI221_X4 g108(.A(new_n307), .B1(KEYINPUT33), .B2(new_n304), .C1(new_n286), .C2(new_n285), .ZN(new_n310));
  OR2_X1    g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n297), .A2(new_n301), .A3(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT36), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n291), .A2(new_n296), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n309), .A2(new_n310), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n298), .A2(new_n300), .A3(new_n284), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n318), .A2(new_n311), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT73), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n283), .B(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n299), .A2(KEYINPUT34), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n321), .B1(new_n322), .B2(new_n295), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n315), .B1(new_n323), .B2(new_n300), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n313), .B1(new_n319), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n317), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT30), .ZN(new_n327));
  XNOR2_X1  g126(.A(G197gat), .B(G204gat), .ZN(new_n328));
  INV_X1    g127(.A(G211gat), .ZN(new_n329));
  OR2_X1    g128(.A1(KEYINPUT75), .A2(G218gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(KEYINPUT75), .A2(G218gat), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n328), .B1(new_n332), .B2(KEYINPUT22), .ZN(new_n333));
  XNOR2_X1  g132(.A(G211gat), .B(G218gat), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n328), .B(new_n334), .C1(new_n332), .C2(KEYINPUT22), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(G226gat), .A2(G233gat), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n275), .B1(new_n228), .B2(new_n237), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n339), .B1(new_n340), .B2(KEYINPUT29), .ZN(new_n341));
  INV_X1    g140(.A(new_n339), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n342), .B1(new_n279), .B2(new_n275), .ZN(new_n343));
  AOI211_X1 g142(.A(KEYINPUT76), .B(new_n338), .C1(new_n341), .C2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT76), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n341), .A2(new_n343), .ZN(new_n346));
  INV_X1    g145(.A(new_n338), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n238), .A2(new_n276), .ZN(new_n349));
  AOI21_X1  g148(.A(KEYINPUT77), .B1(new_n349), .B2(new_n342), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT77), .ZN(new_n351));
  NOR3_X1   g150(.A1(new_n340), .A2(new_n351), .A3(new_n339), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n338), .B(new_n341), .C1(new_n350), .C2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n344), .B1(new_n348), .B2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G8gat), .B(G36gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(G64gat), .B(G92gat), .ZN(new_n356));
  XOR2_X1   g155(.A(new_n355), .B(new_n356), .Z(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n327), .B1(new_n354), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n354), .A2(new_n358), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n348), .A2(new_n353), .ZN(new_n362));
  INV_X1    g161(.A(new_n344), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(new_n357), .ZN(new_n365));
  OAI21_X1  g164(.A(KEYINPUT78), .B1(new_n365), .B2(new_n327), .ZN(new_n366));
  NAND2_X1  g165(.A1(G225gat), .A2(G233gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(KEYINPUT81), .B(G155gat), .ZN(new_n369));
  INV_X1    g168(.A(G162gat), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT2), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(G141gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(KEYINPUT79), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT79), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(G141gat), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(new_n375), .A3(G148gat), .ZN(new_n376));
  INV_X1    g175(.A(G148gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(G141gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  AND2_X1   g178(.A1(new_n370), .A2(G155gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n370), .A2(G155gat), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT80), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G155gat), .B(G162gat), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT80), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n371), .A2(new_n379), .A3(new_n382), .A4(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G141gat), .B(G148gat), .ZN(new_n387));
  OAI22_X1  g186(.A1(new_n387), .A2(KEYINPUT2), .B1(new_n380), .B2(new_n381), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT82), .B1(new_n389), .B2(KEYINPUT3), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT83), .B(KEYINPUT3), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n386), .A2(new_n388), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n253), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT3), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n395), .B1(new_n386), .B2(new_n388), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT82), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n368), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT5), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT85), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT1), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n243), .A2(new_n401), .ZN(new_n402));
  AND2_X1   g201(.A1(new_n247), .A2(KEYINPUT68), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n247), .A2(KEYINPUT68), .ZN(new_n404));
  OAI21_X1  g203(.A(G134gat), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n402), .A2(new_n405), .A3(new_n249), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n386), .A2(new_n388), .A3(new_n406), .A4(new_n246), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n400), .B1(new_n407), .B2(KEYINPUT4), .ZN(new_n408));
  AND2_X1   g207(.A1(new_n386), .A2(new_n388), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n409), .A2(new_n254), .A3(new_n256), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n408), .B1(new_n410), .B2(KEYINPUT4), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n407), .A2(new_n400), .A3(KEYINPUT4), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n398), .A2(new_n399), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n389), .A2(new_n253), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n407), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n368), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n253), .B(new_n392), .C1(new_n396), .C2(KEYINPUT82), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n396), .A2(KEYINPUT82), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n367), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT4), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n407), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n421), .B1(new_n410), .B2(new_n420), .ZN(new_n422));
  OAI211_X1 g221(.A(KEYINPUT5), .B(new_n416), .C1(new_n419), .C2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n413), .A2(new_n423), .ZN(new_n424));
  XOR2_X1   g223(.A(G1gat), .B(G29gat), .Z(new_n425));
  XNOR2_X1  g224(.A(G57gat), .B(G85gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(KEYINPUT84), .B(KEYINPUT0), .ZN(new_n428));
  XOR2_X1   g227(.A(new_n427), .B(new_n428), .Z(new_n429));
  NAND2_X1  g228(.A1(new_n424), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT6), .ZN(new_n431));
  INV_X1    g230(.A(new_n429), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n413), .A2(new_n423), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n430), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n416), .A2(KEYINPUT5), .ZN(new_n435));
  INV_X1    g234(.A(new_n422), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n435), .B1(new_n398), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n411), .A2(new_n412), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n399), .B(new_n367), .C1(new_n417), .C2(new_n418), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI211_X1 g239(.A(KEYINPUT6), .B(new_n429), .C1(new_n437), .C2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n434), .A2(new_n441), .ZN(new_n442));
  NOR3_X1   g241(.A1(new_n354), .A2(new_n327), .A3(new_n358), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT78), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n361), .A2(new_n366), .A3(new_n442), .A4(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT29), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n338), .B1(new_n392), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(G228gat), .A2(G233gat), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n389), .A2(KEYINPUT3), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT86), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n338), .A2(new_n447), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n451), .B(new_n452), .C1(new_n453), .C2(new_n409), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT29), .B1(new_n336), .B2(new_n337), .ZN(new_n455));
  OAI211_X1 g254(.A(KEYINPUT86), .B(new_n389), .C1(new_n455), .C2(KEYINPUT3), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n450), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n409), .B1(new_n453), .B2(new_n391), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n449), .B1(new_n458), .B2(new_n448), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(G22gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(G78gat), .B(G106gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(KEYINPUT31), .B(G50gat), .ZN(new_n463));
  XOR2_X1   g262(.A(new_n462), .B(new_n463), .Z(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n465), .A2(KEYINPUT87), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n461), .B(new_n466), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n460), .A2(G22gat), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  OR2_X1    g268(.A1(new_n468), .A2(KEYINPUT88), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n464), .B1(new_n468), .B2(KEYINPUT88), .ZN(new_n471));
  AOI22_X1  g270(.A1(new_n467), .A2(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n446), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n326), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT89), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT37), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n364), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n358), .B1(new_n354), .B2(KEYINPUT37), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT38), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT90), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n441), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n424), .A2(KEYINPUT90), .A3(KEYINPUT6), .A4(new_n429), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT6), .B1(new_n424), .B2(new_n429), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n482), .A2(new_n483), .B1(new_n484), .B2(new_n433), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n477), .B1(new_n346), .B2(new_n338), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n347), .B(new_n341), .C1(new_n350), .C2(new_n352), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT38), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n358), .B(new_n488), .C1(new_n354), .C2(KEYINPUT37), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n480), .A2(new_n485), .A3(new_n365), .A4(new_n489), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n490), .A2(new_n472), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT40), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n411), .B(new_n412), .C1(new_n418), .C2(new_n417), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT39), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(new_n494), .A3(new_n368), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n432), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n414), .A2(new_n367), .A3(new_n407), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT39), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n498), .B1(new_n493), .B2(new_n368), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n492), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n499), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n501), .A2(KEYINPUT40), .A3(new_n432), .A4(new_n495), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n500), .A2(new_n502), .A3(new_n430), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n360), .B(new_n359), .C1(new_n443), .C2(new_n444), .ZN(new_n504));
  NOR3_X1   g303(.A1(new_n365), .A2(KEYINPUT78), .A3(new_n327), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n475), .A2(new_n476), .B1(new_n491), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n326), .A2(new_n474), .A3(KEYINPUT89), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n318), .A2(new_n311), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n323), .A2(new_n300), .A3(new_n315), .ZN(new_n510));
  AND3_X1   g309(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT91), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT91), .B1(new_n509), .B2(new_n510), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n472), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n504), .A2(new_n505), .ZN(new_n514));
  XNOR2_X1  g313(.A(KEYINPUT92), .B(KEYINPUT35), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n485), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  OR2_X1    g316(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n312), .A2(new_n510), .A3(new_n472), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT35), .B1(new_n519), .B2(new_n446), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n507), .A2(new_n508), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(G43gat), .B(G50gat), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n522), .A2(KEYINPUT15), .ZN(new_n523));
  NOR2_X1   g322(.A1(G29gat), .A2(G36gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n524), .B(KEYINPUT14), .ZN(new_n525));
  INV_X1    g324(.A(G29gat), .ZN(new_n526));
  INV_X1    g325(.A(G36gat), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT94), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR3_X1   g327(.A1(new_n523), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n522), .A2(KEYINPUT15), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT17), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT95), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n531), .B(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n533), .B1(new_n535), .B2(new_n532), .ZN(new_n536));
  INV_X1    g335(.A(G8gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(G15gat), .B(G22gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(KEYINPUT96), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n539), .A2(G1gat), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n537), .B1(new_n540), .B2(KEYINPUT97), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT16), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n539), .B1(new_n542), .B2(G1gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n541), .A2(new_n544), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n536), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(G229gat), .A2(G233gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n547), .A2(new_n535), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT18), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n547), .B(new_n535), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n550), .B(KEYINPUT13), .Z(new_n555));
  AOI22_X1  g354(.A1(new_n552), .A2(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n549), .A2(KEYINPUT18), .A3(new_n550), .A4(new_n551), .ZN(new_n557));
  XNOR2_X1  g356(.A(G113gat), .B(G141gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(KEYINPUT93), .B(G197gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(KEYINPUT11), .B(G169gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n562), .B(KEYINPUT12), .Z(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n556), .A2(new_n557), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n564), .B1(new_n556), .B2(new_n557), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n521), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G85gat), .A2(G92gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT7), .ZN(new_n571));
  NAND2_X1  g370(.A1(G99gat), .A2(G106gat), .ZN(new_n572));
  INV_X1    g371(.A(G85gat), .ZN(new_n573));
  INV_X1    g372(.A(G92gat), .ZN(new_n574));
  AOI22_X1  g373(.A1(KEYINPUT8), .A2(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G99gat), .B(G106gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n536), .A2(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(G190gat), .B(G218gat), .Z(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT100), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT101), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT41), .ZN(new_n584));
  NAND2_X1  g383(.A1(G232gat), .A2(G233gat), .ZN(new_n585));
  OAI22_X1  g384(.A1(new_n582), .A2(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n586), .B1(new_n535), .B2(new_n578), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n580), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n588), .A2(new_n583), .A3(new_n582), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n582), .A2(new_n583), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n580), .A2(new_n590), .A3(new_n587), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G134gat), .B(G162gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n585), .A2(new_n584), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n593), .B(new_n594), .Z(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n589), .A2(new_n595), .A3(new_n591), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT21), .ZN(new_n600));
  XOR2_X1   g399(.A(G57gat), .B(G64gat), .Z(new_n601));
  INV_X1    g400(.A(KEYINPUT9), .ZN(new_n602));
  INV_X1    g401(.A(G71gat), .ZN(new_n603));
  INV_X1    g402(.A(G78gat), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(G71gat), .B(G78gat), .Z(new_n607));
  OR2_X1    g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n548), .B1(new_n600), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n600), .ZN(new_n612));
  XOR2_X1   g411(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n611), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G127gat), .B(G155gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT99), .ZN(new_n617));
  NAND2_X1  g416(.A1(G231gat), .A2(G233gat), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n618), .B(KEYINPUT98), .Z(new_n619));
  XNOR2_X1  g418(.A(new_n617), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G183gat), .B(G211gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n615), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n615), .A2(new_n622), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n599), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n578), .A2(KEYINPUT10), .A3(new_n609), .A4(new_n608), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n578), .B(new_n610), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n627), .B1(new_n629), .B2(KEYINPUT10), .ZN(new_n630));
  AND2_X1   g429(.A1(G230gat), .A2(G233gat), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n633), .B1(new_n628), .B2(new_n632), .ZN(new_n634));
  XNOR2_X1  g433(.A(G120gat), .B(G148gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(G176gat), .B(G204gat), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n635), .B(new_n636), .Z(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n634), .A2(new_n638), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n626), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n569), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT102), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n569), .A2(KEYINPUT102), .A3(new_n642), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n442), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(G1gat), .ZN(G1324gat));
  NAND3_X1  g449(.A1(new_n361), .A2(new_n366), .A3(new_n445), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n537), .B1(new_n647), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT103), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(G8gat), .ZN(new_n654));
  AOI211_X1 g453(.A(new_n514), .B(new_n654), .C1(new_n645), .C2(new_n646), .ZN(new_n655));
  OAI21_X1  g454(.A(KEYINPUT42), .B1(new_n652), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n656), .B1(KEYINPUT42), .B2(new_n655), .ZN(G1325gat));
  INV_X1    g456(.A(new_n511), .ZN(new_n658));
  INV_X1    g457(.A(new_n512), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(G15gat), .B1(new_n647), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(KEYINPUT36), .B1(new_n318), .B2(new_n311), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n315), .B1(new_n318), .B2(new_n202), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n662), .B1(new_n301), .B2(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(KEYINPUT36), .B1(new_n509), .B2(new_n510), .ZN(new_n665));
  OAI21_X1  g464(.A(KEYINPUT104), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT104), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n317), .A2(new_n325), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(G15gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT105), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n661), .B1(new_n647), .B2(new_n671), .ZN(G1326gat));
  INV_X1    g471(.A(new_n646), .ZN(new_n673));
  AOI21_X1  g472(.A(KEYINPUT102), .B1(new_n569), .B2(new_n642), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n473), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(KEYINPUT106), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT106), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n647), .A2(new_n677), .A3(new_n473), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT43), .B(G22gat), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n676), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n679), .B1(new_n676), .B2(new_n678), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n680), .A2(new_n681), .ZN(G1327gat));
  INV_X1    g481(.A(new_n599), .ZN(new_n683));
  INV_X1    g482(.A(new_n625), .ZN(new_n684));
  INV_X1    g483(.A(new_n641), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n521), .A2(new_n568), .A3(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n687), .A2(new_n526), .A3(new_n648), .ZN(new_n688));
  XOR2_X1   g487(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n506), .A2(new_n490), .A3(new_n472), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n666), .A2(new_n691), .A3(new_n474), .A4(new_n668), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT110), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n520), .B1(new_n513), .B2(new_n517), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n693), .B1(new_n692), .B2(new_n694), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n599), .A2(KEYINPUT44), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n697), .A2(KEYINPUT111), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n692), .A2(new_n694), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(KEYINPUT110), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n692), .A2(new_n694), .A3(new_n693), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n701), .A2(new_n702), .A3(new_n698), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT111), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n507), .A2(new_n508), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(new_n694), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n683), .ZN(new_n708));
  AOI22_X1  g507(.A1(new_n699), .A2(new_n705), .B1(KEYINPUT44), .B2(new_n708), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n641), .B(KEYINPUT108), .Z(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n556), .A2(new_n557), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(new_n563), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n565), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n711), .A2(new_n714), .A3(new_n684), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT109), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n709), .A2(new_n442), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n690), .B1(new_n717), .B2(new_n526), .ZN(G1328gat));
  NAND3_X1  g517(.A1(new_n687), .A2(new_n527), .A3(new_n651), .ZN(new_n719));
  XOR2_X1   g518(.A(new_n719), .B(KEYINPUT46), .Z(new_n720));
  NOR3_X1   g519(.A1(new_n709), .A2(new_n514), .A3(new_n716), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT112), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(G36gat), .B1(new_n721), .B2(new_n722), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n720), .B1(new_n723), .B2(new_n724), .ZN(G1329gat));
  INV_X1    g524(.A(KEYINPUT47), .ZN(new_n726));
  INV_X1    g525(.A(G43gat), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n699), .A2(new_n705), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n708), .A2(KEYINPUT44), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n716), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n727), .B1(new_n730), .B2(new_n669), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n687), .A2(new_n727), .A3(new_n660), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n726), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n669), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n709), .A2(new_n735), .A3(new_n716), .ZN(new_n736));
  OAI211_X1 g535(.A(KEYINPUT47), .B(new_n732), .C1(new_n736), .C2(new_n727), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n734), .A2(new_n737), .ZN(G1330gat));
  INV_X1    g537(.A(KEYINPUT48), .ZN(new_n739));
  INV_X1    g538(.A(G50gat), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n740), .B1(new_n730), .B2(new_n473), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n472), .A2(G50gat), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n687), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n739), .B1(new_n741), .B2(new_n744), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n709), .A2(new_n472), .A3(new_n716), .ZN(new_n746));
  OAI211_X1 g545(.A(KEYINPUT48), .B(new_n743), .C1(new_n746), .C2(new_n740), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(G1331gat));
  NOR3_X1   g547(.A1(new_n711), .A2(new_n714), .A3(new_n626), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n697), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n648), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n651), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n753), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n754));
  XOR2_X1   g553(.A(KEYINPUT49), .B(G64gat), .Z(new_n755));
  OAI21_X1  g554(.A(new_n754), .B1(new_n753), .B2(new_n755), .ZN(G1333gat));
  NAND3_X1  g555(.A1(new_n750), .A2(new_n603), .A3(new_n660), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n750), .A2(new_n669), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n757), .B1(new_n758), .B2(new_n603), .ZN(new_n759));
  XNOR2_X1  g558(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n759), .B(new_n760), .Z(G1334gat));
  NAND2_X1  g560(.A1(new_n750), .A2(new_n473), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(G78gat), .ZN(G1335gat));
  AOI21_X1  g562(.A(KEYINPUT111), .B1(new_n697), .B2(new_n698), .ZN(new_n764));
  AND4_X1   g563(.A1(KEYINPUT111), .A2(new_n701), .A3(new_n702), .A4(new_n698), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n729), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n714), .A2(new_n625), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n641), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(G85gat), .B1(new_n770), .B2(new_n442), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n700), .A2(new_n683), .A3(new_n767), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT51), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n773), .A2(new_n685), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n774), .A2(new_n573), .A3(new_n648), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n771), .A2(new_n775), .ZN(G1336gat));
  NOR2_X1   g575(.A1(KEYINPUT115), .A2(KEYINPUT52), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n766), .A2(new_n651), .A3(new_n769), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(G92gat), .ZN(new_n780));
  NAND2_X1  g579(.A1(KEYINPUT115), .A2(KEYINPUT52), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n710), .A2(new_n574), .A3(new_n651), .ZN(new_n782));
  XOR2_X1   g581(.A(new_n782), .B(KEYINPUT114), .Z(new_n783));
  OAI21_X1  g582(.A(new_n781), .B1(new_n773), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n778), .B1(new_n780), .B2(new_n785), .ZN(new_n786));
  AOI211_X1 g585(.A(new_n784), .B(new_n777), .C1(new_n779), .C2(G92gat), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n786), .A2(new_n787), .ZN(G1337gat));
  OAI21_X1  g587(.A(G99gat), .B1(new_n770), .B2(new_n735), .ZN(new_n789));
  INV_X1    g588(.A(G99gat), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n774), .A2(new_n790), .A3(new_n660), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n789), .A2(new_n791), .ZN(G1338gat));
  INV_X1    g591(.A(G106gat), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n768), .B1(new_n728), .B2(new_n729), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n793), .B1(new_n794), .B2(new_n473), .ZN(new_n795));
  NOR4_X1   g594(.A1(new_n773), .A2(G106gat), .A3(new_n472), .A4(new_n711), .ZN(new_n796));
  OAI21_X1  g595(.A(KEYINPUT53), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(G106gat), .B1(new_n770), .B2(new_n472), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n799));
  INV_X1    g598(.A(new_n796), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n797), .A2(new_n801), .ZN(G1339gat));
  NOR3_X1   g601(.A1(new_n626), .A2(new_n714), .A3(new_n641), .ZN(new_n803));
  INV_X1    g602(.A(new_n633), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n637), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OR2_X1    g605(.A1(new_n630), .A2(new_n632), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n807), .A2(KEYINPUT54), .A3(new_n633), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n806), .A2(new_n808), .A3(KEYINPUT55), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n811), .A2(new_n639), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n813), .B1(new_n713), .B2(new_n565), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n554), .A2(new_n555), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n550), .B1(new_n549), .B2(new_n551), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n562), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n565), .A2(new_n641), .A3(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n599), .B1(new_n814), .B2(new_n819), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n565), .A2(new_n817), .ZN(new_n821));
  INV_X1    g620(.A(new_n813), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n683), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n803), .B1(new_n824), .B2(new_n684), .ZN(new_n825));
  NOR4_X1   g624(.A1(new_n825), .A2(new_n442), .A3(new_n651), .A4(new_n519), .ZN(new_n826));
  AOI21_X1  g625(.A(G113gat), .B1(new_n826), .B2(new_n714), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n714), .A2(new_n822), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n683), .B1(new_n828), .B2(new_n818), .ZN(new_n829));
  INV_X1    g628(.A(new_n823), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n684), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n803), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n513), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n833), .A2(new_n648), .A3(new_n514), .A4(new_n834), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(KEYINPUT116), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n568), .A2(new_n241), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n827), .B1(new_n836), .B2(new_n837), .ZN(G1340gat));
  AOI21_X1  g637(.A(G120gat), .B1(new_n826), .B2(new_n641), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n711), .A2(new_n239), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n839), .B1(new_n836), .B2(new_n840), .ZN(G1341gat));
  INV_X1    g640(.A(new_n836), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n842), .A2(new_n250), .A3(new_n684), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n826), .A2(new_n625), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n844), .B(KEYINPUT117), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n843), .B1(new_n845), .B2(new_n250), .ZN(G1342gat));
  NAND3_X1  g645(.A1(new_n826), .A2(new_n248), .A3(new_n683), .ZN(new_n847));
  XOR2_X1   g646(.A(new_n847), .B(KEYINPUT56), .Z(new_n848));
  OAI21_X1  g647(.A(G134gat), .B1(new_n842), .B2(new_n599), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(G1343gat));
  NAND2_X1  g649(.A1(new_n373), .A2(new_n375), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n852), .B1(new_n825), .B2(new_n472), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n809), .A2(KEYINPUT118), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT118), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n806), .A2(new_n808), .A3(new_n855), .ZN(new_n856));
  XNOR2_X1  g655(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n854), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n812), .A2(new_n639), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n818), .B1(new_n568), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n599), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n625), .B1(new_n862), .B2(new_n823), .ZN(new_n863));
  OAI211_X1 g662(.A(KEYINPUT57), .B(new_n473), .C1(new_n863), .C2(new_n803), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n853), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n714), .A2(new_n859), .A3(new_n858), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n683), .B1(new_n867), .B2(new_n818), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n684), .B1(new_n868), .B2(new_n830), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n472), .B1(new_n869), .B2(new_n832), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n870), .A2(KEYINPUT120), .A3(KEYINPUT57), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n669), .A2(new_n442), .A3(new_n651), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n866), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n851), .B1(new_n873), .B2(new_n568), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n651), .A2(new_n472), .ZN(new_n875));
  AND4_X1   g674(.A1(new_n648), .A2(new_n833), .A3(new_n735), .A4(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n876), .A2(new_n372), .A3(new_n714), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g677(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n874), .A2(new_n877), .A3(new_n879), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(G1344gat));
  NAND3_X1  g682(.A1(new_n833), .A2(KEYINPUT57), .A3(new_n473), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n884), .B1(KEYINPUT57), .B2(new_n870), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n885), .A2(new_n641), .A3(new_n872), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT59), .B1(new_n886), .B2(new_n377), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n866), .A2(new_n641), .A3(new_n871), .A4(new_n872), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT122), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n377), .A2(KEYINPUT59), .ZN(new_n890));
  AND3_X1   g689(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n889), .B1(new_n888), .B2(new_n890), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n887), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n876), .A2(new_n377), .A3(new_n641), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(G1345gat));
  NAND3_X1  g694(.A1(new_n876), .A2(new_n369), .A3(new_n625), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n873), .A2(new_n684), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n896), .B1(new_n897), .B2(new_n369), .ZN(G1346gat));
  NAND3_X1  g697(.A1(new_n876), .A2(new_n370), .A3(new_n683), .ZN(new_n899));
  XOR2_X1   g698(.A(new_n899), .B(KEYINPUT123), .Z(new_n900));
  OAI21_X1  g699(.A(G162gat), .B1(new_n873), .B2(new_n599), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(G1347gat));
  NOR3_X1   g701(.A1(new_n825), .A2(new_n648), .A3(new_n514), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n834), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n904), .A2(new_n221), .A3(new_n568), .ZN(new_n905));
  INV_X1    g704(.A(new_n519), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n714), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n905), .B1(new_n221), .B2(new_n909), .ZN(G1348gat));
  OAI21_X1  g709(.A(G176gat), .B1(new_n904), .B2(new_n711), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n641), .A2(new_n222), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n911), .B1(new_n907), .B2(new_n912), .ZN(G1349gat));
  OAI21_X1  g712(.A(G183gat), .B1(new_n904), .B2(new_n684), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n625), .A2(new_n272), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n914), .B1(new_n907), .B2(new_n915), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g716(.A1(new_n908), .A2(new_n269), .A3(new_n683), .ZN(new_n918));
  OAI21_X1  g717(.A(G190gat), .B1(new_n904), .B2(new_n599), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n919), .A2(KEYINPUT61), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n919), .A2(KEYINPUT61), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(G1351gat));
  NAND3_X1  g721(.A1(new_n735), .A2(new_n442), .A3(new_n651), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n885), .A2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(G197gat), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n925), .A2(new_n926), .A3(new_n568), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n825), .A2(new_n472), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(new_n924), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT124), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n928), .A2(KEYINPUT124), .A3(new_n924), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(new_n714), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n927), .B1(new_n934), .B2(new_n926), .ZN(G1352gat));
  NOR3_X1   g734(.A1(new_n929), .A2(G204gat), .A3(new_n685), .ZN(new_n936));
  XNOR2_X1  g735(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n936), .B(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(G204gat), .B1(new_n925), .B2(new_n711), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(G1353gat));
  OAI21_X1  g739(.A(G211gat), .B1(new_n925), .B2(new_n684), .ZN(new_n941));
  NOR2_X1   g740(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI221_X1 g742(.A(G211gat), .B1(KEYINPUT126), .B2(KEYINPUT63), .C1(new_n925), .C2(new_n684), .ZN(new_n944));
  NAND2_X1  g743(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n933), .A2(new_n329), .A3(new_n625), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(G1354gat));
  AOI211_X1 g747(.A(new_n599), .B(new_n925), .C1(new_n330), .C2(new_n331), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n931), .A2(new_n683), .A3(new_n932), .ZN(new_n950));
  INV_X1    g749(.A(G218gat), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT127), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n950), .A2(KEYINPUT127), .A3(new_n951), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n949), .B1(new_n954), .B2(new_n955), .ZN(G1355gat));
endmodule


