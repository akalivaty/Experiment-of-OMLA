

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U551 ( .A1(n544), .A2(n543), .ZN(n677) );
  XOR2_X1 U552 ( .A(KEYINPUT17), .B(n540), .Z(n880) );
  AND2_X2 U553 ( .A1(n536), .A2(G2104), .ZN(n879) );
  NOR2_X1 U554 ( .A1(n747), .A2(n765), .ZN(n516) );
  INV_X1 U555 ( .A(KEYINPUT26), .ZN(n689) );
  XNOR2_X1 U556 ( .A(n690), .B(n689), .ZN(n692) );
  XNOR2_X1 U557 ( .A(n716), .B(KEYINPUT30), .ZN(n717) );
  INV_X1 U558 ( .A(KEYINPUT102), .ZN(n720) );
  XNOR2_X1 U559 ( .A(n720), .B(KEYINPUT31), .ZN(n721) );
  XNOR2_X1 U560 ( .A(n722), .B(n721), .ZN(n723) );
  INV_X1 U561 ( .A(G40), .ZN(n676) );
  XNOR2_X1 U562 ( .A(n733), .B(KEYINPUT32), .ZN(n742) );
  NOR2_X2 U563 ( .A1(n769), .A2(n770), .ZN(n713) );
  NOR2_X1 U564 ( .A1(n758), .A2(n757), .ZN(n767) );
  NOR2_X1 U565 ( .A1(G651), .A2(n634), .ZN(n644) );
  XNOR2_X1 U566 ( .A(G543), .B(KEYINPUT0), .ZN(n517) );
  XNOR2_X1 U567 ( .A(n517), .B(KEYINPUT67), .ZN(n634) );
  NAND2_X1 U568 ( .A1(n644), .A2(G51), .ZN(n522) );
  INV_X1 U569 ( .A(G651), .ZN(n526) );
  NOR2_X1 U570 ( .A1(G543), .A2(n526), .ZN(n519) );
  XNOR2_X1 U571 ( .A(KEYINPUT69), .B(KEYINPUT1), .ZN(n518) );
  XNOR2_X1 U572 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U573 ( .A(KEYINPUT68), .B(n520), .ZN(n647) );
  NAND2_X1 U574 ( .A1(G63), .A2(n647), .ZN(n521) );
  NAND2_X1 U575 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U576 ( .A(KEYINPUT6), .B(n523), .ZN(n531) );
  XOR2_X1 U577 ( .A(KEYINPUT4), .B(KEYINPUT75), .Z(n525) );
  NOR2_X1 U578 ( .A1(G651), .A2(G543), .ZN(n643) );
  NAND2_X1 U579 ( .A1(G89), .A2(n643), .ZN(n524) );
  XNOR2_X1 U580 ( .A(n525), .B(n524), .ZN(n528) );
  NOR2_X1 U581 ( .A1(n634), .A2(n526), .ZN(n641) );
  NAND2_X1 U582 ( .A1(n641), .A2(G76), .ZN(n527) );
  NAND2_X1 U583 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U584 ( .A(n529), .B(KEYINPUT5), .Z(n530) );
  NOR2_X1 U585 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U586 ( .A(KEYINPUT76), .B(n532), .Z(n533) );
  XNOR2_X1 U587 ( .A(KEYINPUT7), .B(n533), .ZN(G168) );
  XOR2_X1 U588 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  INV_X1 U589 ( .A(KEYINPUT23), .ZN(n535) );
  INV_X1 U590 ( .A(G2105), .ZN(n536) );
  NAND2_X1 U591 ( .A1(n879), .A2(G101), .ZN(n534) );
  XNOR2_X1 U592 ( .A(n535), .B(n534), .ZN(n538) );
  NOR2_X1 U593 ( .A1(G2104), .A2(n536), .ZN(n883) );
  NAND2_X1 U594 ( .A1(n883), .A2(G125), .ZN(n537) );
  NAND2_X1 U595 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U596 ( .A(KEYINPUT66), .B(n539), .ZN(n544) );
  AND2_X1 U597 ( .A1(G2104), .A2(G2105), .ZN(n885) );
  NAND2_X1 U598 ( .A1(n885), .A2(G113), .ZN(n542) );
  NOR2_X1 U599 ( .A1(G2104), .A2(G2105), .ZN(n540) );
  NAND2_X1 U600 ( .A1(n880), .A2(G137), .ZN(n541) );
  NAND2_X1 U601 ( .A1(n542), .A2(n541), .ZN(n543) );
  INV_X1 U602 ( .A(n677), .ZN(G160) );
  NAND2_X1 U603 ( .A1(G72), .A2(n641), .ZN(n546) );
  NAND2_X1 U604 ( .A1(G60), .A2(n647), .ZN(n545) );
  NAND2_X1 U605 ( .A1(n546), .A2(n545), .ZN(n550) );
  NAND2_X1 U606 ( .A1(G85), .A2(n643), .ZN(n548) );
  NAND2_X1 U607 ( .A1(G47), .A2(n644), .ZN(n547) );
  NAND2_X1 U608 ( .A1(n548), .A2(n547), .ZN(n549) );
  OR2_X1 U609 ( .A1(n550), .A2(n549), .ZN(G290) );
  AND2_X1 U610 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U611 ( .A(G132), .ZN(G219) );
  INV_X1 U612 ( .A(G82), .ZN(G220) );
  INV_X1 U613 ( .A(G57), .ZN(G237) );
  NAND2_X1 U614 ( .A1(G90), .A2(n643), .ZN(n552) );
  NAND2_X1 U615 ( .A1(G77), .A2(n641), .ZN(n551) );
  NAND2_X1 U616 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U617 ( .A(KEYINPUT9), .B(n553), .ZN(n557) );
  NAND2_X1 U618 ( .A1(n647), .A2(G64), .ZN(n555) );
  NAND2_X1 U619 ( .A1(n644), .A2(G52), .ZN(n554) );
  AND2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n556) );
  NAND2_X1 U621 ( .A1(n557), .A2(n556), .ZN(G301) );
  INV_X1 U622 ( .A(G301), .ZN(G171) );
  NAND2_X1 U623 ( .A1(n880), .A2(G138), .ZN(n560) );
  NAND2_X1 U624 ( .A1(G114), .A2(n885), .ZN(n558) );
  XOR2_X1 U625 ( .A(KEYINPUT91), .B(n558), .Z(n559) );
  NAND2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n564) );
  NAND2_X1 U627 ( .A1(G102), .A2(n879), .ZN(n562) );
  NAND2_X1 U628 ( .A1(G126), .A2(n883), .ZN(n561) );
  NAND2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U630 ( .A1(n564), .A2(n563), .ZN(G164) );
  NAND2_X1 U631 ( .A1(G7), .A2(G661), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U633 ( .A(G223), .ZN(n824) );
  NAND2_X1 U634 ( .A1(n824), .A2(G567), .ZN(n566) );
  XNOR2_X1 U635 ( .A(n566), .B(KEYINPUT71), .ZN(n567) );
  XNOR2_X1 U636 ( .A(KEYINPUT11), .B(n567), .ZN(G234) );
  NAND2_X1 U637 ( .A1(G56), .A2(n647), .ZN(n568) );
  XOR2_X1 U638 ( .A(KEYINPUT14), .B(n568), .Z(n576) );
  NAND2_X1 U639 ( .A1(n643), .A2(G81), .ZN(n569) );
  XOR2_X1 U640 ( .A(KEYINPUT12), .B(n569), .Z(n572) );
  NAND2_X1 U641 ( .A1(n641), .A2(G68), .ZN(n570) );
  XOR2_X1 U642 ( .A(n570), .B(KEYINPUT72), .Z(n571) );
  NOR2_X1 U643 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U644 ( .A(KEYINPUT13), .B(n573), .Z(n574) );
  XNOR2_X1 U645 ( .A(n574), .B(KEYINPUT73), .ZN(n575) );
  NOR2_X1 U646 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U647 ( .A1(n644), .A2(G43), .ZN(n577) );
  NAND2_X1 U648 ( .A1(n578), .A2(n577), .ZN(n967) );
  INV_X1 U649 ( .A(G860), .ZN(n829) );
  OR2_X1 U650 ( .A1(n967), .A2(n829), .ZN(G153) );
  NAND2_X1 U651 ( .A1(G79), .A2(n641), .ZN(n580) );
  NAND2_X1 U652 ( .A1(G66), .A2(n647), .ZN(n579) );
  NAND2_X1 U653 ( .A1(n580), .A2(n579), .ZN(n584) );
  NAND2_X1 U654 ( .A1(G92), .A2(n643), .ZN(n582) );
  NAND2_X1 U655 ( .A1(G54), .A2(n644), .ZN(n581) );
  NAND2_X1 U656 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U657 ( .A1(n584), .A2(n583), .ZN(n586) );
  XNOR2_X1 U658 ( .A(KEYINPUT74), .B(KEYINPUT15), .ZN(n585) );
  XNOR2_X1 U659 ( .A(n586), .B(n585), .ZN(n948) );
  NOR2_X1 U660 ( .A1(n948), .A2(G868), .ZN(n588) );
  INV_X1 U661 ( .A(G868), .ZN(n659) );
  NOR2_X1 U662 ( .A1(n659), .A2(G301), .ZN(n587) );
  NOR2_X1 U663 ( .A1(n588), .A2(n587), .ZN(G284) );
  NAND2_X1 U664 ( .A1(G91), .A2(n643), .ZN(n590) );
  NAND2_X1 U665 ( .A1(G78), .A2(n641), .ZN(n589) );
  NAND2_X1 U666 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U667 ( .A(KEYINPUT70), .B(n591), .Z(n595) );
  NAND2_X1 U668 ( .A1(n647), .A2(G65), .ZN(n593) );
  NAND2_X1 U669 ( .A1(n644), .A2(G53), .ZN(n592) );
  AND2_X1 U670 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U671 ( .A1(n595), .A2(n594), .ZN(G299) );
  XNOR2_X1 U672 ( .A(KEYINPUT77), .B(G868), .ZN(n596) );
  NOR2_X1 U673 ( .A1(G286), .A2(n596), .ZN(n598) );
  NOR2_X1 U674 ( .A1(G868), .A2(G299), .ZN(n597) );
  NOR2_X1 U675 ( .A1(n598), .A2(n597), .ZN(G297) );
  NAND2_X1 U676 ( .A1(n829), .A2(G559), .ZN(n599) );
  INV_X1 U677 ( .A(n948), .ZN(n699) );
  NAND2_X1 U678 ( .A1(n599), .A2(n699), .ZN(n600) );
  XNOR2_X1 U679 ( .A(n600), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U680 ( .A1(G868), .A2(n967), .ZN(n603) );
  NAND2_X1 U681 ( .A1(n699), .A2(G868), .ZN(n601) );
  NOR2_X1 U682 ( .A1(G559), .A2(n601), .ZN(n602) );
  NOR2_X1 U683 ( .A1(n603), .A2(n602), .ZN(G282) );
  NAND2_X1 U684 ( .A1(G111), .A2(n885), .ZN(n612) );
  NAND2_X1 U685 ( .A1(G123), .A2(n883), .ZN(n604) );
  XNOR2_X1 U686 ( .A(n604), .B(KEYINPUT78), .ZN(n605) );
  XNOR2_X1 U687 ( .A(n605), .B(KEYINPUT18), .ZN(n607) );
  NAND2_X1 U688 ( .A1(G135), .A2(n880), .ZN(n606) );
  NAND2_X1 U689 ( .A1(n607), .A2(n606), .ZN(n610) );
  NAND2_X1 U690 ( .A1(G99), .A2(n879), .ZN(n608) );
  XNOR2_X1 U691 ( .A(KEYINPUT79), .B(n608), .ZN(n609) );
  NOR2_X1 U692 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U693 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U694 ( .A(n613), .B(KEYINPUT80), .ZN(n922) );
  XOR2_X1 U695 ( .A(n922), .B(G2096), .Z(n615) );
  XNOR2_X1 U696 ( .A(G2100), .B(KEYINPUT81), .ZN(n614) );
  NAND2_X1 U697 ( .A1(n615), .A2(n614), .ZN(G156) );
  NAND2_X1 U698 ( .A1(n641), .A2(G75), .ZN(n618) );
  NAND2_X1 U699 ( .A1(G50), .A2(n644), .ZN(n616) );
  XOR2_X1 U700 ( .A(KEYINPUT87), .B(n616), .Z(n617) );
  NAND2_X1 U701 ( .A1(n618), .A2(n617), .ZN(n622) );
  NAND2_X1 U702 ( .A1(G88), .A2(n643), .ZN(n620) );
  NAND2_X1 U703 ( .A1(G62), .A2(n647), .ZN(n619) );
  NAND2_X1 U704 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U705 ( .A1(n622), .A2(n621), .ZN(G166) );
  NAND2_X1 U706 ( .A1(G48), .A2(n644), .ZN(n623) );
  XNOR2_X1 U707 ( .A(n623), .B(KEYINPUT86), .ZN(n630) );
  NAND2_X1 U708 ( .A1(G86), .A2(n643), .ZN(n625) );
  NAND2_X1 U709 ( .A1(G61), .A2(n647), .ZN(n624) );
  NAND2_X1 U710 ( .A1(n625), .A2(n624), .ZN(n628) );
  NAND2_X1 U711 ( .A1(n641), .A2(G73), .ZN(n626) );
  XOR2_X1 U712 ( .A(KEYINPUT2), .B(n626), .Z(n627) );
  NOR2_X1 U713 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U714 ( .A1(n630), .A2(n629), .ZN(G305) );
  NAND2_X1 U715 ( .A1(G49), .A2(n644), .ZN(n632) );
  NAND2_X1 U716 ( .A1(G74), .A2(G651), .ZN(n631) );
  NAND2_X1 U717 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U718 ( .A1(n647), .A2(n633), .ZN(n637) );
  NAND2_X1 U719 ( .A1(G87), .A2(n634), .ZN(n635) );
  XOR2_X1 U720 ( .A(KEYINPUT85), .B(n635), .Z(n636) );
  NAND2_X1 U721 ( .A1(n637), .A2(n636), .ZN(G288) );
  NAND2_X1 U722 ( .A1(n699), .A2(G559), .ZN(n638) );
  XOR2_X1 U723 ( .A(n967), .B(n638), .Z(n828) );
  XNOR2_X1 U724 ( .A(KEYINPUT88), .B(G305), .ZN(n639) );
  XNOR2_X1 U725 ( .A(n639), .B(G288), .ZN(n640) );
  XOR2_X1 U726 ( .A(n640), .B(KEYINPUT19), .Z(n655) );
  INV_X1 U727 ( .A(G299), .ZN(n952) );
  NAND2_X1 U728 ( .A1(G80), .A2(n641), .ZN(n642) );
  XNOR2_X1 U729 ( .A(n642), .B(KEYINPUT82), .ZN(n652) );
  NAND2_X1 U730 ( .A1(G93), .A2(n643), .ZN(n646) );
  NAND2_X1 U731 ( .A1(G55), .A2(n644), .ZN(n645) );
  NAND2_X1 U732 ( .A1(n646), .A2(n645), .ZN(n650) );
  NAND2_X1 U733 ( .A1(G67), .A2(n647), .ZN(n648) );
  XNOR2_X1 U734 ( .A(KEYINPUT83), .B(n648), .ZN(n649) );
  NOR2_X1 U735 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U736 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U737 ( .A(KEYINPUT84), .B(n653), .ZN(n830) );
  XNOR2_X1 U738 ( .A(n952), .B(n830), .ZN(n654) );
  XNOR2_X1 U739 ( .A(n655), .B(n654), .ZN(n656) );
  XOR2_X1 U740 ( .A(G166), .B(n656), .Z(n657) );
  XNOR2_X1 U741 ( .A(G290), .B(n657), .ZN(n900) );
  XNOR2_X1 U742 ( .A(n828), .B(n900), .ZN(n658) );
  NAND2_X1 U743 ( .A1(n658), .A2(G868), .ZN(n661) );
  NAND2_X1 U744 ( .A1(n659), .A2(n830), .ZN(n660) );
  NAND2_X1 U745 ( .A1(n661), .A2(n660), .ZN(G295) );
  XOR2_X1 U746 ( .A(KEYINPUT89), .B(KEYINPUT21), .Z(n665) );
  NAND2_X1 U747 ( .A1(G2084), .A2(G2078), .ZN(n662) );
  XOR2_X1 U748 ( .A(KEYINPUT20), .B(n662), .Z(n663) );
  NAND2_X1 U749 ( .A1(n663), .A2(G2090), .ZN(n664) );
  XNOR2_X1 U750 ( .A(n665), .B(n664), .ZN(n666) );
  NAND2_X1 U751 ( .A1(G2072), .A2(n666), .ZN(G158) );
  XNOR2_X1 U752 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U753 ( .A1(G120), .A2(G69), .ZN(n667) );
  NOR2_X1 U754 ( .A1(G237), .A2(n667), .ZN(n668) );
  XNOR2_X1 U755 ( .A(KEYINPUT90), .B(n668), .ZN(n669) );
  NAND2_X1 U756 ( .A1(n669), .A2(G108), .ZN(n833) );
  NAND2_X1 U757 ( .A1(n833), .A2(G567), .ZN(n674) );
  NOR2_X1 U758 ( .A1(G220), .A2(G219), .ZN(n670) );
  XOR2_X1 U759 ( .A(KEYINPUT22), .B(n670), .Z(n671) );
  NOR2_X1 U760 ( .A1(G218), .A2(n671), .ZN(n672) );
  NAND2_X1 U761 ( .A1(G96), .A2(n672), .ZN(n832) );
  NAND2_X1 U762 ( .A1(n832), .A2(G2106), .ZN(n673) );
  NAND2_X1 U763 ( .A1(n674), .A2(n673), .ZN(n835) );
  NAND2_X1 U764 ( .A1(G661), .A2(G483), .ZN(n675) );
  NOR2_X1 U765 ( .A1(n835), .A2(n675), .ZN(n827) );
  NAND2_X1 U766 ( .A1(n827), .A2(G36), .ZN(G176) );
  XOR2_X1 U767 ( .A(KEYINPUT92), .B(G166), .Z(G303) );
  INV_X1 U768 ( .A(KEYINPUT94), .ZN(n679) );
  NOR2_X1 U769 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U770 ( .A(n679), .B(n678), .ZN(n769) );
  NOR2_X1 U771 ( .A1(G164), .A2(G1384), .ZN(n680) );
  XOR2_X1 U772 ( .A(KEYINPUT64), .B(n680), .Z(n770) );
  INV_X1 U773 ( .A(n713), .ZN(n725) );
  NAND2_X1 U774 ( .A1(G8), .A2(n725), .ZN(n765) );
  NOR2_X1 U775 ( .A1(G1976), .A2(G288), .ZN(n744) );
  NAND2_X1 U776 ( .A1(n744), .A2(KEYINPUT33), .ZN(n681) );
  NOR2_X1 U777 ( .A1(n765), .A2(n681), .ZN(n751) );
  NOR2_X1 U778 ( .A1(n713), .A2(G1961), .ZN(n682) );
  XNOR2_X1 U779 ( .A(n682), .B(KEYINPUT100), .ZN(n684) );
  XOR2_X1 U780 ( .A(KEYINPUT25), .B(G2078), .Z(n978) );
  NOR2_X1 U781 ( .A1(n725), .A2(n978), .ZN(n683) );
  NOR2_X1 U782 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U783 ( .A(KEYINPUT101), .B(n685), .ZN(n712) );
  NAND2_X1 U784 ( .A1(n712), .A2(G171), .ZN(n711) );
  NAND2_X1 U785 ( .A1(n713), .A2(G2072), .ZN(n686) );
  XNOR2_X1 U786 ( .A(n686), .B(KEYINPUT27), .ZN(n688) );
  INV_X1 U787 ( .A(G1956), .ZN(n1001) );
  NOR2_X1 U788 ( .A1(n1001), .A2(n713), .ZN(n687) );
  NOR2_X1 U789 ( .A1(n688), .A2(n687), .ZN(n705) );
  NAND2_X1 U790 ( .A1(n705), .A2(n952), .ZN(n704) );
  AND2_X1 U791 ( .A1(n713), .A2(G1996), .ZN(n690) );
  NAND2_X1 U792 ( .A1(n725), .A2(G1341), .ZN(n691) );
  NAND2_X1 U793 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U794 ( .A1(n967), .A2(n693), .ZN(n694) );
  XNOR2_X1 U795 ( .A(n694), .B(KEYINPUT65), .ZN(n698) );
  INV_X1 U796 ( .A(G2067), .ZN(n972) );
  NOR2_X1 U797 ( .A1(n725), .A2(n972), .ZN(n696) );
  INV_X1 U798 ( .A(G1348), .ZN(n1004) );
  NOR2_X1 U799 ( .A1(n713), .A2(n1004), .ZN(n695) );
  NOR2_X1 U800 ( .A1(n696), .A2(n695), .ZN(n700) );
  NAND2_X1 U801 ( .A1(n699), .A2(n700), .ZN(n697) );
  NAND2_X1 U802 ( .A1(n698), .A2(n697), .ZN(n702) );
  OR2_X1 U803 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U804 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U805 ( .A1(n704), .A2(n703), .ZN(n708) );
  NOR2_X1 U806 ( .A1(n705), .A2(n952), .ZN(n706) );
  XOR2_X1 U807 ( .A(n706), .B(KEYINPUT28), .Z(n707) );
  NAND2_X1 U808 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U809 ( .A(KEYINPUT29), .B(n709), .Z(n710) );
  NAND2_X1 U810 ( .A1(n711), .A2(n710), .ZN(n724) );
  NOR2_X1 U811 ( .A1(G171), .A2(n712), .ZN(n719) );
  NOR2_X1 U812 ( .A1(G1966), .A2(n765), .ZN(n736) );
  INV_X1 U813 ( .A(G2084), .ZN(n714) );
  NAND2_X1 U814 ( .A1(n714), .A2(n713), .ZN(n734) );
  NAND2_X1 U815 ( .A1(G8), .A2(n734), .ZN(n715) );
  OR2_X1 U816 ( .A1(n736), .A2(n715), .ZN(n716) );
  NOR2_X1 U817 ( .A1(n717), .A2(G168), .ZN(n718) );
  NOR2_X1 U818 ( .A1(n719), .A2(n718), .ZN(n722) );
  NAND2_X1 U819 ( .A1(n724), .A2(n723), .ZN(n737) );
  NAND2_X1 U820 ( .A1(n737), .A2(G286), .ZN(n731) );
  NOR2_X1 U821 ( .A1(G2090), .A2(n725), .ZN(n728) );
  NOR2_X1 U822 ( .A1(G1971), .A2(n765), .ZN(n726) );
  XOR2_X1 U823 ( .A(KEYINPUT103), .B(n726), .Z(n727) );
  NOR2_X1 U824 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U825 ( .A1(n729), .A2(G303), .ZN(n730) );
  NAND2_X1 U826 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U827 ( .A1(n732), .A2(G8), .ZN(n733) );
  INV_X1 U828 ( .A(n734), .ZN(n735) );
  NAND2_X1 U829 ( .A1(G8), .A2(n735), .ZN(n740) );
  INV_X1 U830 ( .A(n737), .ZN(n738) );
  NOR2_X1 U831 ( .A1(n736), .A2(n738), .ZN(n739) );
  NAND2_X1 U832 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U833 ( .A1(n742), .A2(n741), .ZN(n761) );
  NOR2_X1 U834 ( .A1(G303), .A2(G1971), .ZN(n743) );
  NOR2_X1 U835 ( .A1(n744), .A2(n743), .ZN(n947) );
  INV_X1 U836 ( .A(KEYINPUT33), .ZN(n745) );
  AND2_X1 U837 ( .A1(n947), .A2(n745), .ZN(n746) );
  NAND2_X1 U838 ( .A1(n761), .A2(n746), .ZN(n749) );
  NAND2_X1 U839 ( .A1(G1976), .A2(G288), .ZN(n946) );
  INV_X1 U840 ( .A(n946), .ZN(n747) );
  OR2_X1 U841 ( .A1(KEYINPUT33), .A2(n516), .ZN(n748) );
  NAND2_X1 U842 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U843 ( .A1(n751), .A2(n750), .ZN(n753) );
  XOR2_X1 U844 ( .A(G1981), .B(KEYINPUT104), .Z(n752) );
  XNOR2_X1 U845 ( .A(G305), .B(n752), .ZN(n961) );
  NAND2_X1 U846 ( .A1(n753), .A2(n961), .ZN(n754) );
  XNOR2_X1 U847 ( .A(n754), .B(KEYINPUT105), .ZN(n758) );
  NOR2_X1 U848 ( .A1(G1981), .A2(G305), .ZN(n755) );
  XOR2_X1 U849 ( .A(n755), .B(KEYINPUT24), .Z(n756) );
  NOR2_X1 U850 ( .A1(n765), .A2(n756), .ZN(n757) );
  NOR2_X1 U851 ( .A1(G303), .A2(G2090), .ZN(n759) );
  XNOR2_X1 U852 ( .A(n759), .B(KEYINPUT106), .ZN(n760) );
  NAND2_X1 U853 ( .A1(n760), .A2(G8), .ZN(n762) );
  NAND2_X1 U854 ( .A1(n762), .A2(n761), .ZN(n763) );
  XOR2_X1 U855 ( .A(KEYINPUT107), .B(n763), .Z(n764) );
  NAND2_X1 U856 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U857 ( .A1(n767), .A2(n766), .ZN(n806) );
  XOR2_X1 U858 ( .A(KEYINPUT93), .B(G1986), .Z(n768) );
  XNOR2_X1 U859 ( .A(G290), .B(n768), .ZN(n956) );
  INV_X1 U860 ( .A(n769), .ZN(n771) );
  NAND2_X1 U861 ( .A1(n771), .A2(n770), .ZN(n772) );
  XOR2_X1 U862 ( .A(n772), .B(KEYINPUT95), .Z(n801) );
  INV_X1 U863 ( .A(n801), .ZN(n818) );
  NAND2_X1 U864 ( .A1(n956), .A2(n818), .ZN(n804) );
  XNOR2_X1 U865 ( .A(G2067), .B(KEYINPUT37), .ZN(n815) );
  NAND2_X1 U866 ( .A1(G104), .A2(n879), .ZN(n774) );
  NAND2_X1 U867 ( .A1(G140), .A2(n880), .ZN(n773) );
  NAND2_X1 U868 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U869 ( .A(KEYINPUT34), .B(n775), .ZN(n781) );
  NAND2_X1 U870 ( .A1(G128), .A2(n883), .ZN(n777) );
  NAND2_X1 U871 ( .A1(G116), .A2(n885), .ZN(n776) );
  NAND2_X1 U872 ( .A1(n777), .A2(n776), .ZN(n778) );
  XOR2_X1 U873 ( .A(KEYINPUT35), .B(n778), .Z(n779) );
  XNOR2_X1 U874 ( .A(KEYINPUT96), .B(n779), .ZN(n780) );
  NOR2_X1 U875 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U876 ( .A(KEYINPUT36), .B(n782), .ZN(n891) );
  NOR2_X1 U877 ( .A1(n815), .A2(n891), .ZN(n920) );
  NAND2_X1 U878 ( .A1(n818), .A2(n920), .ZN(n813) );
  NAND2_X1 U879 ( .A1(n883), .A2(G119), .ZN(n783) );
  XOR2_X1 U880 ( .A(KEYINPUT97), .B(n783), .Z(n785) );
  NAND2_X1 U881 ( .A1(n885), .A2(G107), .ZN(n784) );
  NAND2_X1 U882 ( .A1(n785), .A2(n784), .ZN(n786) );
  XOR2_X1 U883 ( .A(KEYINPUT98), .B(n786), .Z(n790) );
  NAND2_X1 U884 ( .A1(n879), .A2(G95), .ZN(n788) );
  NAND2_X1 U885 ( .A1(G131), .A2(n880), .ZN(n787) );
  AND2_X1 U886 ( .A1(n788), .A2(n787), .ZN(n789) );
  NAND2_X1 U887 ( .A1(n790), .A2(n789), .ZN(n894) );
  AND2_X1 U888 ( .A1(n894), .A2(G1991), .ZN(n800) );
  NAND2_X1 U889 ( .A1(n885), .A2(G117), .ZN(n797) );
  NAND2_X1 U890 ( .A1(G129), .A2(n883), .ZN(n792) );
  NAND2_X1 U891 ( .A1(G141), .A2(n880), .ZN(n791) );
  NAND2_X1 U892 ( .A1(n792), .A2(n791), .ZN(n795) );
  NAND2_X1 U893 ( .A1(n879), .A2(G105), .ZN(n793) );
  XOR2_X1 U894 ( .A(KEYINPUT38), .B(n793), .Z(n794) );
  NOR2_X1 U895 ( .A1(n795), .A2(n794), .ZN(n796) );
  NAND2_X1 U896 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U897 ( .A(KEYINPUT99), .B(n798), .ZN(n874) );
  INV_X1 U898 ( .A(G1996), .ZN(n807) );
  NOR2_X1 U899 ( .A1(n874), .A2(n807), .ZN(n799) );
  NOR2_X1 U900 ( .A1(n800), .A2(n799), .ZN(n927) );
  NOR2_X1 U901 ( .A1(n927), .A2(n801), .ZN(n810) );
  INV_X1 U902 ( .A(n810), .ZN(n802) );
  AND2_X1 U903 ( .A1(n813), .A2(n802), .ZN(n803) );
  AND2_X1 U904 ( .A1(n804), .A2(n803), .ZN(n805) );
  NAND2_X1 U905 ( .A1(n806), .A2(n805), .ZN(n821) );
  AND2_X1 U906 ( .A1(n807), .A2(n874), .ZN(n930) );
  NOR2_X1 U907 ( .A1(G1986), .A2(G290), .ZN(n808) );
  NOR2_X1 U908 ( .A1(G1991), .A2(n894), .ZN(n919) );
  NOR2_X1 U909 ( .A1(n808), .A2(n919), .ZN(n809) );
  NOR2_X1 U910 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U911 ( .A1(n930), .A2(n811), .ZN(n812) );
  XNOR2_X1 U912 ( .A(KEYINPUT39), .B(n812), .ZN(n814) );
  NAND2_X1 U913 ( .A1(n814), .A2(n813), .ZN(n817) );
  NAND2_X1 U914 ( .A1(n891), .A2(n815), .ZN(n816) );
  XNOR2_X1 U915 ( .A(n816), .B(KEYINPUT108), .ZN(n941) );
  NAND2_X1 U916 ( .A1(n817), .A2(n941), .ZN(n819) );
  NAND2_X1 U917 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U918 ( .A1(n821), .A2(n820), .ZN(n823) );
  XOR2_X1 U919 ( .A(KEYINPUT109), .B(KEYINPUT40), .Z(n822) );
  XNOR2_X1 U920 ( .A(n823), .B(n822), .ZN(G329) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n824), .ZN(G217) );
  AND2_X1 U922 ( .A1(G15), .A2(G2), .ZN(n825) );
  NAND2_X1 U923 ( .A1(G661), .A2(n825), .ZN(G259) );
  NAND2_X1 U924 ( .A1(G3), .A2(G1), .ZN(n826) );
  NAND2_X1 U925 ( .A1(n827), .A2(n826), .ZN(G188) );
  XOR2_X1 U926 ( .A(G96), .B(KEYINPUT110), .Z(G221) );
  NAND2_X1 U928 ( .A1(n829), .A2(n828), .ZN(n831) );
  XNOR2_X1 U929 ( .A(n831), .B(n830), .ZN(G145) );
  INV_X1 U930 ( .A(G120), .ZN(G236) );
  INV_X1 U931 ( .A(G108), .ZN(G238) );
  INV_X1 U932 ( .A(G69), .ZN(G235) );
  NOR2_X1 U933 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U934 ( .A(n834), .B(KEYINPUT111), .ZN(G261) );
  INV_X1 U935 ( .A(G261), .ZN(G325) );
  INV_X1 U936 ( .A(n835), .ZN(G319) );
  XOR2_X1 U937 ( .A(KEYINPUT112), .B(KEYINPUT114), .Z(n837) );
  XNOR2_X1 U938 ( .A(G2678), .B(G2096), .ZN(n836) );
  XNOR2_X1 U939 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U940 ( .A(n838), .B(KEYINPUT113), .Z(n840) );
  XNOR2_X1 U941 ( .A(G2078), .B(G2072), .ZN(n839) );
  XNOR2_X1 U942 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U943 ( .A(G2100), .B(G2090), .Z(n842) );
  XNOR2_X1 U944 ( .A(G2084), .B(G2067), .ZN(n841) );
  XNOR2_X1 U945 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U946 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U947 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n845) );
  XNOR2_X1 U948 ( .A(n846), .B(n845), .ZN(G227) );
  XOR2_X1 U949 ( .A(G1981), .B(G1956), .Z(n848) );
  XNOR2_X1 U950 ( .A(G1966), .B(G1961), .ZN(n847) );
  XNOR2_X1 U951 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U952 ( .A(n849), .B(KEYINPUT41), .Z(n851) );
  XNOR2_X1 U953 ( .A(G1996), .B(G1991), .ZN(n850) );
  XNOR2_X1 U954 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U955 ( .A(G2474), .B(G1986), .Z(n853) );
  XNOR2_X1 U956 ( .A(G1971), .B(G1976), .ZN(n852) );
  XNOR2_X1 U957 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U958 ( .A(n855), .B(n854), .ZN(G229) );
  NAND2_X1 U959 ( .A1(G124), .A2(n883), .ZN(n856) );
  XOR2_X1 U960 ( .A(KEYINPUT44), .B(n856), .Z(n857) );
  XNOR2_X1 U961 ( .A(n857), .B(KEYINPUT115), .ZN(n859) );
  NAND2_X1 U962 ( .A1(G112), .A2(n885), .ZN(n858) );
  NAND2_X1 U963 ( .A1(n859), .A2(n858), .ZN(n863) );
  NAND2_X1 U964 ( .A1(G100), .A2(n879), .ZN(n861) );
  NAND2_X1 U965 ( .A1(G136), .A2(n880), .ZN(n860) );
  NAND2_X1 U966 ( .A1(n861), .A2(n860), .ZN(n862) );
  NOR2_X1 U967 ( .A1(n863), .A2(n862), .ZN(G162) );
  NAND2_X1 U968 ( .A1(G130), .A2(n883), .ZN(n865) );
  NAND2_X1 U969 ( .A1(G118), .A2(n885), .ZN(n864) );
  NAND2_X1 U970 ( .A1(n865), .A2(n864), .ZN(n870) );
  NAND2_X1 U971 ( .A1(G106), .A2(n879), .ZN(n867) );
  NAND2_X1 U972 ( .A1(G142), .A2(n880), .ZN(n866) );
  NAND2_X1 U973 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U974 ( .A(KEYINPUT45), .B(n868), .Z(n869) );
  NOR2_X1 U975 ( .A1(n870), .A2(n869), .ZN(n878) );
  XOR2_X1 U976 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n872) );
  XNOR2_X1 U977 ( .A(G164), .B(KEYINPUT116), .ZN(n871) );
  XNOR2_X1 U978 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U979 ( .A(n873), .B(G162), .Z(n876) );
  XNOR2_X1 U980 ( .A(n874), .B(n922), .ZN(n875) );
  XNOR2_X1 U981 ( .A(n876), .B(n875), .ZN(n877) );
  XNOR2_X1 U982 ( .A(n878), .B(n877), .ZN(n893) );
  NAND2_X1 U983 ( .A1(G103), .A2(n879), .ZN(n882) );
  NAND2_X1 U984 ( .A1(G139), .A2(n880), .ZN(n881) );
  NAND2_X1 U985 ( .A1(n882), .A2(n881), .ZN(n890) );
  NAND2_X1 U986 ( .A1(n883), .A2(G127), .ZN(n884) );
  XOR2_X1 U987 ( .A(KEYINPUT117), .B(n884), .Z(n887) );
  NAND2_X1 U988 ( .A1(n885), .A2(G115), .ZN(n886) );
  NAND2_X1 U989 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U990 ( .A(KEYINPUT47), .B(n888), .Z(n889) );
  NOR2_X1 U991 ( .A1(n890), .A2(n889), .ZN(n923) );
  XNOR2_X1 U992 ( .A(n891), .B(n923), .ZN(n892) );
  XNOR2_X1 U993 ( .A(n893), .B(n892), .ZN(n896) );
  XNOR2_X1 U994 ( .A(n894), .B(G160), .ZN(n895) );
  XNOR2_X1 U995 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U996 ( .A1(G37), .A2(n897), .ZN(G395) );
  XNOR2_X1 U997 ( .A(G286), .B(KEYINPUT118), .ZN(n899) );
  XNOR2_X1 U998 ( .A(G171), .B(n948), .ZN(n898) );
  XNOR2_X1 U999 ( .A(n899), .B(n898), .ZN(n902) );
  XOR2_X1 U1000 ( .A(n967), .B(n900), .Z(n901) );
  XNOR2_X1 U1001 ( .A(n902), .B(n901), .ZN(n903) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n903), .ZN(G397) );
  XOR2_X1 U1003 ( .A(G2451), .B(G2430), .Z(n905) );
  XNOR2_X1 U1004 ( .A(G2438), .B(G2443), .ZN(n904) );
  XNOR2_X1 U1005 ( .A(n905), .B(n904), .ZN(n911) );
  XOR2_X1 U1006 ( .A(G2435), .B(G2454), .Z(n907) );
  XNOR2_X1 U1007 ( .A(G1348), .B(G1341), .ZN(n906) );
  XNOR2_X1 U1008 ( .A(n907), .B(n906), .ZN(n909) );
  XOR2_X1 U1009 ( .A(G2446), .B(G2427), .Z(n908) );
  XNOR2_X1 U1010 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1011 ( .A(n911), .B(n910), .Z(n912) );
  NAND2_X1 U1012 ( .A1(G14), .A2(n912), .ZN(n918) );
  NAND2_X1 U1013 ( .A1(G319), .A2(n918), .ZN(n915) );
  NOR2_X1 U1014 ( .A1(G227), .A2(G229), .ZN(n913) );
  XNOR2_X1 U1015 ( .A(KEYINPUT49), .B(n913), .ZN(n914) );
  NOR2_X1 U1016 ( .A1(n915), .A2(n914), .ZN(n917) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n916) );
  NAND2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(n918), .ZN(G401) );
  NOR2_X1 U1021 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(n939) );
  XOR2_X1 U1023 ( .A(G2072), .B(n923), .Z(n925) );
  XOR2_X1 U1024 ( .A(G164), .B(G2078), .Z(n924) );
  NOR2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1026 ( .A(KEYINPUT50), .B(n926), .ZN(n937) );
  XNOR2_X1 U1027 ( .A(G160), .B(G2084), .ZN(n928) );
  NAND2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n935) );
  XOR2_X1 U1029 ( .A(G2090), .B(G162), .Z(n929) );
  NOR2_X1 U1030 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1031 ( .A(KEYINPUT51), .B(n931), .Z(n933) );
  XNOR2_X1 U1032 ( .A(KEYINPUT120), .B(KEYINPUT119), .ZN(n932) );
  XNOR2_X1 U1033 ( .A(n933), .B(n932), .ZN(n934) );
  NOR2_X1 U1034 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1035 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1037 ( .A1(n941), .A2(n940), .ZN(n942) );
  XOR2_X1 U1038 ( .A(KEYINPUT52), .B(n942), .Z(n944) );
  INV_X1 U1039 ( .A(KEYINPUT55), .ZN(n943) );
  NAND2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1041 ( .A1(n945), .A2(G29), .ZN(n998) );
  NAND2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n950) );
  XNOR2_X1 U1043 ( .A(G1348), .B(n948), .ZN(n949) );
  NOR2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n966) );
  XNOR2_X1 U1045 ( .A(G1961), .B(G171), .ZN(n951) );
  XNOR2_X1 U1046 ( .A(n951), .B(KEYINPUT124), .ZN(n958) );
  XNOR2_X1 U1047 ( .A(n952), .B(G1956), .ZN(n954) );
  NAND2_X1 U1048 ( .A1(G1971), .A2(G303), .ZN(n953) );
  NAND2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1051 ( .A1(n958), .A2(n957), .ZN(n964) );
  XOR2_X1 U1052 ( .A(G1966), .B(KEYINPUT123), .Z(n959) );
  XNOR2_X1 U1053 ( .A(G168), .B(n959), .ZN(n960) );
  NAND2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1055 ( .A(KEYINPUT57), .B(n962), .Z(n963) );
  NOR2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1057 ( .A1(n966), .A2(n965), .ZN(n969) );
  XNOR2_X1 U1058 ( .A(G1341), .B(n967), .ZN(n968) );
  NOR2_X1 U1059 ( .A1(n969), .A2(n968), .ZN(n971) );
  XOR2_X1 U1060 ( .A(G16), .B(KEYINPUT56), .Z(n970) );
  NOR2_X1 U1061 ( .A1(n971), .A2(n970), .ZN(n996) );
  XOR2_X1 U1062 ( .A(G1991), .B(G25), .Z(n974) );
  XNOR2_X1 U1063 ( .A(n972), .B(G26), .ZN(n973) );
  NAND2_X1 U1064 ( .A1(n974), .A2(n973), .ZN(n976) );
  XNOR2_X1 U1065 ( .A(G32), .B(G1996), .ZN(n975) );
  NOR2_X1 U1066 ( .A1(n976), .A2(n975), .ZN(n983) );
  XOR2_X1 U1067 ( .A(G2072), .B(G33), .Z(n977) );
  NAND2_X1 U1068 ( .A1(n977), .A2(G28), .ZN(n981) );
  XOR2_X1 U1069 ( .A(G27), .B(n978), .Z(n979) );
  XNOR2_X1 U1070 ( .A(KEYINPUT121), .B(n979), .ZN(n980) );
  NOR2_X1 U1071 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1072 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1073 ( .A(n984), .B(KEYINPUT53), .ZN(n987) );
  XOR2_X1 U1074 ( .A(G2084), .B(KEYINPUT54), .Z(n985) );
  XNOR2_X1 U1075 ( .A(G34), .B(n985), .ZN(n986) );
  NAND2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n989) );
  XNOR2_X1 U1077 ( .A(G35), .B(G2090), .ZN(n988) );
  NOR2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1079 ( .A(n990), .B(KEYINPUT55), .ZN(n992) );
  INV_X1 U1080 ( .A(G29), .ZN(n991) );
  NAND2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1082 ( .A1(G11), .A2(n993), .ZN(n994) );
  XNOR2_X1 U1083 ( .A(KEYINPUT122), .B(n994), .ZN(n995) );
  NOR2_X1 U1084 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1085 ( .A1(n998), .A2(n997), .ZN(n1026) );
  XNOR2_X1 U1086 ( .A(G1966), .B(G21), .ZN(n1000) );
  XNOR2_X1 U1087 ( .A(G5), .B(G1961), .ZN(n999) );
  NOR2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1013) );
  XOR2_X1 U1089 ( .A(G1341), .B(G19), .Z(n1003) );
  XNOR2_X1 U1090 ( .A(n1001), .B(G20), .ZN(n1002) );
  NAND2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1010) );
  XOR2_X1 U1092 ( .A(G1981), .B(G6), .Z(n1008) );
  XNOR2_X1 U1093 ( .A(KEYINPUT125), .B(G4), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(n1005), .B(n1004), .ZN(n1006) );
  XNOR2_X1 U1095 ( .A(n1006), .B(KEYINPUT59), .ZN(n1007) );
  NAND2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1098 ( .A(n1011), .B(KEYINPUT60), .ZN(n1012) );
  NAND2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1021) );
  XOR2_X1 U1100 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n1019) );
  XOR2_X1 U1101 ( .A(G1986), .B(G24), .Z(n1017) );
  XNOR2_X1 U1102 ( .A(G1971), .B(G22), .ZN(n1015) );
  XNOR2_X1 U1103 ( .A(G23), .B(G1976), .ZN(n1014) );
  NOR2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1106 ( .A(n1019), .B(n1018), .Z(n1020) );
  NOR2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1108 ( .A(KEYINPUT61), .B(n1022), .Z(n1023) );
  NOR2_X1 U1109 ( .A1(G16), .A2(n1023), .ZN(n1024) );
  XOR2_X1 U1110 ( .A(KEYINPUT127), .B(n1024), .Z(n1025) );
  NOR2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1112 ( .A(n1027), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

