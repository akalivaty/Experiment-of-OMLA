//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 1 1 0 0 1 1 0 0 1 1 1 1 0 0 0 1 0 0 1 0 0 0 0 0 0 0 0 0 0 1 0 1 1 1 1 0 1 1 1 0 1 0 1 1 1 0 1 1 0 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n876, new_n877,
    new_n879, new_n880, new_n881, new_n882, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n975, new_n976, new_n977, new_n978, new_n979;
  INV_X1    g000(.A(G120gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G113gat), .ZN(new_n203));
  INV_X1    g002(.A(G113gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G120gat), .ZN(new_n205));
  AOI21_X1  g004(.A(KEYINPUT1), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G127gat), .B(G134gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(KEYINPUT65), .A2(G127gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(KEYINPUT65), .A2(G127gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n210), .A2(G134gat), .A3(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(G127gat), .A2(G134gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  AND3_X1   g013(.A1(new_n212), .A2(KEYINPUT66), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(KEYINPUT66), .B1(new_n212), .B2(new_n214), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n206), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n209), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT27), .B(G183gat), .ZN(new_n220));
  INV_X1    g019(.A(G190gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT28), .ZN(new_n223));
  NAND2_X1  g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT64), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n230));
  OR3_X1    g029(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT28), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n220), .A2(new_n233), .A3(new_n221), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n223), .A2(new_n224), .A3(new_n232), .A4(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT23), .ZN(new_n236));
  INV_X1    g035(.A(G169gat), .ZN(new_n237));
  INV_X1    g036(.A(G176gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(G183gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(new_n221), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n243), .A2(KEYINPUT24), .A3(new_n224), .ZN(new_n244));
  OR2_X1    g043(.A1(new_n224), .A2(KEYINPUT24), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n241), .A2(new_n244), .A3(new_n229), .A4(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT25), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n224), .A2(KEYINPUT24), .ZN(new_n249));
  AND2_X1   g048(.A1(G183gat), .A2(G190gat), .ZN(new_n250));
  NOR2_X1   g049(.A1(G183gat), .A2(G190gat), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n249), .B1(new_n252), .B2(KEYINPUT24), .ZN(new_n253));
  AOI22_X1  g052(.A1(new_n240), .A2(new_n239), .B1(new_n227), .B2(new_n228), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT25), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n235), .B1(new_n248), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n219), .A2(new_n256), .ZN(new_n257));
  AND2_X1   g056(.A1(G227gat), .A2(G233gat), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n259));
  AND2_X1   g058(.A1(KEYINPUT65), .A2(G127gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(KEYINPUT65), .A2(G127gat), .ZN(new_n261));
  INV_X1    g060(.A(G134gat), .ZN(new_n262));
  NOR3_X1   g061(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n259), .B1(new_n263), .B2(new_n213), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n212), .A2(KEYINPUT66), .A3(new_n214), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n264), .A2(new_n218), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(new_n208), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n246), .A2(new_n247), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n253), .A2(new_n254), .A3(KEYINPUT25), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n267), .A2(new_n270), .A3(new_n235), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n257), .A2(new_n258), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT67), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n257), .A2(new_n271), .A3(KEYINPUT67), .A4(new_n258), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT32), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT68), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G15gat), .B(G43gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(G71gat), .ZN(new_n281));
  INV_X1    g080(.A(G99gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT33), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n284), .B1(new_n276), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n276), .A2(KEYINPUT68), .A3(KEYINPUT32), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n279), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(KEYINPUT33), .B1(new_n283), .B2(KEYINPUT69), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n289), .B1(KEYINPUT69), .B2(new_n283), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n277), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n258), .B1(new_n257), .B2(new_n271), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT70), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT34), .ZN(new_n295));
  AND3_X1   g094(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n294), .B1(new_n293), .B2(new_n295), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n293), .A2(new_n295), .ZN(new_n298));
  NOR3_X1   g097(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n288), .A2(new_n292), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n299), .B1(new_n288), .B2(new_n292), .ZN(new_n301));
  XNOR2_X1  g100(.A(G78gat), .B(G106gat), .ZN(new_n302));
  XOR2_X1   g101(.A(new_n302), .B(G22gat), .Z(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G141gat), .ZN(new_n305));
  INV_X1    g104(.A(G148gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(G141gat), .A2(G148gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT2), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n310), .B1(G155gat), .B2(G162gat), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT75), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G155gat), .B(G162gat), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(G155gat), .ZN(new_n316));
  INV_X1    g115(.A(G162gat), .ZN(new_n317));
  OAI21_X1  g116(.A(KEYINPUT2), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n318), .A2(new_n307), .A3(new_n308), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n319), .A2(KEYINPUT75), .A3(new_n313), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT29), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT72), .ZN(new_n323));
  OR2_X1    g122(.A1(KEYINPUT71), .A2(G204gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(KEYINPUT71), .A2(G204gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G197gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT22), .ZN(new_n329));
  INV_X1    g128(.A(G211gat), .ZN(new_n330));
  INV_X1    g129(.A(G218gat), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n324), .A2(G197gat), .A3(new_n325), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n328), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  XOR2_X1   g133(.A(G211gat), .B(G218gat), .Z(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n335), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n337), .A2(new_n328), .A3(new_n332), .A4(new_n333), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n323), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT72), .B1(new_n334), .B2(new_n335), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n322), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n321), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n336), .A2(new_n338), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT72), .ZN(new_n345));
  INV_X1    g144(.A(new_n340), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT29), .B1(new_n321), .B2(new_n342), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G228gat), .A2(G233gat), .ZN(new_n350));
  NOR3_X1   g149(.A1(new_n343), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(KEYINPUT31), .B(G50gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n350), .B(KEYINPUT79), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  OR3_X1    g153(.A1(new_n348), .A2(new_n339), .A3(new_n340), .ZN(new_n355));
  INV_X1    g154(.A(new_n321), .ZN(new_n356));
  AOI21_X1  g155(.A(KEYINPUT29), .B1(new_n336), .B2(new_n338), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n356), .B1(new_n357), .B2(KEYINPUT3), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n354), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  NOR3_X1   g158(.A1(new_n351), .A2(new_n352), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n352), .ZN(new_n361));
  INV_X1    g160(.A(new_n350), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT3), .B1(new_n347), .B2(new_n322), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n355), .B(new_n362), .C1(new_n363), .C2(new_n321), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n355), .A2(new_n358), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n353), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n361), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n304), .B1(new_n360), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n352), .B1(new_n351), .B2(new_n359), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n364), .A2(new_n366), .A3(new_n361), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n369), .A2(new_n303), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  NOR3_X1   g171(.A1(new_n300), .A2(new_n301), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n267), .A2(new_n356), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n321), .A2(new_n266), .A3(new_n208), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n374), .A2(KEYINPUT76), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(G225gat), .A2(G233gat), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT76), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n267), .A2(new_n356), .A3(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n376), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT4), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n375), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n375), .A2(new_n378), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n321), .A2(new_n342), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n315), .A2(KEYINPUT3), .A3(new_n320), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n385), .A2(new_n267), .A3(new_n386), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n321), .A2(new_n266), .A3(KEYINPUT4), .A4(new_n208), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n383), .A2(new_n384), .A3(new_n387), .A4(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n381), .A2(KEYINPUT5), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n383), .A2(new_n388), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT77), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n375), .A2(KEYINPUT77), .A3(KEYINPUT4), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n394), .A2(new_n387), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n378), .A2(KEYINPUT5), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n393), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(KEYINPUT0), .B(G57gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n398), .B(G85gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(G1gat), .B(G29gat), .ZN(new_n400));
  XOR2_X1   g199(.A(new_n399), .B(new_n400), .Z(new_n401));
  NAND3_X1  g200(.A1(new_n390), .A2(new_n397), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT78), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n390), .A2(new_n397), .ZN(new_n404));
  INV_X1    g203(.A(new_n401), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT6), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT78), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n390), .A2(new_n397), .A3(new_n408), .A4(new_n401), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n403), .A2(new_n406), .A3(new_n407), .A4(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n401), .B1(new_n390), .B2(new_n397), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT6), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT30), .ZN(new_n414));
  INV_X1    g213(.A(G226gat), .ZN(new_n415));
  INV_X1    g214(.A(G233gat), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n418), .B1(new_n270), .B2(new_n235), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n256), .A2(new_n322), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n419), .B1(new_n420), .B2(new_n418), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n347), .ZN(new_n422));
  XNOR2_X1  g221(.A(G8gat), .B(G36gat), .ZN(new_n423));
  INV_X1    g222(.A(G64gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(G92gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT73), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n429), .B1(new_n420), .B2(new_n418), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n256), .A2(new_n417), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT29), .B1(new_n270), .B2(new_n235), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n431), .B1(new_n432), .B2(new_n417), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n430), .B1(new_n433), .B2(new_n429), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n422), .B(new_n428), .C1(new_n434), .C2(new_n347), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT74), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n414), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n422), .B1(new_n434), .B2(new_n347), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n427), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n435), .A2(new_n436), .A3(new_n414), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n438), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n413), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n373), .A2(new_n443), .A3(KEYINPUT35), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT35), .ZN(new_n445));
  INV_X1    g244(.A(new_n299), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n276), .A2(new_n285), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n283), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT68), .B1(new_n276), .B2(KEYINPUT32), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT32), .ZN(new_n450));
  AOI211_X1 g249(.A(new_n278), .B(new_n450), .C1(new_n274), .C2(new_n275), .ZN(new_n451));
  NOR3_X1   g250(.A1(new_n448), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n446), .B1(new_n452), .B2(new_n291), .ZN(new_n453));
  AND3_X1   g252(.A1(new_n369), .A2(new_n303), .A3(new_n370), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n303), .B1(new_n369), .B2(new_n370), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n288), .A2(new_n292), .A3(new_n299), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n453), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n410), .A2(new_n412), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n435), .A2(new_n436), .A3(new_n414), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n460), .A2(new_n437), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n459), .A2(new_n461), .A3(new_n440), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n445), .B1(new_n458), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n444), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT77), .B1(new_n383), .B2(new_n388), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n394), .A2(new_n387), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n378), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n375), .A2(KEYINPUT76), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n321), .B1(new_n208), .B2(new_n266), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n380), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n377), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n467), .A2(KEYINPUT39), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT39), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n474), .B(new_n378), .C1(new_n465), .C2(new_n466), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n473), .A2(new_n401), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT40), .ZN(new_n477));
  AND3_X1   g276(.A1(new_n476), .A2(KEYINPUT80), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n477), .B1(new_n476), .B2(KEYINPUT80), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n478), .A2(new_n479), .A3(new_n411), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n372), .B1(new_n480), .B2(new_n442), .ZN(new_n481));
  INV_X1    g280(.A(new_n435), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n439), .A2(KEYINPUT37), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT37), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n484), .B(new_n422), .C1(new_n434), .C2(new_n347), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n427), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n482), .B1(new_n486), .B2(KEYINPUT38), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT38), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n485), .A2(new_n488), .A3(new_n427), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT73), .B1(new_n432), .B2(new_n417), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n347), .B(new_n490), .C1(new_n421), .C2(KEYINPUT73), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT81), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n433), .A2(new_n429), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n494), .A2(KEYINPUT81), .A3(new_n347), .A4(new_n490), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n421), .A2(new_n347), .ZN(new_n497));
  OAI21_X1  g296(.A(KEYINPUT37), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT82), .ZN(new_n499));
  AND3_X1   g298(.A1(new_n489), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n499), .B1(new_n489), .B2(new_n498), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n413), .B(new_n487), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n481), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT83), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n481), .A2(new_n502), .A3(KEYINPUT83), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n505), .A2(new_n506), .B1(new_n372), .B2(new_n462), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT36), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n508), .B1(new_n300), .B2(new_n301), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n453), .A2(KEYINPUT36), .A3(new_n457), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n464), .B1(new_n507), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(G8gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(G15gat), .B(G22gat), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT88), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n515), .A2(G1gat), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT16), .B1(new_n515), .B2(G1gat), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT89), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n513), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n518), .B1(G1gat), .B2(new_n514), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n520), .B(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(KEYINPUT90), .ZN(new_n523));
  XNOR2_X1  g322(.A(G43gat), .B(G50gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT15), .ZN(new_n525));
  XNOR2_X1  g324(.A(KEYINPUT86), .B(G29gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(G36gat), .ZN(new_n527));
  OR3_X1    g326(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n525), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n524), .A2(KEYINPUT15), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n529), .A2(KEYINPUT85), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n529), .A2(KEYINPUT85), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n534), .A2(new_n535), .A3(new_n528), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n525), .B1(new_n536), .B2(new_n527), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n523), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(KEYINPUT91), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT87), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n541), .B1(new_n533), .B2(new_n537), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n542), .B(KEYINPUT17), .Z(new_n543));
  INV_X1    g342(.A(new_n522), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AND2_X1   g344(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(G229gat), .A2(G233gat), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n546), .A2(KEYINPUT18), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n523), .A2(new_n538), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n540), .A2(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n547), .B(KEYINPUT13), .Z(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n540), .A2(new_n547), .A3(new_n545), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT18), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n548), .A2(new_n552), .A3(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(KEYINPUT11), .B(G169gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(G197gat), .ZN(new_n558));
  XOR2_X1   g357(.A(G113gat), .B(G141gat), .Z(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n560), .B(KEYINPUT84), .Z(new_n561));
  XOR2_X1   g360(.A(new_n561), .B(KEYINPUT12), .Z(new_n562));
  NAND2_X1  g361(.A1(new_n556), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n562), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n548), .A2(new_n564), .A3(new_n552), .A4(new_n555), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT92), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n563), .A2(KEYINPUT92), .A3(new_n565), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n512), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT21), .ZN(new_n573));
  XNOR2_X1  g372(.A(G71gat), .B(G78gat), .ZN(new_n574));
  OR2_X1    g373(.A1(new_n424), .A2(G57gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n424), .A2(G57gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n574), .B1(new_n577), .B2(KEYINPUT9), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT93), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AND2_X1   g379(.A1(G71gat), .A2(G78gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n576), .B(KEYINPUT94), .ZN(new_n582));
  INV_X1    g381(.A(new_n575), .ZN(new_n583));
  OAI221_X1 g382(.A(new_n574), .B1(KEYINPUT9), .B2(new_n581), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n578), .A2(new_n579), .ZN(new_n585));
  AND3_X1   g384(.A1(new_n580), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n523), .B1(new_n573), .B2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(new_n242), .ZN(new_n589));
  XOR2_X1   g388(.A(KEYINPUT95), .B(KEYINPUT21), .Z(new_n590));
  NOR2_X1   g389(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n589), .A2(new_n591), .ZN(new_n593));
  XOR2_X1   g392(.A(G127gat), .B(G155gat), .Z(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT20), .ZN(new_n595));
  OR3_X1    g394(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n595), .B1(new_n592), .B2(new_n593), .ZN(new_n597));
  XNOR2_X1  g396(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(new_n330), .ZN(new_n599));
  NAND2_X1  g398(.A1(G231gat), .A2(G233gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  AND3_X1   g400(.A1(new_n596), .A2(new_n597), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n601), .B1(new_n596), .B2(new_n597), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT104), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT98), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n607), .A2(G85gat), .A3(G92gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT7), .ZN(new_n609));
  INV_X1    g408(.A(G106gat), .ZN(new_n610));
  OAI21_X1  g409(.A(KEYINPUT99), .B1(new_n282), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT99), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n612), .A2(G99gat), .A3(G106gat), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n611), .A2(KEYINPUT8), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT100), .B(G92gat), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n609), .B(new_n614), .C1(G85gat), .C2(new_n615), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n616), .A2(KEYINPUT101), .ZN(new_n617));
  XOR2_X1   g416(.A(G99gat), .B(G106gat), .Z(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(KEYINPUT101), .ZN(new_n619));
  AND3_X1   g418(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n618), .B1(new_n617), .B2(new_n619), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n538), .ZN(new_n623));
  NAND2_X1  g422(.A1(G232gat), .A2(G233gat), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  AOI22_X1  g424(.A1(new_n622), .A2(new_n623), .B1(KEYINPUT41), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT102), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n627), .B1(new_n620), .B2(new_n621), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n616), .B(KEYINPUT101), .ZN(new_n629));
  INV_X1    g428(.A(new_n618), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n631), .A2(KEYINPUT102), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n628), .A2(new_n543), .A3(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT103), .ZN(new_n635));
  AND3_X1   g434(.A1(new_n626), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n635), .B1(new_n626), .B2(new_n634), .ZN(new_n637));
  XOR2_X1   g436(.A(G190gat), .B(G218gat), .Z(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NOR3_X1   g438(.A1(new_n636), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n626), .A2(new_n634), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(KEYINPUT103), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n626), .A2(new_n634), .A3(new_n635), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n638), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n606), .B1(new_n640), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n639), .B1(new_n636), .B2(new_n637), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n642), .A2(new_n638), .A3(new_n643), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n646), .A2(new_n647), .A3(KEYINPUT104), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n625), .A2(KEYINPUT41), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT97), .ZN(new_n650));
  XNOR2_X1  g449(.A(G134gat), .B(G162gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n645), .A2(new_n648), .A3(new_n653), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n648), .A2(new_n653), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n605), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n622), .A2(KEYINPUT10), .A3(new_n586), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n631), .A2(new_n632), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(new_n587), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n659), .B1(new_n661), .B2(KEYINPUT10), .ZN(new_n662));
  INV_X1    g461(.A(G230gat), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n663), .A2(new_n416), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  AND2_X1   g465(.A1(new_n661), .A2(new_n664), .ZN(new_n667));
  XNOR2_X1  g466(.A(G176gat), .B(G204gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(G148gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT105), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(new_n202), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  OR3_X1    g471(.A1(new_n666), .A2(new_n667), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n672), .B1(new_n666), .B2(new_n667), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n658), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n572), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(new_n413), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(G1gat), .ZN(G1324gat));
  INV_X1    g481(.A(new_n442), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  OR2_X1    g483(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n686), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n687), .A2(KEYINPUT42), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(KEYINPUT42), .ZN(new_n689));
  OAI211_X1 g488(.A(new_n688), .B(new_n689), .C1(new_n513), .C2(new_n684), .ZN(G1325gat));
  INV_X1    g489(.A(G15gat), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT106), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n300), .A2(new_n301), .A3(new_n508), .ZN(new_n693));
  AOI21_X1  g492(.A(KEYINPUT36), .B1(new_n453), .B2(new_n457), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT106), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT107), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n679), .A2(new_n691), .A3(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n300), .A2(new_n301), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n680), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n699), .B1(new_n691), .B2(new_n701), .ZN(G1326gat));
  NOR2_X1   g501(.A1(new_n679), .A2(new_n456), .ZN(new_n703));
  XOR2_X1   g502(.A(KEYINPUT43), .B(G22gat), .Z(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(G1327gat));
  NAND3_X1  g504(.A1(new_n605), .A2(new_n676), .A3(new_n657), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n706), .A2(KEYINPUT108), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(KEYINPUT108), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n572), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(new_n459), .A3(new_n526), .ZN(new_n710));
  XOR2_X1   g509(.A(new_n710), .B(KEYINPUT45), .Z(new_n711));
  OAI21_X1  g510(.A(KEYINPUT44), .B1(new_n512), .B2(new_n656), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n462), .A2(new_n372), .ZN(new_n713));
  AOI21_X1  g512(.A(KEYINPUT83), .B1(new_n481), .B2(new_n502), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n481), .A2(new_n502), .A3(KEYINPUT83), .ZN(new_n715));
  OAI211_X1 g514(.A(new_n697), .B(new_n713), .C1(new_n714), .C2(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(KEYINPUT35), .B1(new_n373), .B2(new_n443), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n458), .A2(new_n462), .A3(new_n445), .ZN(new_n718));
  OAI21_X1  g517(.A(KEYINPUT110), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT110), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n444), .A2(new_n463), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n716), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n656), .A2(KEYINPUT111), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT111), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n654), .A2(new_n655), .A3(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n724), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT112), .B1(new_n723), .B2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT112), .ZN(new_n731));
  AOI211_X1 g530(.A(new_n731), .B(new_n728), .C1(new_n716), .C2(new_n722), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n712), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  XOR2_X1   g532(.A(new_n675), .B(KEYINPUT109), .Z(new_n734));
  NAND4_X1  g533(.A1(new_n733), .A2(new_n566), .A3(new_n605), .A4(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n526), .B1(new_n735), .B2(new_n459), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n711), .A2(new_n736), .ZN(G1328gat));
  NOR3_X1   g536(.A1(new_n709), .A2(G36gat), .A3(new_n683), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT46), .ZN(new_n739));
  OAI21_X1  g538(.A(G36gat), .B1(new_n735), .B2(new_n683), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT113), .ZN(G1329gat));
  OAI21_X1  g541(.A(G43gat), .B1(new_n735), .B2(new_n697), .ZN(new_n743));
  INV_X1    g542(.A(new_n700), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n709), .A2(G43gat), .A3(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n743), .A2(KEYINPUT47), .A3(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT114), .ZN(new_n748));
  OR2_X1    g547(.A1(new_n735), .A2(new_n698), .ZN(new_n749));
  AOI211_X1 g548(.A(new_n748), .B(new_n745), .C1(new_n749), .C2(G43gat), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n749), .A2(new_n748), .A3(G43gat), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT47), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n747), .B1(new_n750), .B2(new_n753), .ZN(G1330gat));
  OAI21_X1  g553(.A(G50gat), .B1(new_n735), .B2(new_n456), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n456), .A2(G50gat), .ZN(new_n756));
  XOR2_X1   g555(.A(new_n756), .B(KEYINPUT115), .Z(new_n757));
  OAI21_X1  g556(.A(new_n755), .B1(new_n709), .B2(new_n757), .ZN(new_n758));
  XOR2_X1   g557(.A(new_n758), .B(KEYINPUT48), .Z(G1331gat));
  INV_X1    g558(.A(new_n566), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n723), .A2(new_n760), .A3(new_n658), .ZN(new_n761));
  INV_X1    g560(.A(new_n734), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n413), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g565(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n734), .A2(new_n683), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n761), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(KEYINPUT116), .ZN(new_n770));
  NOR2_X1   g569(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n770), .B(new_n771), .ZN(G1333gat));
  OAI21_X1  g571(.A(G71gat), .B1(new_n763), .B2(new_n698), .ZN(new_n773));
  OR2_X1    g572(.A1(new_n763), .A2(G71gat), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n773), .B1(new_n774), .B2(new_n744), .ZN(new_n775));
  XOR2_X1   g574(.A(new_n775), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g575(.A1(new_n764), .A2(new_n372), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(G78gat), .ZN(G1335gat));
  OAI211_X1 g577(.A(new_n563), .B(new_n565), .C1(new_n602), .C2(new_n603), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(new_n676), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n733), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(G85gat), .B1(new_n782), .B2(new_n459), .ZN(new_n783));
  INV_X1    g582(.A(new_n779), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n723), .A2(KEYINPUT51), .A3(new_n657), .A4(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(KEYINPUT117), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n779), .B1(new_n716), .B2(new_n722), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT117), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n787), .A2(new_n788), .A3(KEYINPUT51), .A4(new_n657), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT51), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n723), .A2(new_n657), .A3(new_n784), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n786), .A2(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n792), .A2(new_n676), .ZN(new_n793));
  INV_X1    g592(.A(G85gat), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n793), .A2(new_n794), .A3(new_n413), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n783), .A2(new_n795), .ZN(G1336gat));
  INV_X1    g595(.A(KEYINPUT121), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT120), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT119), .ZN(new_n800));
  AOI211_X1 g599(.A(new_n656), .B(new_n779), .C1(new_n716), .C2(new_n722), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n800), .B1(new_n801), .B2(KEYINPUT51), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n791), .A2(KEYINPUT119), .A3(new_n790), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n786), .A2(new_n789), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n768), .A2(new_n426), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n799), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  AOI22_X1  g608(.A1(new_n802), .A2(new_n803), .B1(new_n786), .B2(new_n789), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n810), .A2(KEYINPUT120), .A3(new_n807), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n733), .A2(new_n442), .A3(new_n780), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n813), .A2(KEYINPUT118), .A3(new_n615), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT118), .B1(new_n813), .B2(new_n615), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n798), .B1(new_n812), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n813), .A2(new_n615), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n798), .B1(new_n792), .B2(new_n807), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n797), .B1(new_n817), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n815), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n806), .A2(new_n799), .A3(new_n808), .ZN(new_n824));
  OAI21_X1  g623(.A(KEYINPUT120), .B1(new_n810), .B2(new_n807), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n813), .A2(KEYINPUT118), .A3(new_n615), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n823), .A2(new_n824), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT52), .ZN(new_n828));
  INV_X1    g627(.A(new_n821), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n828), .A2(KEYINPUT121), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n822), .A2(new_n830), .ZN(G1337gat));
  OAI21_X1  g630(.A(G99gat), .B1(new_n782), .B2(new_n698), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n793), .A2(new_n282), .A3(new_n700), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(G1338gat));
  AOI21_X1  g633(.A(new_n610), .B1(new_n781), .B2(new_n372), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n734), .A2(G106gat), .A3(new_n456), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n835), .B1(new_n806), .B2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n838));
  INV_X1    g637(.A(new_n836), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n838), .B1(new_n792), .B2(new_n839), .ZN(new_n840));
  OAI22_X1  g639(.A1(new_n837), .A2(new_n838), .B1(new_n835), .B2(new_n840), .ZN(G1339gat));
  NOR4_X1   g640(.A1(new_n605), .A2(new_n566), .A3(new_n675), .A4(new_n657), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n724), .A2(new_n727), .ZN(new_n843));
  OAI21_X1  g642(.A(KEYINPUT54), .B1(new_n662), .B2(new_n665), .ZN(new_n844));
  OR2_X1    g643(.A1(new_n666), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n671), .B1(new_n666), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT55), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n845), .A2(KEYINPUT55), .A3(new_n847), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n850), .A2(new_n673), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n852), .A2(new_n760), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n546), .A2(new_n547), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n550), .A2(new_n551), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n560), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n565), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n676), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n843), .B1(new_n853), .B2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n843), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n852), .A2(new_n857), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n842), .B1(new_n863), .B2(new_n605), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n442), .A2(new_n459), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n373), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n869), .A2(new_n204), .A3(new_n566), .ZN(new_n870));
  OAI21_X1  g669(.A(G113gat), .B1(new_n868), .B2(new_n571), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(G1340gat));
  NAND3_X1  g671(.A1(new_n869), .A2(new_n202), .A3(new_n675), .ZN(new_n873));
  OAI21_X1  g672(.A(G120gat), .B1(new_n868), .B2(new_n734), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(G1341gat));
  NOR2_X1   g674(.A1(new_n868), .A2(new_n605), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n210), .A2(new_n211), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n876), .B(new_n877), .ZN(G1342gat));
  NAND3_X1  g677(.A1(new_n869), .A2(new_n262), .A3(new_n657), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n879), .A2(KEYINPUT56), .ZN(new_n880));
  OAI21_X1  g679(.A(G134gat), .B1(new_n868), .B2(new_n656), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(KEYINPUT56), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(G1343gat));
  AND3_X1   g682(.A1(new_n867), .A2(new_n372), .A3(new_n698), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n884), .A2(new_n305), .A3(new_n570), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(KEYINPUT58), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n852), .B1(new_n568), .B2(new_n569), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n656), .B1(new_n887), .B2(new_n858), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n604), .B1(new_n888), .B2(new_n862), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n372), .B1(new_n889), .B2(new_n842), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(KEYINPUT57), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n866), .B1(new_n695), .B2(new_n696), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT57), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n604), .B1(new_n859), .B2(new_n862), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n893), .B(new_n372), .C1(new_n894), .C2(new_n842), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n891), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(G141gat), .B1(new_n896), .B2(new_n571), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n886), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n891), .A2(new_n566), .A3(new_n892), .A4(new_n895), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n899), .A2(KEYINPUT122), .A3(G141gat), .ZN(new_n900));
  AOI21_X1  g699(.A(KEYINPUT122), .B1(new_n899), .B2(G141gat), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n900), .A2(new_n901), .A3(new_n885), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT58), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n898), .B1(new_n902), .B2(new_n903), .ZN(G1344gat));
  NAND3_X1  g703(.A1(new_n884), .A2(new_n306), .A3(new_n675), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n906), .B1(new_n896), .B2(new_n676), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n907), .A2(new_n306), .ZN(new_n908));
  OAI21_X1  g707(.A(KEYINPUT57), .B1(new_n864), .B2(new_n456), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n861), .A2(new_n657), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n604), .B1(new_n888), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n677), .A2(new_n570), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n893), .B(new_n372), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n909), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n675), .A3(new_n892), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n906), .B1(new_n915), .B2(G148gat), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n905), .B1(new_n908), .B2(new_n916), .ZN(G1345gat));
  NOR3_X1   g716(.A1(new_n896), .A2(new_n316), .A3(new_n605), .ZN(new_n918));
  AOI21_X1  g717(.A(G155gat), .B1(new_n884), .B2(new_n604), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n918), .A2(new_n919), .ZN(G1346gat));
  NOR3_X1   g719(.A1(new_n896), .A2(new_n317), .A3(new_n843), .ZN(new_n921));
  AOI21_X1  g720(.A(G162gat), .B1(new_n884), .B2(new_n657), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n921), .A2(new_n922), .ZN(G1347gat));
  NOR3_X1   g722(.A1(new_n864), .A2(new_n413), .A3(new_n683), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(new_n373), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n926), .A2(new_n237), .A3(new_n566), .ZN(new_n927));
  OAI21_X1  g726(.A(G169gat), .B1(new_n925), .B2(new_n571), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(G1348gat));
  NOR3_X1   g728(.A1(new_n925), .A2(new_n238), .A3(new_n734), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n926), .A2(new_n675), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n930), .B1(new_n238), .B2(new_n931), .ZN(G1349gat));
  INV_X1    g731(.A(KEYINPUT60), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(KEYINPUT123), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n242), .B1(new_n925), .B2(new_n605), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n926), .A2(new_n604), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n934), .B(new_n935), .C1(new_n936), .C2(new_n220), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n933), .A2(KEYINPUT123), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n937), .B(new_n938), .ZN(G1350gat));
  NAND3_X1  g738(.A1(new_n926), .A2(new_n221), .A3(new_n860), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n926), .A2(new_n657), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT61), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n941), .A2(new_n942), .A3(G190gat), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n942), .B1(new_n941), .B2(G190gat), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n940), .B1(new_n944), .B2(new_n945), .ZN(G1351gat));
  AND3_X1   g745(.A1(new_n698), .A2(new_n459), .A3(new_n442), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n914), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g747(.A(G197gat), .B1(new_n948), .B2(new_n571), .ZN(new_n949));
  INV_X1    g748(.A(new_n864), .ZN(new_n950));
  AND3_X1   g749(.A1(new_n950), .A2(new_n372), .A3(new_n947), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n951), .A2(new_n327), .A3(new_n566), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n949), .A2(new_n952), .ZN(G1352gat));
  OAI21_X1  g752(.A(G204gat), .B1(new_n948), .B2(new_n734), .ZN(new_n954));
  INV_X1    g753(.A(G204gat), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n951), .A2(new_n955), .A3(new_n675), .ZN(new_n956));
  AND2_X1   g755(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n957));
  NOR2_X1   g756(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OAI211_X1 g758(.A(new_n954), .B(new_n959), .C1(new_n957), .C2(new_n956), .ZN(G1353gat));
  NAND4_X1  g759(.A1(new_n909), .A2(new_n913), .A3(new_n604), .A4(new_n947), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT63), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(KEYINPUT125), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n961), .A2(G211gat), .A3(new_n963), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n962), .A2(KEYINPUT125), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n951), .A2(new_n330), .A3(new_n604), .ZN(new_n967));
  INV_X1    g766(.A(new_n965), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n961), .A2(G211gat), .A3(new_n968), .A4(new_n963), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n966), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n966), .A2(new_n967), .A3(KEYINPUT126), .A4(new_n969), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(G1354gat));
  NAND3_X1  g773(.A1(new_n951), .A2(new_n331), .A3(new_n860), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n948), .A2(KEYINPUT127), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT127), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n977), .B1(new_n914), .B2(new_n947), .ZN(new_n978));
  NOR3_X1   g777(.A1(new_n976), .A2(new_n656), .A3(new_n978), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n975), .B1(new_n979), .B2(new_n331), .ZN(G1355gat));
endmodule


