//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 1 1 0 0 0 0 1 0 1 1 0 1 0 0 0 1 1 0 0 1 1 0 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n448, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n561, new_n562, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n614, new_n616, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1147, new_n1148,
    new_n1149;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  NAND2_X1  g022(.A1(G94), .A2(G452), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT65), .Z(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(new_n462), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n470), .B1(new_n465), .B2(G125), .ZN(new_n471));
  AND2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  OAI211_X1 g048(.A(new_n470), .B(G125), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n469), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n468), .B1(new_n476), .B2(G2105), .ZN(G160));
  NOR2_X1   g052(.A1(new_n472), .A2(new_n473), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n478), .A2(new_n462), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OAI21_X1  g057(.A(KEYINPUT67), .B1(G100), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NOR3_X1   g059(.A1(KEYINPUT67), .A2(G100), .A3(G2105), .ZN(new_n485));
  OAI221_X1 g060(.A(G2104), .B1(G112), .B2(new_n462), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n480), .A2(new_n482), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  OAI211_X1 g063(.A(G138), .B(new_n462), .C1(new_n472), .C2(new_n473), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n465), .A2(new_n491), .A3(G138), .A4(new_n462), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n462), .A2(G114), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n498), .A2(new_n500), .A3(KEYINPUT69), .A4(G2104), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT68), .ZN(new_n503));
  AND2_X1   g078(.A1(G126), .A2(G2105), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n503), .B1(new_n465), .B2(new_n504), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n503), .B(new_n504), .C1(new_n472), .C2(new_n473), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n502), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n493), .A2(new_n508), .ZN(G164));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT5), .B(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G62), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n512), .A2(KEYINPUT70), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n512), .A2(KEYINPUT70), .B1(G75), .B2(G543), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n510), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  OR2_X1    g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G50), .ZN(new_n520));
  INV_X1    g095(.A(G88), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  AND2_X1   g097(.A1(KEYINPUT5), .A2(G543), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n522), .A2(new_n523), .B1(new_n516), .B2(new_n517), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n515), .A2(new_n525), .ZN(G166));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  INV_X1    g103(.A(G51), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n528), .B1(new_n519), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n523), .A2(new_n522), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n518), .A2(G89), .ZN(new_n532));
  NAND2_X1  g107(.A1(G63), .A2(G651), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n530), .A2(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  INV_X1    g111(.A(G52), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n519), .A2(new_n537), .B1(new_n538), .B2(new_n524), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n510), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n539), .A2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n531), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G651), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT71), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n546), .A2(KEYINPUT71), .A3(G651), .ZN(new_n550));
  INV_X1    g125(.A(new_n524), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n516), .A2(new_n517), .ZN(new_n552));
  INV_X1    g127(.A(G543), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(G81), .A2(new_n551), .B1(new_n554), .B2(G43), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n549), .A2(new_n550), .A3(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(G860), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT72), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  XOR2_X1   g138(.A(KEYINPUT73), .B(G65), .Z(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(new_n511), .ZN(new_n565));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(KEYINPUT74), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT74), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n565), .A2(new_n569), .A3(new_n566), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(G651), .A3(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(G53), .ZN(new_n572));
  OAI21_X1  g147(.A(KEYINPUT9), .B1(new_n519), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT9), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n554), .A2(new_n574), .A3(G53), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n573), .A2(new_n575), .B1(G91), .B2(new_n551), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n571), .A2(new_n576), .ZN(G299));
  INV_X1    g152(.A(G166), .ZN(G303));
  NAND2_X1  g153(.A1(new_n551), .A2(G87), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT75), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n511), .A2(G74), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n581), .A2(G651), .B1(new_n554), .B2(G49), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n580), .A2(new_n582), .ZN(G288));
  OAI211_X1 g158(.A(G48), .B(G543), .C1(new_n516), .C2(new_n517), .ZN(new_n584));
  INV_X1    g159(.A(G86), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n524), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g161(.A(G61), .B1(new_n523), .B2(new_n522), .ZN(new_n587));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n510), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G305));
  AND2_X1   g166(.A1(new_n511), .A2(G60), .ZN(new_n592));
  AND2_X1   g167(.A1(G72), .A2(G543), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT76), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n595), .ZN(new_n597));
  AOI22_X1  g172(.A1(G85), .A2(new_n551), .B1(new_n554), .B2(G47), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n551), .A2(G92), .ZN(new_n601));
  XOR2_X1   g176(.A(new_n601), .B(KEYINPUT10), .Z(new_n602));
  NAND2_X1  g177(.A1(G79), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G66), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n531), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n605), .A2(G651), .B1(new_n554), .B2(G54), .ZN(new_n606));
  AND2_X1   g181(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n600), .B1(new_n607), .B2(G868), .ZN(G284));
  OAI21_X1  g183(.A(new_n600), .B1(new_n607), .B2(G868), .ZN(G321));
  NAND2_X1  g184(.A1(G286), .A2(G868), .ZN(new_n610));
  INV_X1    g185(.A(G299), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G297));
  OAI21_X1  g187(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G280));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n607), .B1(new_n614), .B2(G860), .ZN(G148));
  NAND2_X1  g190(.A1(new_n607), .A2(new_n614), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G868), .ZN(new_n617));
  INV_X1    g192(.A(new_n556), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(G868), .B2(new_n618), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g195(.A1(new_n465), .A2(new_n463), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT12), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT77), .B(KEYINPUT13), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(G2100), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT78), .Z(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  INV_X1    g203(.A(G111), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(G2105), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n481), .A2(G123), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT79), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  AOI211_X1 g208(.A(new_n630), .B(new_n633), .C1(G135), .C2(new_n479), .ZN(new_n634));
  INV_X1    g209(.A(G2096), .ZN(new_n635));
  AOI22_X1  g210(.A1(new_n634), .A2(new_n635), .B1(new_n625), .B2(new_n624), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n627), .B(new_n636), .C1(new_n635), .C2(new_n634), .ZN(G156));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2430), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(KEYINPUT14), .ZN(new_n642));
  AND2_X1   g217(.A1(new_n642), .A2(KEYINPUT80), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n642), .A2(KEYINPUT80), .ZN(new_n644));
  OAI22_X1  g219(.A1(new_n643), .A2(new_n644), .B1(new_n639), .B2(new_n640), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2451), .B(G2454), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n647), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT81), .ZN(new_n653));
  INV_X1    g228(.A(G14), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n654), .B1(new_n650), .B2(new_n651), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G401));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT82), .ZN(new_n659));
  XOR2_X1   g234(.A(G2072), .B(G2078), .Z(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  NOR3_X1   g237(.A1(new_n659), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT18), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n659), .A2(new_n660), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n660), .B(KEYINPUT17), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n665), .B(new_n662), .C1(new_n659), .C2(new_n666), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n666), .A2(new_n659), .A3(new_n661), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n664), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G2096), .B(G2100), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(G227));
  XOR2_X1   g246(.A(G1971), .B(G1976), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  XOR2_X1   g248(.A(G1956), .B(G2474), .Z(new_n674));
  XOR2_X1   g249(.A(G1961), .B(G1966), .Z(new_n675));
  AND2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT20), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n674), .A2(new_n675), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  MUX2_X1   g256(.A(new_n681), .B(new_n680), .S(new_n673), .Z(new_n682));
  NOR2_X1   g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(G1981), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G1986), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT83), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n686), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(G229));
  INV_X1    g267(.A(KEYINPUT30), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n693), .A2(G28), .ZN(new_n694));
  INV_X1    g269(.A(G29), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(new_n693), .B2(G28), .ZN(new_n696));
  AND2_X1   g271(.A1(KEYINPUT31), .A2(G11), .ZN(new_n697));
  NOR2_X1   g272(.A1(KEYINPUT31), .A2(G11), .ZN(new_n698));
  OAI22_X1  g273(.A1(new_n694), .A2(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(new_n634), .B2(G29), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G21), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G168), .B2(new_n701), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n700), .B1(G1966), .B2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(G33), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n705), .A2(G29), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT87), .B(KEYINPUT25), .Z(new_n707));
  NAND3_X1  g282(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n479), .A2(G139), .ZN(new_n710));
  AOI22_X1  g285(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n709), .B(new_n710), .C1(new_n462), .C2(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n706), .B1(new_n712), .B2(G29), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(new_n442), .ZN(new_n714));
  NAND2_X1  g289(.A1(G301), .A2(G16), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n701), .A2(G5), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n714), .B1(new_n717), .B2(G1961), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(G1961), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(new_n442), .B2(new_n713), .ZN(new_n720));
  NOR3_X1   g295(.A1(new_n704), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n695), .B1(KEYINPUT24), .B2(G34), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(KEYINPUT24), .B2(G34), .ZN(new_n723));
  INV_X1    g298(.A(G160), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(G29), .ZN(new_n725));
  INV_X1    g300(.A(G2084), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT93), .Z(new_n728));
  NAND2_X1  g303(.A1(new_n703), .A2(G1966), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT92), .ZN(new_n730));
  NOR2_X1   g305(.A1(G27), .A2(G29), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G164), .B2(G29), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G2078), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n721), .A2(new_n728), .A3(new_n730), .A4(new_n734), .ZN(new_n735));
  NAND3_X1  g310(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT89), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT26), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n479), .A2(G141), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n481), .A2(G129), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n463), .A2(G105), .ZN(new_n741));
  NAND4_X1  g316(.A1(new_n738), .A2(new_n739), .A3(new_n740), .A4(new_n741), .ZN(new_n742));
  MUX2_X1   g317(.A(G32), .B(new_n742), .S(G29), .Z(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT90), .Z(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT27), .B(G1996), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT91), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n744), .B(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n725), .A2(new_n726), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT88), .Z(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  NOR3_X1   g325(.A1(new_n735), .A2(new_n747), .A3(new_n750), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n751), .A2(KEYINPUT94), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n751), .A2(KEYINPUT94), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n701), .A2(G4), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n607), .B2(new_n701), .ZN(new_n755));
  INV_X1    g330(.A(G1348), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n479), .A2(G140), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n481), .A2(G128), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n462), .A2(G116), .ZN(new_n760));
  OAI21_X1  g335(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n758), .B(new_n759), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(G29), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n695), .A2(G26), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT28), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(G2067), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(G29), .A2(G35), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G162), .B2(G29), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n772), .A2(G2090), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n757), .B(new_n768), .C1(new_n773), .C2(KEYINPUT96), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(KEYINPUT96), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n701), .A2(G20), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT23), .Z(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G299), .B2(G16), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G1956), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n774), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(G1341), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n618), .A2(G16), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G16), .B2(G19), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n772), .A2(G2090), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n781), .B(new_n785), .C1(new_n782), .C2(new_n784), .ZN(new_n786));
  NOR3_X1   g361(.A1(new_n752), .A2(new_n753), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n701), .A2(G23), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n580), .A2(new_n582), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(new_n789), .B2(new_n701), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT33), .B(G1976), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n701), .A2(G22), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G166), .B2(new_n701), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(G1971), .Z(new_n795));
  NOR2_X1   g370(.A1(G6), .A2(G16), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n590), .B2(G16), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT32), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(new_n684), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n792), .A2(new_n795), .A3(new_n799), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n800), .A2(KEYINPUT34), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(KEYINPUT34), .ZN(new_n802));
  MUX2_X1   g377(.A(G24), .B(G290), .S(G16), .Z(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(G1986), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n479), .A2(G131), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n481), .A2(G119), .ZN(new_n806));
  OAI21_X1  g381(.A(KEYINPUT85), .B1(G95), .B2(G2105), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  NOR3_X1   g383(.A1(KEYINPUT85), .A2(G95), .A3(G2105), .ZN(new_n809));
  OAI221_X1 g384(.A(G2104), .B1(G107), .B2(new_n462), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n805), .A2(new_n806), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(G29), .ZN(new_n812));
  INV_X1    g387(.A(G25), .ZN(new_n813));
  OR3_X1    g388(.A1(new_n813), .A2(KEYINPUT84), .A3(G29), .ZN(new_n814));
  OAI21_X1  g389(.A(KEYINPUT84), .B1(new_n813), .B2(G29), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n812), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT35), .B(G1991), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n801), .A2(new_n802), .A3(new_n804), .A4(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT36), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n820), .A2(KEYINPUT86), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n819), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n787), .A2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(G311));
  XNOR2_X1  g399(.A(new_n823), .B(KEYINPUT97), .ZN(G150));
  NAND2_X1  g400(.A1(new_n554), .A2(G55), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT99), .B(G93), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n828));
  OAI221_X1 g403(.A(new_n826), .B1(new_n524), .B2(new_n827), .C1(new_n510), .C2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(G860), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT37), .Z(new_n831));
  NAND2_X1  g406(.A1(new_n607), .A2(G559), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n556), .B(new_n829), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n834), .B(new_n835), .Z(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n557), .B1(new_n837), .B2(KEYINPUT39), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n831), .B1(new_n838), .B2(new_n839), .ZN(G145));
  XNOR2_X1  g415(.A(new_n742), .B(new_n712), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n762), .ZN(new_n842));
  OAI21_X1  g417(.A(KEYINPUT100), .B1(new_n493), .B2(new_n508), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n504), .B1(new_n472), .B2(new_n473), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(KEYINPUT68), .ZN(new_n845));
  AOI22_X1  g420(.A1(new_n845), .A2(new_n506), .B1(new_n497), .B2(new_n501), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT100), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n490), .A2(new_n492), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n843), .A2(new_n849), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n842), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n842), .A2(new_n850), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n811), .B(KEYINPUT101), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n622), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n481), .A2(G130), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n462), .A2(G118), .ZN(new_n857));
  OAI21_X1  g432(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n859), .B1(G142), .B2(new_n479), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n855), .B(new_n860), .ZN(new_n861));
  OR3_X1    g436(.A1(new_n853), .A2(KEYINPUT102), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n853), .B1(KEYINPUT102), .B2(new_n861), .ZN(new_n863));
  XNOR2_X1  g438(.A(G160), .B(G162), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n634), .B(new_n864), .Z(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n862), .A2(new_n863), .A3(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(G37), .ZN(new_n868));
  NOR3_X1   g443(.A1(new_n851), .A2(new_n861), .A3(new_n852), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n861), .B1(new_n851), .B2(new_n852), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(new_n865), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n867), .B(new_n868), .C1(new_n869), .C2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g448(.A(KEYINPUT106), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n607), .A2(G299), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n875), .A2(KEYINPUT103), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(KEYINPUT103), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n607), .A2(G299), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT41), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n607), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n611), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n878), .ZN(new_n884));
  OR3_X1    g459(.A1(new_n884), .A2(KEYINPUT104), .A3(new_n880), .ZN(new_n885));
  OAI21_X1  g460(.A(KEYINPUT104), .B1(new_n884), .B2(new_n880), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n881), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n616), .B(new_n835), .Z(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n889), .A2(KEYINPUT105), .ZN(new_n890));
  INV_X1    g465(.A(new_n884), .ZN(new_n891));
  OAI211_X1 g466(.A(new_n889), .B(KEYINPUT105), .C1(new_n888), .C2(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n874), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n890), .A2(new_n892), .A3(new_n874), .ZN(new_n894));
  XNOR2_X1  g469(.A(G288), .B(G166), .ZN(new_n895));
  XNOR2_X1  g470(.A(G290), .B(new_n590), .ZN(new_n896));
  XOR2_X1   g471(.A(new_n895), .B(new_n896), .Z(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT42), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n893), .B1(new_n894), .B2(new_n899), .ZN(new_n900));
  AOI211_X1 g475(.A(new_n874), .B(new_n898), .C1(new_n890), .C2(new_n892), .ZN(new_n901));
  OAI21_X1  g476(.A(G868), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(G868), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n829), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(G295));
  NAND2_X1  g480(.A1(new_n902), .A2(new_n904), .ZN(G331));
  XNOR2_X1  g481(.A(new_n835), .B(G301), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n907), .A2(G168), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(G168), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(new_n891), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n911), .B1(new_n887), .B2(new_n910), .ZN(new_n912));
  INV_X1    g487(.A(new_n897), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(G37), .B1(new_n912), .B2(new_n913), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n916), .A2(KEYINPUT43), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n891), .B1(new_n910), .B2(new_n880), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT107), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n908), .A2(new_n879), .A3(KEYINPUT41), .A4(new_n909), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n918), .A2(new_n919), .A3(new_n897), .A4(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n918), .A2(new_n897), .A3(new_n920), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(KEYINPUT107), .ZN(new_n923));
  AND4_X1   g498(.A1(KEYINPUT43), .A2(new_n915), .A3(new_n921), .A4(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT44), .B1(new_n917), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT43), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n915), .A2(new_n923), .A3(new_n926), .A4(new_n921), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n927), .B1(new_n916), .B2(new_n926), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n925), .A2(new_n930), .ZN(G397));
  AOI22_X1  g506(.A1(new_n479), .A2(G137), .B1(G101), .B2(new_n463), .ZN(new_n932));
  XOR2_X1   g507(.A(KEYINPUT109), .B(G40), .Z(new_n933));
  INV_X1    g508(.A(new_n469), .ZN(new_n934));
  OAI21_X1  g509(.A(G125), .B1(new_n472), .B2(new_n473), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT66), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n934), .B1(new_n936), .B2(new_n474), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n932), .B(new_n933), .C1(new_n937), .C2(new_n462), .ZN(new_n938));
  XNOR2_X1  g513(.A(KEYINPUT108), .B(G1384), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  AOI211_X1 g515(.A(KEYINPUT45), .B(new_n938), .C1(new_n850), .C2(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n742), .B(G1996), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n762), .B(new_n767), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n811), .B(new_n817), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(G290), .B(G1986), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n941), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT125), .ZN(new_n950));
  INV_X1    g525(.A(G1966), .ZN(new_n951));
  AOI21_X1  g526(.A(G1384), .B1(new_n846), .B2(new_n848), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT45), .ZN(new_n953));
  OAI211_X1 g528(.A(G160), .B(new_n933), .C1(new_n952), .C2(KEYINPUT45), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT114), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(G1384), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n957), .B1(new_n493), .B2(new_n508), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT45), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n938), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT114), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n951), .B1(new_n956), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT115), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n938), .B1(new_n958), .B2(new_n959), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT114), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n954), .A2(new_n955), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n966), .A2(new_n967), .A3(new_n953), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT115), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n968), .A2(new_n969), .A3(new_n951), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT50), .ZN(new_n971));
  OAI211_X1 g546(.A(G160), .B(new_n933), .C1(new_n952), .C2(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n958), .A2(KEYINPUT50), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  XOR2_X1   g549(.A(KEYINPUT116), .B(G2084), .Z(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n964), .A2(G168), .A3(new_n970), .A4(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT51), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n977), .A2(new_n978), .A3(G8), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n958), .A2(new_n959), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n980), .B1(new_n965), .B2(KEYINPUT114), .ZN(new_n981));
  AOI21_X1  g556(.A(G1966), .B1(new_n981), .B2(new_n967), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n976), .B1(new_n982), .B2(new_n969), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n963), .A2(KEYINPUT115), .ZN(new_n984));
  OAI21_X1  g559(.A(G286), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n985), .A2(G8), .A3(new_n977), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n979), .B1(KEYINPUT51), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT62), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n950), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n789), .A2(G1976), .ZN(new_n990));
  INV_X1    g565(.A(G1976), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT52), .B1(G288), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(G160), .A2(new_n952), .A3(new_n933), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT112), .B1(new_n993), .B2(G8), .ZN(new_n994));
  OAI211_X1 g569(.A(KEYINPUT112), .B(G8), .C1(new_n958), .C2(new_n938), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n990), .B(new_n992), .C1(new_n994), .C2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n589), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n518), .A2(G86), .A3(new_n511), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n998), .A2(new_n999), .A3(new_n684), .A4(new_n584), .ZN(new_n1000));
  OAI21_X1  g575(.A(G1981), .B1(new_n586), .B2(new_n589), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT113), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT49), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1000), .A2(new_n1001), .A3(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n1005), .B(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(new_n994), .B2(new_n996), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n1009));
  OAI21_X1  g584(.A(G8), .B1(new_n958), .B2(new_n938), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT112), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n1012), .A2(new_n995), .B1(G1976), .B2(new_n789), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n997), .B(new_n1008), .C1(new_n1009), .C2(new_n1013), .ZN(new_n1014));
  AND2_X1   g589(.A1(G303), .A2(G8), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n1015), .B(KEYINPUT55), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G2090), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n974), .A2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n939), .A2(new_n959), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n843), .A2(new_n849), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT110), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n843), .A2(KEYINPUT110), .A3(new_n849), .A4(new_n1020), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n954), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1019), .B1(new_n1025), .B2(G1971), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(G8), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1014), .B1(new_n1017), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(KEYINPUT111), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT111), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1030), .B(new_n1019), .C1(new_n1025), .C2(G1971), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1029), .A2(G8), .A3(new_n1016), .A4(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n974), .A2(G1961), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1025), .A2(new_n443), .ZN(new_n1034));
  XOR2_X1   g609(.A(KEYINPUT123), .B(KEYINPUT53), .Z(new_n1035));
  AOI21_X1  g610(.A(new_n1033), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n443), .A2(KEYINPUT53), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1036), .B1(new_n968), .B2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1028), .A2(new_n1032), .A3(new_n1038), .A4(G171), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1039), .B1(new_n987), .B2(new_n988), .ZN(new_n1040));
  INV_X1    g615(.A(new_n979), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n977), .A2(G8), .ZN(new_n1042));
  AOI22_X1  g617(.A1(new_n963), .A2(KEYINPUT115), .B1(new_n974), .B2(new_n975), .ZN(new_n1043));
  AOI21_X1  g618(.A(G168), .B1(new_n1043), .B2(new_n970), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT51), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1041), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1046), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n989), .A2(new_n1040), .A3(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g623(.A(G301), .B(KEYINPUT54), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n443), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n937), .A2(KEYINPUT124), .ZN(new_n1051));
  OAI21_X1  g626(.A(G2105), .B1(new_n937), .B2(KEYINPUT124), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n932), .B(new_n1050), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n850), .A2(new_n940), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1053), .B1(new_n1054), .B2(new_n959), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1049), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AOI22_X1  g632(.A1(new_n1038), .A2(new_n1049), .B1(new_n1057), .B2(new_n1036), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1058), .A2(new_n1032), .A3(new_n1028), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n987), .A2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n756), .B1(new_n972), .B2(new_n973), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n961), .A2(new_n767), .A3(new_n952), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(KEYINPUT60), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT122), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1063), .A2(new_n1064), .A3(new_n882), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n882), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1066));
  OAI22_X1  g641(.A1(new_n1065), .A2(new_n1066), .B1(new_n1064), .B2(new_n1063), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT60), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1067), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(G1996), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1025), .A2(new_n1072), .ZN(new_n1073));
  XOR2_X1   g648(.A(KEYINPUT58), .B(G1341), .Z(new_n1074));
  NAND2_X1  g649(.A1(new_n993), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT59), .B1(new_n1076), .B2(new_n618), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT59), .ZN(new_n1078));
  AOI211_X1 g653(.A(new_n1078), .B(new_n556), .C1(new_n1073), .C2(new_n1075), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT61), .ZN(new_n1081));
  XNOR2_X1  g656(.A(KEYINPUT56), .B(G2072), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1025), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n1084));
  OR2_X1    g659(.A1(new_n1084), .A2(KEYINPUT57), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(KEYINPUT57), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n611), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(G299), .A2(new_n1084), .A3(KEYINPUT57), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  OR2_X1    g664(.A1(new_n974), .A2(G1956), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1083), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1089), .B1(new_n1083), .B2(new_n1090), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1081), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1071), .A2(new_n1080), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1091), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1083), .A2(new_n1089), .A3(new_n1090), .A4(KEYINPUT120), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1097), .A2(new_n1098), .A3(KEYINPUT61), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT121), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1097), .A2(new_n1098), .A3(new_n1101), .A4(KEYINPUT61), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1095), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1093), .B1(new_n607), .B2(new_n1068), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1104), .A2(new_n1092), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1060), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1008), .A2(new_n991), .A3(new_n789), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n1000), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(new_n996), .B2(new_n994), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(new_n1032), .B2(new_n1014), .ZN(new_n1110));
  NAND2_X1  g685(.A1(G168), .A2(G8), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1111), .B1(new_n1043), .B2(new_n970), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1028), .A2(new_n1032), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT63), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT117), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1029), .A2(G8), .A3(new_n1031), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n1017), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1014), .A2(new_n1114), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1032), .A2(new_n1112), .A3(new_n1119), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1115), .A2(new_n1116), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1113), .A2(KEYINPUT117), .A3(new_n1114), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1110), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1048), .B(new_n1106), .C1(new_n1123), .C2(KEYINPUT118), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT118), .ZN(new_n1125));
  AOI211_X1 g700(.A(new_n1125), .B(new_n1110), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n949), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n941), .A2(new_n1072), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n1128), .B(KEYINPUT46), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n941), .B1(new_n742), .B2(new_n944), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  XOR2_X1   g706(.A(new_n1131), .B(KEYINPUT126), .Z(new_n1132));
  OR2_X1    g707(.A1(new_n1132), .A2(KEYINPUT47), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(KEYINPUT47), .ZN(new_n1134));
  NOR2_X1   g709(.A1(G290), .A2(G1986), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n941), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1136), .ZN(new_n1137));
  OR2_X1    g712(.A1(new_n1137), .A2(KEYINPUT48), .ZN(new_n1138));
  AOI22_X1  g713(.A1(new_n1137), .A2(KEYINPUT48), .B1(new_n947), .B2(new_n941), .ZN(new_n1139));
  INV_X1    g714(.A(new_n811), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n945), .A2(new_n817), .A3(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1141), .B1(G2067), .B2(new_n762), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1138), .A2(new_n1139), .B1(new_n941), .B2(new_n1142), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1133), .A2(new_n1134), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1127), .A2(new_n1144), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g720(.A(G319), .ZN(new_n1147));
  NOR2_X1   g721(.A1(G227), .A2(new_n1147), .ZN(new_n1148));
  AND2_X1   g722(.A1(new_n691), .A2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g723(.A1(new_n928), .A2(new_n656), .A3(new_n1149), .A4(new_n872), .ZN(G225));
  INV_X1    g724(.A(G225), .ZN(G308));
endmodule


