//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 1 0 1 0 0 1 0 1 0 0 1 0 0 1 0 1 0 0 0 1 0 0 1 1 0 0 0 0 0 1 1 1 1 0 0 0 0 1 0 0 0 1 1 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017;
  XNOR2_X1  g000(.A(KEYINPUT71), .B(G237), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G210), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT27), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT26), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT27), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n189), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT26), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  AND3_X1   g009(.A1(new_n191), .A2(new_n195), .A3(G101), .ZN(new_n196));
  AOI21_X1  g010(.A(G101), .B1(new_n191), .B2(new_n195), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(KEYINPUT72), .B(KEYINPUT28), .ZN(new_n199));
  INV_X1    g013(.A(G143), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT64), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G146), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n200), .B1(new_n202), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT0), .ZN(new_n206));
  INV_X1    g020(.A(G128), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n201), .A2(G143), .ZN(new_n208));
  NOR4_X1   g022(.A1(new_n205), .A2(new_n206), .A3(new_n207), .A4(new_n208), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n206), .A2(new_n207), .ZN(new_n210));
  NOR2_X1   g024(.A1(KEYINPUT0), .A2(G128), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n202), .A2(new_n204), .A3(new_n200), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n200), .A2(G146), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  AOI211_X1 g028(.A(new_n210), .B(new_n211), .C1(new_n212), .C2(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n209), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT11), .ZN(new_n217));
  INV_X1    g031(.A(G134), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n217), .B1(new_n218), .B2(G137), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(G137), .ZN(new_n220));
  INV_X1    g034(.A(G137), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(KEYINPUT11), .A3(G134), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n219), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G131), .ZN(new_n224));
  INV_X1    g038(.A(G131), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n219), .A2(new_n222), .A3(new_n225), .A4(new_n220), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n227));
  AND2_X1   g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n226), .A2(new_n227), .ZN(new_n229));
  OAI211_X1 g043(.A(KEYINPUT70), .B(new_n224), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  AND2_X1   g045(.A1(new_n219), .A2(new_n222), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n232), .A2(KEYINPUT66), .A3(new_n225), .A4(new_n220), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n226), .A2(new_n227), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT70), .B1(new_n235), .B2(new_n224), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n216), .B1(new_n231), .B2(new_n236), .ZN(new_n237));
  XOR2_X1   g051(.A(KEYINPUT2), .B(G113), .Z(new_n238));
  INV_X1    g052(.A(G116), .ZN(new_n239));
  NOR3_X1   g053(.A1(new_n239), .A2(KEYINPUT69), .A3(G119), .ZN(new_n240));
  INV_X1    g054(.A(G119), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G116), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n243), .B1(new_n241), .B2(G116), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n240), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n238), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n244), .A2(new_n242), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n243), .A2(new_n241), .A3(G116), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n238), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n250), .A2(new_n251), .A3(KEYINPUT68), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n247), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  AND2_X1   g068(.A1(KEYINPUT67), .A2(G128), .ZN(new_n255));
  NOR2_X1   g069(.A1(KEYINPUT67), .A2(G128), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT1), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n257), .B1(new_n205), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n212), .A2(new_n214), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n205), .A2(new_n208), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n207), .A2(KEYINPUT1), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  XOR2_X1   g079(.A(G134), .B(G137), .Z(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G131), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n265), .A2(new_n235), .A3(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n237), .A2(new_n254), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT65), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n270), .B1(new_n209), .B2(new_n215), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n224), .B1(new_n228), .B2(new_n229), .ZN(new_n272));
  INV_X1    g086(.A(new_n210), .ZN(new_n273));
  INV_X1    g087(.A(new_n211), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n260), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n202), .A2(new_n204), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G143), .ZN(new_n277));
  INV_X1    g091(.A(new_n208), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n277), .A2(new_n278), .A3(new_n210), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n275), .A2(KEYINPUT65), .A3(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n271), .A2(new_n272), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n268), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n253), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n199), .B1(new_n269), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n275), .A2(new_n279), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT70), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n272), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n285), .B1(new_n287), .B2(new_n230), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n265), .A2(new_n235), .A3(new_n267), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT28), .B1(new_n290), .B2(new_n254), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n198), .B1(new_n284), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n237), .A2(KEYINPUT30), .A3(new_n268), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT30), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n282), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n293), .A2(new_n253), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n191), .A2(new_n195), .ZN(new_n297));
  INV_X1    g111(.A(G101), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n191), .A2(new_n195), .A3(G101), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n296), .A2(new_n301), .A3(new_n269), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT29), .B1(new_n292), .B2(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n254), .B1(new_n237), .B2(new_n268), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n288), .A2(new_n253), .A3(new_n289), .ZN(new_n305));
  OAI21_X1  g119(.A(KEYINPUT28), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n299), .A2(KEYINPUT29), .A3(new_n300), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT28), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n269), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n306), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G902), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(G472), .B1(new_n303), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT73), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n296), .A2(new_n198), .A3(new_n269), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT31), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n301), .B1(new_n284), .B2(new_n291), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT31), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n296), .A2(new_n198), .A3(new_n319), .A4(new_n269), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n317), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  NOR2_X1   g135(.A1(G472), .A2(G902), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT32), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n321), .A2(KEYINPUT32), .A3(new_n322), .ZN(new_n326));
  OAI211_X1 g140(.A(KEYINPUT73), .B(G472), .C1(new_n303), .C2(new_n312), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n315), .A2(new_n325), .A3(new_n326), .A4(new_n327), .ZN(new_n328));
  XOR2_X1   g142(.A(KEYINPUT71), .B(G237), .Z(new_n329));
  INV_X1    g143(.A(G953), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(G214), .A3(new_n330), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n331), .A2(new_n200), .ZN(new_n332));
  AOI21_X1  g146(.A(G143), .B1(new_n188), .B2(G214), .ZN(new_n333));
  OAI21_X1  g147(.A(G131), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT17), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n331), .A2(new_n200), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n188), .A2(G143), .A3(G214), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n225), .A3(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n334), .A2(new_n335), .A3(new_n338), .ZN(new_n339));
  OAI211_X1 g153(.A(KEYINPUT17), .B(G131), .C1(new_n332), .C2(new_n333), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT89), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(G125), .B(G140), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT16), .ZN(new_n344));
  INV_X1    g158(.A(G125), .ZN(new_n345));
  OR3_X1    g159(.A1(new_n345), .A2(KEYINPUT16), .A3(G140), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n201), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n344), .A2(G146), .A3(new_n346), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n225), .B1(new_n336), .B2(new_n337), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n352), .A2(KEYINPUT89), .A3(KEYINPUT17), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n339), .A2(new_n342), .A3(new_n351), .A4(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(G113), .B(G122), .ZN(new_n355));
  INV_X1    g169(.A(G104), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n355), .B(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT18), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n336), .B(new_n337), .C1(new_n358), .C2(new_n225), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n276), .A2(new_n343), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n360), .B1(new_n201), .B2(new_n343), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n359), .B(new_n361), .C1(new_n334), .C2(new_n358), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n354), .A2(new_n357), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n349), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT19), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n365), .A2(KEYINPUT87), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n343), .A2(new_n366), .ZN(new_n367));
  XOR2_X1   g181(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n368));
  OAI21_X1  g182(.A(new_n367), .B1(new_n343), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n276), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n364), .B1(new_n370), .B2(KEYINPUT88), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT88), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n369), .A2(new_n372), .A3(new_n276), .ZN(new_n373));
  INV_X1    g187(.A(new_n338), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n371), .B(new_n373), .C1(new_n374), .C2(new_n352), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n362), .ZN(new_n376));
  INV_X1    g190(.A(new_n357), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n363), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G475), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(new_n311), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT20), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n363), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n357), .B1(new_n354), .B2(new_n362), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n311), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G475), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n379), .A2(KEYINPUT20), .A3(new_n380), .A4(new_n311), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n383), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  XOR2_X1   g203(.A(KEYINPUT9), .B(G234), .Z(new_n390));
  NAND3_X1  g204(.A1(new_n390), .A2(G217), .A3(new_n330), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT67), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n207), .ZN(new_n393));
  NAND2_X1  g207(.A1(KEYINPUT67), .A2(G128), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G143), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n207), .A2(G143), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n399), .A2(G134), .ZN(new_n400));
  XOR2_X1   g214(.A(G116), .B(G122), .Z(new_n401));
  INV_X1    g215(.A(G107), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n401), .B(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n396), .A2(KEYINPUT13), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT90), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n404), .A2(new_n405), .A3(new_n398), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT13), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n398), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n407), .B1(new_n395), .B2(G143), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT90), .B1(new_n410), .B2(new_n397), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n406), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  AOI211_X1 g226(.A(new_n400), .B(new_n403), .C1(new_n412), .C2(G134), .ZN(new_n413));
  INV_X1    g227(.A(new_n400), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n399), .A2(G134), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OR2_X1    g230(.A1(new_n239), .A2(G122), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n402), .B1(new_n417), .B2(KEYINPUT14), .ZN(new_n418));
  OR2_X1    g232(.A1(new_n418), .A2(new_n401), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n401), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n416), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n391), .B1(new_n413), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n412), .A2(G134), .ZN(new_n423));
  INV_X1    g237(.A(new_n403), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(new_n414), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n416), .A2(new_n419), .A3(new_n420), .ZN(new_n426));
  INV_X1    g240(.A(new_n391), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n422), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n311), .ZN(new_n430));
  INV_X1    g244(.A(G478), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT91), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n432), .A2(KEYINPUT15), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(KEYINPUT15), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n431), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n430), .B(new_n436), .ZN(new_n437));
  OR2_X1    g251(.A1(new_n389), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(KEYINPUT3), .B1(new_n356), .B2(G107), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT3), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(new_n402), .A3(G104), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n356), .A2(G107), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n439), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT4), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n443), .A2(new_n444), .A3(G101), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT79), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n443), .A2(KEYINPUT79), .A3(new_n444), .A4(G101), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n443), .A2(G101), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n439), .A2(new_n441), .A3(new_n298), .A4(new_n442), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n450), .A2(KEYINPUT4), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n449), .A2(new_n253), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(KEYINPUT69), .B1(new_n239), .B2(G119), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n239), .A2(G119), .ZN(new_n455));
  OAI211_X1 g269(.A(KEYINPUT5), .B(new_n249), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G113), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT5), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n457), .B1(new_n455), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT83), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n442), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n356), .A2(G107), .ZN(new_n464));
  OAI21_X1  g278(.A(G101), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n451), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n245), .A2(new_n238), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n456), .A2(KEYINPUT83), .A3(new_n459), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n462), .A2(new_n467), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n453), .A2(new_n470), .ZN(new_n471));
  XOR2_X1   g285(.A(G110), .B(G122), .Z(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n472), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n453), .A2(new_n470), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n473), .A2(KEYINPUT6), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT6), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n471), .A2(new_n477), .A3(new_n472), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n275), .A2(G125), .A3(new_n279), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(G125), .B1(new_n261), .B2(new_n264), .ZN(new_n481));
  OAI211_X1 g295(.A(G224), .B(new_n330), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n265), .A2(new_n345), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n330), .A2(G224), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(new_n479), .A3(new_n484), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n476), .A2(new_n478), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n456), .A2(KEYINPUT84), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT84), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n248), .A2(new_n489), .A3(KEYINPUT5), .A4(new_n249), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n488), .A2(new_n459), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n468), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT85), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT85), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n491), .A2(new_n494), .A3(new_n468), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n493), .A2(new_n467), .A3(new_n495), .ZN(new_n496));
  XOR2_X1   g310(.A(new_n472), .B(KEYINPUT8), .Z(new_n497));
  NAND4_X1  g311(.A1(new_n462), .A2(new_n466), .A3(new_n468), .A4(new_n469), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n484), .A2(KEYINPUT7), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  OAI22_X1  g315(.A1(new_n480), .A2(new_n481), .B1(KEYINPUT86), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT86), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n502), .B1(new_n503), .B2(new_n500), .ZN(new_n504));
  OAI211_X1 g318(.A(KEYINPUT86), .B(new_n501), .C1(new_n480), .C2(new_n481), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n499), .A2(new_n504), .A3(new_n475), .A4(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n487), .A2(new_n311), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(G210), .B1(G237), .B2(G902), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n487), .A2(new_n311), .A3(new_n506), .A4(new_n508), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(G234), .A2(G237), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n513), .A2(G952), .A3(new_n330), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT21), .B(G898), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n515), .B(KEYINPUT92), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n513), .A2(G902), .A3(G953), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n514), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(G214), .B1(G237), .B2(G902), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n512), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n438), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g337(.A(G110), .B(G140), .ZN(new_n524));
  AND2_X1   g338(.A1(new_n330), .A2(G227), .ZN(new_n525));
  XOR2_X1   g339(.A(new_n524), .B(new_n525), .Z(new_n526));
  OAI21_X1  g340(.A(KEYINPUT1), .B1(new_n200), .B2(G146), .ZN(new_n527));
  OR2_X1    g341(.A1(new_n527), .A2(KEYINPUT80), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n207), .B1(new_n527), .B2(KEYINPUT80), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n528), .A2(new_n529), .B1(new_n277), .B2(new_n278), .ZN(new_n530));
  NOR4_X1   g344(.A1(new_n205), .A2(KEYINPUT1), .A3(new_n207), .A4(new_n208), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n467), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT10), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n216), .A2(new_n449), .A3(new_n452), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n265), .A2(KEYINPUT10), .A3(new_n467), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n287), .A2(new_n230), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n526), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT82), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n261), .A2(new_n466), .A3(new_n264), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n532), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n538), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT12), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n543), .A2(KEYINPUT12), .A3(new_n272), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT81), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n543), .A2(KEYINPUT81), .A3(KEYINPUT12), .A4(new_n272), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n546), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n231), .A2(new_n236), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n552), .A2(new_n534), .A3(new_n535), .A4(new_n536), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n553), .A2(KEYINPUT82), .A3(new_n526), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n541), .A2(new_n551), .A3(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n526), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n537), .A2(new_n538), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n537), .A2(new_n538), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(G902), .B1(new_n555), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(G469), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n557), .A2(new_n558), .A3(new_n556), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n551), .A2(new_n553), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n563), .B1(new_n564), .B2(new_n556), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(G469), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n561), .A2(new_n311), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n562), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n390), .ZN(new_n570));
  OAI21_X1  g384(.A(G221), .B1(new_n570), .B2(G902), .ZN(new_n571));
  XOR2_X1   g385(.A(new_n571), .B(KEYINPUT78), .Z(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n241), .B1(new_n393), .B2(new_n394), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n207), .A2(G119), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT24), .B(G110), .ZN(new_n578));
  OR4_X1    g392(.A1(KEYINPUT74), .A2(new_n576), .A3(new_n577), .A4(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(KEYINPUT23), .B1(new_n207), .B2(G119), .ZN(new_n580));
  OAI21_X1  g394(.A(KEYINPUT75), .B1(new_n241), .B2(G128), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT75), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n582), .A2(new_n207), .A3(G119), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  OAI211_X1 g398(.A(KEYINPUT23), .B(G119), .C1(new_n255), .C2(new_n256), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(G110), .ZN(new_n587));
  INV_X1    g401(.A(new_n578), .ZN(new_n588));
  INV_X1    g402(.A(new_n577), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n588), .B(new_n589), .C1(new_n241), .C2(new_n257), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(KEYINPUT74), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n350), .A2(new_n579), .A3(new_n587), .A4(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT76), .ZN(new_n593));
  INV_X1    g407(.A(G110), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n584), .A2(new_n594), .A3(new_n585), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n578), .B1(new_n576), .B2(new_n577), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AND4_X1   g411(.A1(new_n593), .A2(new_n597), .A3(new_n360), .A4(new_n349), .ZN(new_n598));
  INV_X1    g412(.A(new_n360), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n599), .B1(new_n595), .B2(new_n596), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n593), .B1(new_n600), .B2(new_n349), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n592), .B1(new_n598), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n330), .A2(G221), .A3(G234), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(KEYINPUT22), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G137), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n592), .B(new_n605), .C1(new_n598), .C2(new_n601), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n607), .A2(new_n311), .A3(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT77), .ZN(new_n610));
  AOI21_X1  g424(.A(KEYINPUT25), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(G217), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n613), .B1(G234), .B2(new_n311), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n609), .A2(new_n610), .A3(KEYINPUT25), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n612), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n614), .A2(G902), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n607), .A2(new_n608), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n328), .A2(new_n523), .A3(new_n575), .A4(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G101), .ZN(G3));
  NAND2_X1  g436(.A1(new_n321), .A2(new_n311), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(G472), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n323), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n625), .A2(new_n574), .A3(new_n619), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT93), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n510), .A2(new_n627), .A3(new_n511), .ZN(new_n628));
  OR2_X1    g442(.A1(new_n511), .A2(new_n627), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n628), .A2(new_n629), .A3(new_n520), .A4(new_n521), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT94), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT33), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(KEYINPUT94), .A2(KEYINPUT33), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n429), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n422), .A2(new_n428), .A3(new_n631), .A4(new_n632), .ZN(new_n636));
  AOI211_X1 g450(.A(new_n431), .B(G902), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n430), .A2(new_n431), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n389), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n630), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n626), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT34), .B(G104), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  INV_X1    g458(.A(new_n389), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n437), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n646), .A2(new_n630), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n626), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT35), .B(G107), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  INV_X1    g464(.A(KEYINPUT95), .ZN(new_n651));
  AND3_X1   g465(.A1(new_n609), .A2(new_n610), .A3(KEYINPUT25), .ZN(new_n652));
  INV_X1    g466(.A(new_n614), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n652), .A2(new_n611), .A3(new_n653), .ZN(new_n654));
  OR3_X1    g468(.A1(new_n602), .A2(KEYINPUT36), .A3(new_n606), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n602), .B1(KEYINPUT36), .B2(new_n606), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n657), .A2(G902), .A3(new_n614), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n651), .B1(new_n654), .B2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n658), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n616), .A2(new_n660), .A3(KEYINPUT95), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n574), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n625), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n663), .A2(new_n664), .A3(new_n523), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT37), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(new_n594), .ZN(G12));
  NAND3_X1  g481(.A1(new_n628), .A2(new_n521), .A3(new_n629), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(G900), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n518), .A2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n514), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n645), .A2(new_n437), .A3(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n663), .A2(new_n328), .A3(new_n669), .A4(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G128), .ZN(G30));
  XOR2_X1   g490(.A(new_n673), .B(KEYINPUT39), .Z(new_n677));
  NOR2_X1   g491(.A1(new_n574), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(KEYINPUT96), .B(KEYINPUT40), .ZN(new_n679));
  OR2_X1    g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n512), .B(KEYINPUT38), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n682), .B1(new_n678), .B2(new_n679), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n389), .A2(new_n437), .A3(new_n521), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n321), .A2(KEYINPUT32), .A3(new_n322), .ZN(new_n685));
  AOI21_X1  g499(.A(KEYINPUT32), .B1(new_n321), .B2(new_n322), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n301), .B1(new_n296), .B2(new_n269), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n253), .B1(new_n288), .B2(new_n289), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n269), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n311), .B1(new_n690), .B2(new_n198), .ZN(new_n691));
  OAI21_X1  g505(.A(G472), .B1(new_n688), .B2(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n684), .B1(new_n687), .B2(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n680), .A2(new_n683), .A3(new_n662), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G143), .ZN(G45));
  NAND2_X1  g509(.A1(new_n635), .A2(new_n636), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n696), .A2(G478), .A3(new_n311), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n638), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n698), .A2(new_n389), .A3(new_n673), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n663), .A2(new_n328), .A3(new_n669), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G146), .ZN(G48));
  OR2_X1    g516(.A1(new_n560), .A2(new_n561), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n703), .A2(new_n573), .A3(new_n562), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n328), .A2(new_n620), .A3(new_n641), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(KEYINPUT41), .B(G113), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G15));
  NAND4_X1  g522(.A1(new_n328), .A2(new_n647), .A3(new_n705), .A4(new_n620), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G116), .ZN(G18));
  NOR2_X1   g524(.A1(new_n704), .A2(new_n438), .ZN(new_n711));
  INV_X1    g525(.A(new_n630), .ZN(new_n712));
  INV_X1    g526(.A(new_n662), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n711), .A2(new_n328), .A3(new_n712), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G119), .ZN(G21));
  AOI21_X1  g529(.A(new_n308), .B1(new_n689), .B2(new_n269), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n301), .B1(new_n716), .B2(new_n291), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n317), .A2(new_n320), .A3(new_n717), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n718), .A2(new_n322), .ZN(new_n719));
  XOR2_X1   g533(.A(KEYINPUT97), .B(G472), .Z(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n721), .B1(new_n321), .B2(new_n311), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n719), .A2(new_n722), .A3(new_n619), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n389), .A2(new_n437), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n668), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n723), .A2(new_n705), .A3(new_n520), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(KEYINPUT98), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G122), .ZN(G24));
  NOR3_X1   g542(.A1(new_n662), .A2(new_n719), .A3(new_n722), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n729), .A2(new_n669), .A3(new_n700), .A4(new_n705), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G125), .ZN(G27));
  INV_X1    g545(.A(KEYINPUT42), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n328), .A2(new_n620), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n567), .B1(new_n560), .B2(new_n561), .ZN(new_n734));
  OR2_X1    g548(.A1(new_n563), .A2(KEYINPUT99), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT99), .ZN(new_n736));
  OAI211_X1 g550(.A(G469), .B(new_n735), .C1(new_n565), .C2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n512), .ZN(new_n739));
  INV_X1    g553(.A(new_n521), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n572), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n738), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(KEYINPUT100), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT100), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n738), .A2(new_n744), .A3(new_n739), .A4(new_n741), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n733), .A2(new_n746), .A3(new_n700), .ZN(new_n747));
  AOI211_X1 g561(.A(new_n732), .B(new_n699), .C1(new_n743), .C2(new_n745), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n326), .A2(KEYINPUT101), .ZN(new_n749));
  AND4_X1   g563(.A1(new_n325), .A2(new_n749), .A3(new_n315), .A4(new_n327), .ZN(new_n750));
  OR2_X1    g564(.A1(new_n326), .A2(KEYINPUT101), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n619), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  AOI22_X1  g566(.A1(new_n732), .A2(new_n747), .B1(new_n748), .B2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n225), .ZN(G33));
  NAND3_X1  g568(.A1(new_n733), .A2(new_n746), .A3(new_n674), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G134), .ZN(G36));
  OR2_X1    g570(.A1(new_n389), .A2(KEYINPUT103), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n389), .A2(KEYINPUT103), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n698), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(KEYINPUT43), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n698), .A2(KEYINPUT102), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT43), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT102), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n697), .A2(new_n764), .A3(new_n638), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n762), .A2(new_n763), .A3(new_n645), .A4(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n761), .A2(new_n625), .A3(new_n713), .A4(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT44), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n512), .A2(new_n740), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n637), .A2(new_n639), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n771), .B1(new_n757), .B2(new_n758), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n766), .B1(new_n772), .B2(new_n763), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n774), .A2(KEYINPUT44), .A3(new_n625), .A4(new_n713), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n769), .A2(new_n770), .A3(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT104), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n677), .ZN(new_n779));
  OAI211_X1 g593(.A(KEYINPUT45), .B(new_n735), .C1(new_n565), .C2(new_n736), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n780), .B(G469), .C1(KEYINPUT45), .C2(new_n565), .ZN(new_n781));
  AOI21_X1  g595(.A(KEYINPUT46), .B1(new_n781), .B2(new_n568), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n782), .B1(new_n561), .B2(new_n560), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n781), .A2(KEYINPUT46), .A3(new_n568), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n572), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n769), .A2(new_n775), .A3(KEYINPUT104), .A4(new_n770), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n778), .A2(new_n779), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT105), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G137), .ZN(G39));
  INV_X1    g603(.A(KEYINPUT47), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n785), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n785), .A2(new_n790), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n770), .ZN(new_n794));
  NOR4_X1   g608(.A1(new_n328), .A2(new_n620), .A3(new_n699), .A4(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT106), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G140), .ZN(G42));
  INV_X1    g612(.A(KEYINPUT111), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n761), .A2(new_n799), .A3(new_n514), .A4(new_n766), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n514), .B(new_n766), .C1(new_n772), .C2(new_n763), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT111), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n704), .A2(new_n794), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n803), .A2(new_n752), .A3(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT48), .ZN(new_n806));
  INV_X1    g620(.A(G952), .ZN(new_n807));
  INV_X1    g621(.A(new_n723), .ZN(new_n808));
  AOI211_X1 g622(.A(new_n704), .B(new_n808), .C1(new_n800), .C2(new_n802), .ZN(new_n809));
  AOI211_X1 g623(.A(new_n807), .B(G953), .C1(new_n809), .C2(new_n669), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n325), .A2(new_n326), .A3(new_n692), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n811), .A2(new_n619), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n812), .A2(new_n514), .A3(new_n804), .ZN(new_n813));
  OR2_X1    g627(.A1(new_n813), .A2(new_n640), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n806), .A2(new_n810), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n803), .A2(new_n729), .A3(new_n804), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n813), .A2(new_n389), .A3(new_n698), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT50), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n803), .A2(new_n740), .A3(new_n705), .A4(new_n723), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n819), .B1(new_n820), .B2(new_n681), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n809), .A2(KEYINPUT50), .A3(new_n740), .A4(new_n682), .ZN(new_n822));
  AOI211_X1 g636(.A(new_n817), .B(new_n818), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT51), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n703), .A2(new_n562), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(KEYINPUT112), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n572), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n827), .B1(new_n791), .B2(new_n792), .ZN(new_n828));
  AOI211_X1 g642(.A(new_n808), .B(new_n794), .C1(new_n800), .C2(new_n802), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n824), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n815), .B1(new_n823), .B2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT107), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n832), .B1(new_n640), .B2(new_n522), .ZN(new_n833));
  AOI211_X1 g647(.A(new_n519), .B(new_n740), .C1(new_n510), .C2(new_n511), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n834), .A2(new_n437), .A3(new_n645), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n834), .A2(KEYINPUT107), .A3(new_n698), .A4(new_n389), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n833), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(new_n626), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n838), .A2(new_n621), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n706), .A2(new_n726), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n714), .A2(new_n709), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n839), .A2(new_n665), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n746), .A2(new_n700), .A3(new_n729), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n438), .B1(new_n672), .B2(new_n671), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n844), .A2(new_n663), .A3(new_n328), .A4(new_n770), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n755), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n842), .A2(new_n753), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT53), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n730), .A2(new_n675), .A3(new_n701), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n628), .A2(new_n573), .A3(new_n629), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n616), .A2(new_n660), .A3(new_n673), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n684), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n811), .A2(new_n852), .A3(new_n853), .A4(new_n738), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(KEYINPUT108), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT52), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n849), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n693), .A2(KEYINPUT108), .A3(new_n738), .A4(new_n852), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT108), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n854), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n730), .A2(new_n675), .A3(new_n701), .ZN(new_n862));
  OAI21_X1  g676(.A(KEYINPUT52), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT110), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n857), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n864), .B1(new_n857), .B2(new_n863), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n847), .B(new_n848), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n747), .A2(new_n732), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n748), .A2(new_n752), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(new_n846), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n714), .A2(new_n709), .A3(new_n706), .A4(new_n726), .ZN(new_n872));
  INV_X1    g686(.A(new_n665), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n870), .A2(new_n871), .A3(new_n839), .A4(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n856), .B1(new_n849), .B2(new_n855), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n861), .A2(new_n862), .A3(KEYINPUT52), .ZN(new_n877));
  OAI21_X1  g691(.A(KEYINPUT109), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT109), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n857), .A2(new_n863), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n875), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n867), .B1(new_n881), .B2(new_n848), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n818), .B1(new_n821), .B2(new_n822), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n827), .B(KEYINPUT113), .Z(new_n886));
  OAI21_X1  g700(.A(new_n829), .B1(new_n793), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n885), .A2(new_n887), .A3(new_n816), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n824), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n857), .A2(new_n863), .A3(new_n879), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n879), .B1(new_n857), .B2(new_n863), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n847), .B(new_n848), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(KEYINPUT110), .B1(new_n876), .B2(new_n877), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n857), .A2(new_n863), .A3(new_n864), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n875), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n892), .B(KEYINPUT54), .C1(new_n895), .C2(new_n848), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n831), .A2(new_n884), .A3(new_n889), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n807), .A2(new_n330), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n825), .B(KEYINPUT49), .Z(new_n900));
  NOR3_X1   g714(.A1(new_n681), .A2(new_n740), .A3(new_n572), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n900), .A2(new_n772), .A3(new_n812), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT114), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n899), .A2(KEYINPUT114), .A3(new_n902), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(G75));
  INV_X1    g721(.A(KEYINPUT56), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n847), .B1(new_n890), .B2(new_n891), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT53), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n910), .A2(G902), .A3(new_n867), .ZN(new_n911));
  INV_X1    g725(.A(G210), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n908), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n476), .A2(new_n478), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(new_n486), .Z(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT55), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n913), .A2(KEYINPUT115), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT115), .B1(new_n913), .B2(new_n916), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n911), .A2(KEYINPUT116), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT116), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n910), .A2(new_n920), .A3(G902), .A4(new_n867), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n508), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n916), .A2(KEYINPUT56), .ZN(new_n923));
  OAI22_X1  g737(.A1(new_n917), .A2(new_n918), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n330), .A2(G952), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT117), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n924), .A2(new_n926), .ZN(G51));
  AND2_X1   g741(.A1(new_n919), .A2(new_n921), .ZN(new_n928));
  OR2_X1    g742(.A1(new_n928), .A2(new_n781), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n910), .A2(KEYINPUT54), .A3(new_n867), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n884), .A2(KEYINPUT118), .A3(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT118), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n882), .A2(new_n932), .A3(new_n883), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n567), .B(KEYINPUT57), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n931), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n555), .A2(new_n559), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n925), .B1(new_n929), .B2(new_n937), .ZN(G54));
  INV_X1    g752(.A(KEYINPUT58), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n939), .B1(new_n919), .B2(new_n921), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n940), .A2(G475), .A3(new_n379), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n379), .B1(new_n940), .B2(G475), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n941), .A2(new_n942), .A3(new_n925), .ZN(G60));
  INV_X1    g757(.A(KEYINPUT119), .ZN(new_n944));
  NAND2_X1  g758(.A1(G478), .A2(G902), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT59), .Z(new_n946));
  AOI21_X1  g760(.A(new_n946), .B1(new_n884), .B2(new_n896), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n944), .B1(new_n947), .B2(new_n696), .ZN(new_n948));
  INV_X1    g762(.A(new_n946), .ZN(new_n949));
  INV_X1    g763(.A(new_n896), .ZN(new_n950));
  AOI21_X1  g764(.A(KEYINPUT54), .B1(new_n910), .B2(new_n867), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n696), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n952), .A2(KEYINPUT119), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n948), .A2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n926), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n931), .A2(new_n696), .A3(new_n933), .A4(new_n949), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(G63));
  XNOR2_X1  g772(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n613), .A2(new_n311), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n959), .B(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n910), .A2(new_n867), .A3(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n956), .B1(new_n962), .B2(new_n657), .ZN(new_n963));
  OAI21_X1  g777(.A(KEYINPUT61), .B1(new_n963), .B2(KEYINPUT121), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n607), .A2(new_n608), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n966), .B(new_n956), .C1(new_n657), .C2(new_n962), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n964), .B(new_n967), .ZN(G66));
  INV_X1    g782(.A(KEYINPUT123), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n842), .B(KEYINPUT122), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n330), .ZN(new_n971));
  INV_X1    g785(.A(G224), .ZN(new_n972));
  OAI21_X1  g786(.A(G953), .B1(new_n517), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n969), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n974), .B1(new_n969), .B2(new_n973), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n914), .B1(G898), .B2(new_n330), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT124), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n975), .B(new_n977), .ZN(G69));
  NAND2_X1  g792(.A1(new_n293), .A2(new_n295), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(new_n369), .ZN(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(G900), .A2(G953), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n785), .A2(new_n779), .A3(new_n725), .ZN(new_n983));
  INV_X1    g797(.A(new_n752), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n755), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n985), .B1(new_n793), .B2(new_n796), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n787), .A2(new_n849), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT125), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(KEYINPUT125), .B1(new_n787), .B2(new_n849), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n870), .B(new_n986), .C1(new_n989), .C2(new_n990), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n981), .B(new_n982), .C1(new_n991), .C2(G953), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n849), .A2(new_n694), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT62), .Z(new_n994));
  NAND2_X1  g808(.A1(new_n646), .A2(new_n640), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n733), .A2(new_n678), .A3(new_n770), .A4(new_n995), .ZN(new_n996));
  AND4_X1   g810(.A1(new_n787), .A2(new_n994), .A3(new_n797), .A4(new_n996), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n980), .B1(new_n997), .B2(G953), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n992), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n330), .B1(G227), .B2(G900), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1000), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n992), .A2(new_n1002), .A3(new_n998), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1001), .A2(new_n1003), .ZN(G72));
  XNOR2_X1  g818(.A(new_n987), .B(new_n988), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n302), .B(KEYINPUT126), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n1005), .A2(new_n870), .A3(new_n986), .A4(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n997), .A2(new_n688), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n970), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  OR2_X1    g823(.A1(new_n1006), .A2(new_n688), .ZN(new_n1010));
  NAND2_X1  g824(.A1(G472), .A2(G902), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1011), .B(KEYINPUT63), .ZN(new_n1012));
  AND2_X1   g826(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(new_n302), .ZN(new_n1014));
  NOR3_X1   g828(.A1(new_n1014), .A2(new_n688), .A3(new_n1012), .ZN(new_n1015));
  OAI211_X1 g829(.A(new_n892), .B(new_n1015), .C1(new_n895), .C2(new_n848), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1016), .ZN(new_n1017));
  NOR4_X1   g831(.A1(new_n1009), .A2(new_n925), .A3(new_n1013), .A4(new_n1017), .ZN(G57));
endmodule


