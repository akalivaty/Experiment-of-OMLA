//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 0 0 0 1 0 1 1 0 1 1 1 0 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 0 1 0 0 0 1 1 1 0 0 1 1 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:05 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n560, new_n562, new_n563, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n573, new_n574, new_n575,
    new_n576, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n636, new_n637,
    new_n640, new_n641, new_n643, new_n644, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1219, new_n1220, new_n1221;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT64), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT65), .Z(new_n451));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT66), .Z(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  AOI22_X1  g031(.A1(new_n451), .A2(G567), .B1(new_n453), .B2(G2106), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT67), .Z(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  OR2_X1    g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI22_X1  g037(.A1(new_n462), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g040(.A(G2105), .B1(new_n460), .B2(new_n461), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G137), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n464), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  OR2_X1    g045(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(G160));
  NAND2_X1  g047(.A1(new_n466), .A2(G136), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n464), .A2(G112), .ZN(new_n474));
  OAI21_X1  g049(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n475));
  AND2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  OAI21_X1  g052(.A(G2105), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g055(.A(KEYINPUT68), .B(G2105), .C1(new_n476), .C2(new_n477), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(G124), .ZN(new_n483));
  OAI221_X1 g058(.A(new_n473), .B1(new_n474), .B2(new_n475), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT69), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  OAI21_X1  g061(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT70), .ZN(new_n489));
  OAI21_X1  g064(.A(G2105), .B1(new_n489), .B2(G114), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(KEYINPUT70), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n488), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G126), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n493), .B1(new_n494), .B2(new_n478), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n466), .A2(G138), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n466), .A2(new_n498), .A3(G138), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n495), .B1(new_n497), .B2(new_n499), .ZN(G164));
  AND2_X1   g075(.A1(KEYINPUT6), .A2(G651), .ZN(new_n501));
  NOR2_X1   g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  OAI211_X1 g077(.A(G50), .B(G543), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  XNOR2_X1  g078(.A(new_n503), .B(KEYINPUT71), .ZN(new_n504));
  NAND2_X1  g079(.A1(G75), .A2(G543), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G62), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n505), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OR2_X1    g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  OR2_X1    g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n510), .A2(G651), .B1(new_n515), .B2(G88), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n504), .A2(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n519), .B1(new_n511), .B2(new_n512), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G51), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n513), .A2(new_n514), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n522), .A2(G63), .A3(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT72), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n521), .A2(KEYINPUT72), .A3(new_n523), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n515), .A2(G89), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n526), .A2(new_n527), .A3(new_n529), .A4(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  INV_X1    g107(.A(KEYINPUT73), .ZN(new_n533));
  INV_X1    g108(.A(G64), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n534), .B1(new_n513), .B2(new_n514), .ZN(new_n535));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n533), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  OAI211_X1 g113(.A(KEYINPUT73), .B(new_n536), .C1(new_n508), .C2(new_n534), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n538), .A2(G651), .A3(new_n539), .ZN(new_n540));
  XOR2_X1   g115(.A(KEYINPUT74), .B(G90), .Z(new_n541));
  AOI22_X1  g116(.A1(new_n515), .A2(new_n541), .B1(new_n520), .B2(G52), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(G171));
  XOR2_X1   g119(.A(KEYINPUT76), .B(G43), .Z(new_n545));
  NAND2_X1  g120(.A1(new_n520), .A2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(G81), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n502), .A2(new_n501), .B1(new_n506), .B2(new_n507), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT75), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n522), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G651), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(G68), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G56), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n508), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n556), .A2(KEYINPUT75), .A3(G651), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n549), .B1(new_n553), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n560));
  XOR2_X1   g135(.A(new_n560), .B(KEYINPUT77), .Z(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  AOI22_X1  g139(.A1(new_n522), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G91), .ZN(new_n566));
  OAI22_X1  g141(.A1(new_n565), .A2(new_n552), .B1(new_n566), .B2(new_n548), .ZN(new_n567));
  OAI211_X1 g142(.A(G53), .B(G543), .C1(new_n501), .C2(new_n502), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n568), .B(new_n569), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(G299));
  INV_X1    g147(.A(KEYINPUT78), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n540), .A2(new_n573), .A3(new_n542), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n573), .B1(new_n540), .B2(new_n542), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n575), .A2(new_n576), .ZN(G301));
  NAND2_X1  g152(.A1(new_n515), .A2(G87), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n522), .B2(G74), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n520), .A2(G49), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G288));
  INV_X1    g156(.A(KEYINPUT80), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n515), .A2(new_n582), .A3(G86), .ZN(new_n583));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT79), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n584), .B(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n587), .B1(new_n513), .B2(new_n514), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(G86), .ZN(new_n590));
  OAI21_X1  g165(.A(KEYINPUT80), .B1(new_n548), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n520), .A2(G48), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n583), .A2(new_n589), .A3(new_n591), .A4(new_n592), .ZN(G305));
  INV_X1    g168(.A(KEYINPUT82), .ZN(new_n594));
  INV_X1    g169(.A(G47), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(KEYINPUT81), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT81), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(G47), .ZN(new_n598));
  AND2_X1   g173(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n515), .A2(G85), .B1(new_n520), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G60), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n601), .B1(new_n513), .B2(new_n514), .ZN(new_n602));
  NAND2_X1  g177(.A1(G72), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(G651), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n594), .B1(new_n600), .B2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G85), .ZN(new_n607));
  OAI21_X1  g182(.A(G543), .B1(new_n501), .B2(new_n502), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n596), .A2(new_n598), .ZN(new_n609));
  OAI22_X1  g184(.A1(new_n548), .A2(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(G60), .B1(new_n506), .B2(new_n507), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n552), .B1(new_n611), .B2(new_n603), .ZN(new_n612));
  NOR3_X1   g187(.A1(new_n610), .A2(KEYINPUT82), .A3(new_n612), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n606), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(G290));
  NAND2_X1  g190(.A1(G79), .A2(G543), .ZN(new_n616));
  INV_X1    g191(.A(G66), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n508), .B2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT84), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g195(.A(KEYINPUT84), .B(new_n616), .C1(new_n508), .C2(new_n617), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n620), .A2(G651), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n520), .A2(G54), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n515), .A2(KEYINPUT10), .A3(G92), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT10), .ZN(new_n625));
  INV_X1    g200(.A(G92), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n548), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n622), .A2(new_n623), .A3(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(G868), .ZN(new_n630));
  AOI21_X1  g205(.A(KEYINPUT83), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(G301), .A2(G868), .ZN(new_n632));
  MUX2_X1   g207(.A(KEYINPUT83), .B(new_n631), .S(new_n632), .Z(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(G284));
  INV_X1    g209(.A(new_n633), .ZN(G321));
  NOR2_X1   g210(.A1(G286), .A2(new_n630), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n571), .B(KEYINPUT85), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n636), .B1(new_n637), .B2(new_n630), .ZN(G297));
  AOI21_X1  g213(.A(new_n636), .B1(new_n637), .B2(new_n630), .ZN(G280));
  INV_X1    g214(.A(new_n629), .ZN(new_n640));
  INV_X1    g215(.A(G559), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n640), .B1(new_n641), .B2(G860), .ZN(G148));
  OR2_X1    g217(.A1(new_n558), .A2(G868), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n629), .A2(G559), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n643), .B1(new_n644), .B2(new_n630), .ZN(G323));
  XNOR2_X1  g220(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g221(.A1(new_n462), .A2(new_n468), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT12), .Z(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT13), .Z(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(new_n482), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(G123), .ZN(new_n652));
  OAI21_X1  g227(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n653));
  INV_X1    g228(.A(G111), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n653), .B1(new_n654), .B2(G2105), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n655), .B1(G135), .B2(new_n466), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  AOI22_X1  g232(.A1(new_n650), .A2(G2100), .B1(G2096), .B2(new_n657), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n657), .A2(G2096), .ZN(new_n659));
  OAI211_X1 g234(.A(new_n658), .B(new_n659), .C1(G2100), .C2(new_n650), .ZN(G156));
  XNOR2_X1  g235(.A(KEYINPUT15), .B(G2435), .ZN(new_n661));
  INV_X1    g236(.A(G2438), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2427), .B(G2430), .Z(new_n664));
  OR2_X1    g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(KEYINPUT87), .B(KEYINPUT14), .Z(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n664), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT86), .B(KEYINPUT16), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G2451), .B(G2454), .Z(new_n671));
  XNOR2_X1  g246(.A(G2443), .B(G2446), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n670), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G1341), .B(G1348), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT88), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(G14), .ZN(new_n679));
  OR3_X1    g254(.A1(new_n674), .A2(KEYINPUT89), .A3(new_n677), .ZN(new_n680));
  OAI21_X1  g255(.A(KEYINPUT89), .B1(new_n674), .B2(new_n677), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n679), .B1(new_n680), .B2(new_n681), .ZN(G401));
  XNOR2_X1  g257(.A(G2072), .B(G2078), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT17), .Z(new_n684));
  XNOR2_X1  g259(.A(G2067), .B(G2678), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G2084), .B(G2090), .Z(new_n688));
  INV_X1    g263(.A(new_n683), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n688), .B1(new_n686), .B2(new_n689), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n687), .B1(KEYINPUT90), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(KEYINPUT90), .B2(new_n690), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n688), .A2(new_n685), .A3(new_n683), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT18), .Z(new_n694));
  NAND3_X1  g269(.A1(new_n684), .A2(new_n688), .A3(new_n686), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n692), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(G2096), .B(G2100), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(G227));
  XNOR2_X1  g273(.A(G1971), .B(G1976), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT19), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(G1956), .B(G2474), .Z(new_n702));
  XOR2_X1   g277(.A(G1961), .B(G1966), .Z(new_n703));
  AND2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT20), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n702), .A2(new_n703), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  MUX2_X1   g284(.A(new_n709), .B(new_n708), .S(new_n701), .Z(new_n710));
  NOR2_X1   g285(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n711), .B(new_n713), .ZN(new_n714));
  XOR2_X1   g289(.A(G1991), .B(G1996), .Z(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(G1981), .B(G1986), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n714), .A2(new_n716), .ZN(new_n719));
  AND3_X1   g294(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n718), .B1(new_n717), .B2(new_n719), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n720), .A2(new_n721), .ZN(G229));
  NAND2_X1  g297(.A1(new_n466), .A2(G139), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT93), .Z(new_n724));
  NAND3_X1  g299(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT25), .Z(new_n726));
  AOI22_X1  g301(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n726), .B1(new_n727), .B2(new_n464), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G29), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n730), .B2(G33), .ZN(new_n732));
  INV_X1    g307(.A(G2072), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT94), .ZN(new_n735));
  INV_X1    g310(.A(G16), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G21), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G168), .B2(new_n736), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G1966), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G28), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n741), .A2(KEYINPUT30), .ZN(new_n742));
  AOI21_X1  g317(.A(G29), .B1(new_n741), .B2(KEYINPUT30), .ZN(new_n743));
  OR2_X1    g318(.A1(KEYINPUT31), .A2(G11), .ZN(new_n744));
  NAND2_X1  g319(.A1(KEYINPUT31), .A2(G11), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n742), .A2(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n652), .A2(G29), .A3(new_n656), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT95), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n462), .A2(G141), .A3(new_n464), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT26), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n468), .A2(G105), .ZN(new_n754));
  AND3_X1   g329(.A1(new_n750), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n480), .A2(G129), .A3(new_n481), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n758), .A2(new_n730), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n730), .B2(G32), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT27), .B(G1996), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n749), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI221_X1 g337(.A(new_n762), .B1(new_n760), .B2(new_n761), .C1(new_n733), .C2(new_n732), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n730), .A2(G27), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G164), .B2(new_n730), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT96), .Z(new_n766));
  AND2_X1   g341(.A1(new_n766), .A2(G2078), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n766), .A2(G2078), .ZN(new_n768));
  NOR3_X1   g343(.A1(new_n763), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  AND2_X1   g344(.A1(KEYINPUT24), .A2(G34), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n730), .B1(KEYINPUT24), .B2(G34), .ZN(new_n771));
  OAI22_X1  g346(.A1(G160), .A2(new_n730), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G2084), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n738), .A2(G1966), .ZN(new_n774));
  AOI211_X1 g349(.A(new_n773), .B(new_n774), .C1(new_n748), .C2(new_n747), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n736), .A2(G5), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G171), .B2(new_n736), .ZN(new_n777));
  INV_X1    g352(.A(G1961), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n740), .A2(new_n769), .A3(new_n775), .A4(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT97), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n730), .A2(G25), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n651), .A2(G119), .ZN(new_n784));
  OAI21_X1  g359(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n785));
  INV_X1    g360(.A(G107), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n785), .B1(new_n786), .B2(G2105), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G131), .B2(new_n466), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n784), .A2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n783), .B1(new_n790), .B2(new_n730), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT35), .B(G1991), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(G1986), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n614), .A2(new_n736), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n736), .B2(G24), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n793), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n794), .B2(new_n796), .ZN(new_n798));
  NAND2_X1  g373(.A1(G166), .A2(G16), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G16), .B2(G22), .ZN(new_n800));
  INV_X1    g375(.A(G1971), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT32), .B(G1981), .Z(new_n802));
  AND2_X1   g377(.A1(new_n736), .A2(G6), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G305), .B2(G16), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n800), .A2(new_n801), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(new_n801), .B2(new_n800), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n736), .A2(G23), .ZN(new_n807));
  INV_X1    g382(.A(G288), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n807), .B1(new_n808), .B2(new_n736), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT33), .B(G1976), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n802), .B2(new_n804), .ZN(new_n812));
  OAI21_X1  g387(.A(KEYINPUT34), .B1(new_n806), .B2(new_n812), .ZN(new_n813));
  OR3_X1    g388(.A1(new_n806), .A2(KEYINPUT34), .A3(new_n812), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n798), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT36), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n780), .A2(new_n781), .ZN(new_n817));
  NOR2_X1   g392(.A1(G29), .A2(G35), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(G162), .B2(G29), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT29), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G2090), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n736), .A2(G19), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n558), .B2(new_n736), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(G1341), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n736), .A2(G4), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n640), .B2(new_n736), .ZN(new_n826));
  XOR2_X1   g401(.A(KEYINPUT91), .B(G1348), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT92), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n826), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n736), .A2(G20), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT23), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(new_n571), .B2(new_n736), .ZN(new_n832));
  INV_X1    g407(.A(G1956), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n730), .A2(G26), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT28), .Z(new_n836));
  NAND3_X1  g411(.A1(new_n480), .A2(G128), .A3(new_n481), .ZN(new_n837));
  OAI21_X1  g412(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n838));
  INV_X1    g413(.A(G116), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n838), .B1(new_n839), .B2(G2105), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(G140), .B2(new_n466), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n836), .B1(new_n842), .B2(G29), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(G2067), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n829), .A2(new_n834), .A3(new_n844), .ZN(new_n845));
  NOR3_X1   g420(.A1(new_n821), .A2(new_n824), .A3(new_n845), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n782), .A2(new_n816), .A3(new_n817), .A4(new_n846), .ZN(G150));
  INV_X1    g422(.A(G150), .ZN(G311));
  XOR2_X1   g423(.A(KEYINPUT98), .B(G93), .Z(new_n849));
  INV_X1    g424(.A(G55), .ZN(new_n850));
  OAI22_X1  g425(.A1(new_n548), .A2(new_n849), .B1(new_n608), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(G67), .B1(new_n506), .B2(new_n507), .ZN(new_n852));
  NAND2_X1  g427(.A1(G80), .A2(G543), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n552), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(G860), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT37), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n640), .A2(G559), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT38), .ZN(new_n860));
  INV_X1    g435(.A(new_n549), .ZN(new_n861));
  INV_X1    g436(.A(G67), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n862), .B1(new_n513), .B2(new_n514), .ZN(new_n863));
  INV_X1    g438(.A(new_n853), .ZN(new_n864));
  OAI21_X1  g439(.A(G651), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(KEYINPUT98), .B(G93), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n522), .B(new_n866), .C1(new_n502), .C2(new_n501), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n520), .A2(G55), .ZN(new_n868));
  NAND4_X1  g443(.A1(new_n865), .A2(new_n867), .A3(KEYINPUT99), .A4(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n557), .ZN(new_n870));
  AOI21_X1  g445(.A(KEYINPUT75), .B1(new_n556), .B2(G651), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n861), .B(new_n869), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT99), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT100), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n873), .B(new_n874), .C1(new_n851), .C2(new_n854), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n865), .A2(new_n868), .A3(new_n867), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n874), .B1(new_n877), .B2(new_n873), .ZN(new_n878));
  NOR3_X1   g453(.A1(new_n872), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(KEYINPUT100), .B1(new_n855), .B2(KEYINPUT99), .ZN(new_n880));
  AOI22_X1  g455(.A1(new_n880), .A2(new_n875), .B1(new_n558), .B2(new_n869), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n860), .B(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n884), .A2(KEYINPUT39), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n856), .B1(new_n884), .B2(KEYINPUT39), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n858), .B1(new_n885), .B2(new_n886), .ZN(G145));
  XOR2_X1   g462(.A(KEYINPUT104), .B(G37), .Z(new_n888));
  AND3_X1   g463(.A1(new_n480), .A2(G129), .A3(new_n481), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n750), .A2(new_n753), .A3(new_n754), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n837), .B(new_n841), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n842), .A2(new_n756), .A3(new_n755), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n891), .A2(new_n892), .A3(G164), .ZN(new_n893));
  AOI21_X1  g468(.A(G164), .B1(new_n891), .B2(new_n892), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n729), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT102), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI211_X1 g472(.A(KEYINPUT102), .B(new_n729), .C1(new_n893), .C2(new_n894), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n466), .A2(G142), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n464), .A2(G118), .ZN(new_n901));
  OAI21_X1  g476(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n902));
  INV_X1    g477(.A(G130), .ZN(new_n903));
  OAI221_X1 g478(.A(new_n900), .B1(new_n901), .B2(new_n902), .C1(new_n482), .C2(new_n903), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n904), .A2(new_n648), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(new_n648), .ZN(new_n906));
  OR3_X1    g481(.A1(new_n905), .A2(new_n906), .A3(new_n790), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n790), .B1(new_n905), .B2(new_n906), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n891), .A2(new_n892), .ZN(new_n911));
  INV_X1    g486(.A(G164), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n729), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n891), .A2(new_n892), .A3(G164), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT103), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n913), .A2(new_n914), .A3(new_n918), .A4(new_n915), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n899), .A2(new_n910), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n910), .B1(new_n899), .B2(new_n920), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT101), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n657), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n652), .A2(KEYINPUT101), .A3(new_n656), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(G160), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n924), .A2(new_n471), .A3(new_n925), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n927), .A2(new_n485), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n485), .B1(new_n927), .B2(new_n928), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n921), .A2(new_n922), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n931), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n899), .A2(new_n920), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(new_n909), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n899), .A2(new_n910), .A3(new_n920), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n888), .B1(new_n932), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT105), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n931), .B1(new_n921), .B2(new_n922), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n935), .A2(new_n933), .A3(new_n936), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n943), .A2(KEYINPUT105), .A3(new_n888), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n940), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n945), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g521(.A1(new_n877), .A2(new_n630), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT82), .B1(new_n610), .B2(new_n612), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n515), .A2(G85), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n520), .A2(new_n599), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n949), .A2(new_n605), .A3(new_n594), .A4(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n948), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n952), .B1(new_n948), .B2(new_n951), .ZN(new_n954));
  OAI21_X1  g529(.A(G288), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AND2_X1   g530(.A1(G303), .A2(G305), .ZN(new_n956));
  NOR2_X1   g531(.A1(G303), .A2(G305), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT107), .B1(new_n606), .B2(new_n613), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n948), .A2(new_n951), .A3(new_n952), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n959), .A2(new_n808), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n955), .A2(new_n958), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT109), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT109), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n955), .A2(new_n958), .A3(new_n961), .A4(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n955), .A2(new_n961), .ZN(new_n967));
  INV_X1    g542(.A(new_n958), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n967), .A2(KEYINPUT108), .A3(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT108), .B1(new_n967), .B2(new_n968), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n966), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT110), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n972), .B1(new_n973), .B2(KEYINPUT42), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(KEYINPUT42), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n974), .B(new_n975), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n628), .A2(new_n623), .ZN(new_n977));
  NAND3_X1  g552(.A1(G299), .A2(new_n977), .A3(new_n622), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n629), .A2(KEYINPUT106), .A3(new_n571), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT106), .B1(new_n629), .B2(new_n571), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT41), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n981), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT41), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n983), .A2(new_n984), .A3(new_n978), .A4(new_n979), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n982), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n983), .A2(new_n978), .A3(new_n979), .ZN(new_n988));
  XOR2_X1   g563(.A(new_n882), .B(new_n644), .Z(new_n989));
  MUX2_X1   g564(.A(new_n987), .B(new_n988), .S(new_n989), .Z(new_n990));
  XNOR2_X1  g565(.A(new_n976), .B(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n947), .B1(new_n991), .B2(new_n630), .ZN(G295));
  OAI21_X1  g567(.A(new_n947), .B1(new_n991), .B2(new_n630), .ZN(G331));
  XNOR2_X1  g568(.A(KEYINPUT111), .B(KEYINPUT43), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(G37), .ZN(new_n996));
  OAI21_X1  g571(.A(G168), .B1(new_n575), .B2(new_n576), .ZN(new_n997));
  NAND2_X1  g572(.A1(G286), .A2(new_n543), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n997), .B(new_n998), .C1(new_n879), .C2(new_n881), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n880), .A2(new_n558), .A3(new_n869), .A4(new_n875), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n872), .B1(new_n876), .B2(new_n878), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n543), .A2(KEYINPUT78), .ZN(new_n1002));
  AOI21_X1  g577(.A(G286), .B1(new_n1002), .B2(new_n574), .ZN(new_n1003));
  INV_X1    g578(.A(new_n998), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n1000), .B(new_n1001), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n999), .A2(new_n1005), .A3(new_n988), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n999), .A2(new_n1005), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1006), .B1(new_n987), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT112), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n966), .B(new_n1009), .C1(new_n970), .C2(new_n971), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n996), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n999), .A2(new_n1005), .A3(new_n988), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n999), .A2(new_n1005), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1012), .B1(new_n1013), .B2(new_n986), .ZN(new_n1014));
  INV_X1    g589(.A(new_n971), .ZN(new_n1015));
  AOI22_X1  g590(.A1(new_n1015), .A2(new_n969), .B1(new_n963), .B2(new_n965), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1014), .B1(new_n1009), .B2(new_n1016), .ZN(new_n1017));
  OR2_X1    g592(.A1(new_n1011), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n888), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1008), .A2(new_n1016), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1014), .A2(new_n972), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1019), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1022), .A2(KEYINPUT114), .ZN(new_n1023));
  OAI21_X1  g598(.A(KEYINPUT43), .B1(new_n1022), .B2(KEYINPUT114), .ZN(new_n1024));
  OAI221_X1 g599(.A(KEYINPUT44), .B1(new_n995), .B2(new_n1018), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT113), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n995), .B1(new_n1011), .B2(new_n1017), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n1014), .A2(new_n972), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1014), .A2(new_n972), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n888), .B(new_n994), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT44), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1026), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  AOI211_X1 g608(.A(KEYINPUT113), .B(KEYINPUT44), .C1(new_n1027), .C2(new_n1030), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1025), .B1(new_n1033), .B2(new_n1034), .ZN(G397));
  INV_X1    g610(.A(G40), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n471), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT45), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1039), .B1(G164), .B2(G1384), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(G1996), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g618(.A(new_n1043), .B(KEYINPUT46), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1041), .ZN(new_n1045));
  XOR2_X1   g620(.A(new_n842), .B(G2067), .Z(new_n1046));
  AND2_X1   g621(.A1(new_n1046), .A2(new_n758), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1044), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n1048), .B(KEYINPUT47), .ZN(new_n1049));
  XNOR2_X1  g624(.A(new_n757), .B(new_n1042), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1046), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g627(.A(new_n789), .B(new_n792), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1045), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT48), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n614), .A2(new_n794), .ZN(new_n1056));
  OR2_X1    g631(.A1(new_n1056), .A2(KEYINPUT115), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(KEYINPUT115), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(new_n1041), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1054), .B1(new_n1055), .B2(new_n1059), .ZN(new_n1060));
  OR2_X1    g635(.A1(new_n1059), .A2(new_n1055), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n790), .A2(new_n792), .ZN(new_n1062));
  OAI22_X1  g637(.A1(new_n1051), .A2(new_n1062), .B1(G2067), .B2(new_n842), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1060), .A2(new_n1061), .B1(new_n1041), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1049), .A2(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g640(.A(new_n1065), .B(KEYINPUT126), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n1067));
  NOR2_X1   g642(.A1(G164), .A2(G1384), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT50), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(new_n1071), .A3(new_n1037), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1067), .B1(new_n1072), .B2(G2084), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n1037), .A2(new_n1071), .ZN(new_n1074));
  INV_X1    g649(.A(G2084), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1074), .A2(KEYINPUT120), .A3(new_n1075), .A4(new_n1070), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1068), .A2(KEYINPUT45), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1077), .A2(new_n1040), .A3(new_n1037), .ZN(new_n1078));
  INV_X1    g653(.A(G1966), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1073), .A2(new_n1076), .A3(G168), .A4(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT51), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1081), .A2(new_n1082), .A3(G8), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1073), .A2(new_n1076), .A3(new_n1080), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(G286), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1086), .A2(G8), .A3(new_n1081), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1084), .B1(new_n1087), .B2(KEYINPUT51), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT62), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT125), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  AND2_X1   g665(.A1(new_n1085), .A2(G286), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1081), .A2(G8), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT51), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n1083), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT125), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1094), .A2(new_n1095), .A3(KEYINPUT62), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1078), .A2(KEYINPUT117), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT117), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1077), .A2(new_n1040), .A3(new_n1098), .A4(new_n1037), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1097), .A2(new_n801), .A3(new_n1099), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n1072), .A2(G2090), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(G8), .ZN(new_n1103));
  NAND2_X1  g678(.A1(G303), .A2(G8), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n1104), .B(KEYINPUT55), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  OR2_X1    g681(.A1(G305), .A2(G1981), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n589), .B(new_n592), .C1(new_n590), .C2(new_n548), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(G1981), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT49), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1110), .A2(KEYINPUT119), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(G8), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1113), .B1(new_n1037), .B2(new_n1068), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1111), .A2(KEYINPUT119), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1107), .A2(new_n1109), .A3(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1112), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n808), .A2(G1976), .ZN(new_n1118));
  INV_X1    g693(.A(G1976), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT52), .B1(G288), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1114), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1117), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT52), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(KEYINPUT118), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT118), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1123), .A2(new_n1126), .A3(KEYINPUT52), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1122), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1106), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1078), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT53), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1131), .A2(G2078), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n1130), .A2(new_n1132), .B1(new_n1072), .B2(new_n778), .ZN(new_n1133));
  AOI21_X1  g708(.A(G2078), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1133), .B1(new_n1134), .B2(KEYINPUT53), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1135), .B1(new_n576), .B2(new_n575), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1105), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1102), .A2(G8), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  NOR3_X1   g714(.A1(new_n1129), .A2(new_n1136), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1090), .A2(new_n1096), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1117), .A2(new_n1119), .A3(new_n808), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(new_n1107), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(new_n1114), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1122), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1145), .B1(new_n1148), .B2(new_n1138), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1148), .B1(new_n1105), .B2(new_n1103), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT63), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(KEYINPUT121), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n1085), .A2(G8), .A3(G168), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1150), .A2(new_n1138), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1106), .A2(new_n1138), .A3(new_n1128), .A4(new_n1153), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1155), .A2(KEYINPUT121), .A3(new_n1151), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1149), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n571), .A2(KEYINPUT122), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n1158), .B(KEYINPUT57), .ZN(new_n1159));
  XNOR2_X1  g734(.A(KEYINPUT56), .B(G2072), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1130), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1072), .A2(new_n833), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1159), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1037), .A2(new_n1068), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1164), .A2(G2067), .ZN(new_n1165));
  INV_X1    g740(.A(G1348), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1165), .B1(new_n1166), .B2(new_n1072), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1167), .A2(new_n629), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1161), .A2(new_n1159), .A3(new_n1162), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1163), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1169), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1171), .B1(new_n1172), .B2(new_n1163), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1163), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1174), .A2(KEYINPUT61), .A3(new_n1169), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n640), .A2(KEYINPUT60), .ZN(new_n1177));
  XOR2_X1   g752(.A(new_n1177), .B(KEYINPUT123), .Z(new_n1178));
  INV_X1    g753(.A(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1167), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n640), .A2(KEYINPUT60), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1179), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  OAI211_X1 g757(.A(new_n1178), .B(new_n1167), .C1(KEYINPUT60), .C2(new_n640), .ZN(new_n1183));
  XOR2_X1   g758(.A(KEYINPUT58), .B(G1341), .Z(new_n1184));
  NAND2_X1  g759(.A1(new_n1164), .A2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1185), .B1(new_n1078), .B2(G1996), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1186), .A2(new_n558), .ZN(new_n1187));
  AND2_X1   g762(.A1(new_n1187), .A2(KEYINPUT59), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1187), .A2(KEYINPUT59), .ZN(new_n1189));
  OAI211_X1 g764(.A(new_n1182), .B(new_n1183), .C1(new_n1188), .C2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1170), .B1(new_n1176), .B2(new_n1190), .ZN(new_n1191));
  AND2_X1   g766(.A1(new_n1077), .A2(new_n1040), .ZN(new_n1192));
  XOR2_X1   g767(.A(new_n470), .B(KEYINPUT124), .Z(new_n1193));
  NAND2_X1  g768(.A1(new_n1132), .A2(G40), .ZN(new_n1194));
  NOR3_X1   g769(.A1(new_n1193), .A2(new_n465), .A3(new_n1194), .ZN(new_n1195));
  AOI22_X1  g770(.A1(new_n1192), .A2(new_n1195), .B1(new_n1072), .B2(new_n778), .ZN(new_n1196));
  OAI211_X1 g771(.A(G301), .B(new_n1196), .C1(new_n1134), .C2(KEYINPUT53), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1136), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT54), .ZN(new_n1199));
  OAI211_X1 g774(.A(G301), .B(new_n1133), .C1(new_n1134), .C2(KEYINPUT53), .ZN(new_n1200));
  AND2_X1   g775(.A1(new_n1200), .A2(KEYINPUT54), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1196), .B1(new_n1134), .B2(KEYINPUT53), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1202), .A2(G171), .ZN(new_n1203));
  AOI22_X1  g778(.A1(new_n1198), .A2(new_n1199), .B1(new_n1201), .B2(new_n1203), .ZN(new_n1204));
  NOR2_X1   g779(.A1(new_n1129), .A2(new_n1139), .ZN(new_n1205));
  NAND4_X1  g780(.A1(new_n1191), .A2(new_n1204), .A3(new_n1094), .A4(new_n1205), .ZN(new_n1206));
  AND3_X1   g781(.A1(new_n1142), .A2(new_n1157), .A3(new_n1206), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1041), .A2(G1986), .A3(G290), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1059), .A2(new_n1208), .ZN(new_n1209));
  XOR2_X1   g784(.A(new_n1209), .B(KEYINPUT116), .Z(new_n1210));
  OR2_X1    g785(.A1(new_n1210), .A2(new_n1054), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1066), .B1(new_n1207), .B2(new_n1211), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g787(.A1(G227), .A2(new_n458), .ZN(new_n1214));
  NOR3_X1   g788(.A1(G229), .A2(G401), .A3(new_n1214), .ZN(new_n1215));
  AOI21_X1  g789(.A(KEYINPUT105), .B1(new_n943), .B2(new_n888), .ZN(new_n1216));
  AOI211_X1 g790(.A(new_n939), .B(new_n1019), .C1(new_n941), .C2(new_n942), .ZN(new_n1217));
  OAI211_X1 g791(.A(new_n1031), .B(new_n1215), .C1(new_n1216), .C2(new_n1217), .ZN(G225));
  INV_X1    g792(.A(KEYINPUT127), .ZN(new_n1219));
  NAND2_X1  g793(.A1(G225), .A2(new_n1219), .ZN(new_n1220));
  NAND4_X1  g794(.A1(new_n945), .A2(KEYINPUT127), .A3(new_n1031), .A4(new_n1215), .ZN(new_n1221));
  AND2_X1   g795(.A1(new_n1220), .A2(new_n1221), .ZN(G308));
endmodule


