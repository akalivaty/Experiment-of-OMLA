//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 0 0 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 0 0 1 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n769, new_n770, new_n772,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n850, new_n851, new_n852, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968;
  INV_X1    g000(.A(KEYINPUT15), .ZN(new_n202));
  INV_X1    g001(.A(G43gat), .ZN(new_n203));
  INV_X1    g002(.A(G50gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G43gat), .A2(G50gat), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n202), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n210));
  INV_X1    g009(.A(G36gat), .ZN(new_n211));
  AND3_X1   g010(.A1(new_n210), .A2(KEYINPUT89), .A3(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(KEYINPUT89), .B1(new_n210), .B2(new_n211), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n209), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT90), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g015(.A1(new_n214), .A2(new_n215), .B1(G29gat), .B2(G36gat), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n208), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n207), .B1(G29gat), .B2(G36gat), .ZN(new_n219));
  XOR2_X1   g018(.A(KEYINPUT91), .B(G43gat), .Z(new_n220));
  OAI211_X1 g019(.A(new_n202), .B(new_n206), .C1(new_n220), .C2(G50gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT14), .ZN(new_n222));
  INV_X1    g021(.A(G29gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(new_n223), .A3(new_n211), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(new_n209), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n225), .A2(KEYINPUT92), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n225), .A2(KEYINPUT92), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n219), .B(new_n221), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n218), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G85gat), .A2(G92gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n232), .B(KEYINPUT7), .ZN(new_n233));
  NAND2_X1  g032(.A1(G99gat), .A2(G106gat), .ZN(new_n234));
  INV_X1    g033(.A(G85gat), .ZN(new_n235));
  INV_X1    g034(.A(G92gat), .ZN(new_n236));
  AOI22_X1  g035(.A1(KEYINPUT8), .A2(new_n234), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n233), .A2(new_n237), .ZN(new_n238));
  XOR2_X1   g037(.A(G99gat), .B(G106gat), .Z(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n239), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n241), .A2(new_n233), .A3(new_n237), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT100), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n240), .A2(KEYINPUT100), .A3(new_n242), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AND2_X1   g046(.A1(G232gat), .A2(G233gat), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n231), .A2(new_n247), .B1(KEYINPUT41), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT17), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n231), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n247), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT94), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n254), .B1(new_n230), .B2(KEYINPUT17), .ZN(new_n255));
  NOR4_X1   g054(.A1(new_n218), .A2(new_n229), .A3(KEYINPUT94), .A4(new_n250), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n249), .B1(new_n253), .B2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G190gat), .B(G218gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n259), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n261), .B(new_n249), .C1(new_n253), .C2(new_n257), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT101), .ZN(new_n264));
  AND2_X1   g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT99), .B(G134gat), .ZN(new_n266));
  INV_X1    g065(.A(G162gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n248), .A2(KEYINPUT41), .ZN(new_n269));
  XOR2_X1   g068(.A(new_n268), .B(new_n269), .Z(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n263), .B1(new_n265), .B2(new_n271), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n260), .A2(KEYINPUT101), .A3(new_n262), .A4(new_n270), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  XOR2_X1   g074(.A(G57gat), .B(G64gat), .Z(new_n276));
  NAND2_X1  g075(.A1(G71gat), .A2(G78gat), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT9), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g079(.A1(G71gat), .A2(G78gat), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT96), .ZN(new_n283));
  AOI22_X1  g082(.A1(new_n277), .A2(new_n282), .B1(new_n279), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n280), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n277), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n286), .A2(new_n281), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n276), .B(new_n279), .C1(new_n287), .C2(new_n283), .ZN(new_n288));
  AND2_X1   g087(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT97), .B(KEYINPUT21), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G231gat), .A2(G233gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n293), .B(G127gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(G183gat), .B(G211gat), .ZN(new_n295));
  XOR2_X1   g094(.A(new_n294), .B(new_n295), .Z(new_n296));
  XNOR2_X1  g095(.A(G15gat), .B(G22gat), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT93), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n299), .B(G8gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT16), .ZN(new_n301));
  AOI21_X1  g100(.A(G1gat), .B1(new_n297), .B2(new_n301), .ZN(new_n302));
  XOR2_X1   g101(.A(new_n300), .B(new_n302), .Z(new_n303));
  INV_X1    g102(.A(KEYINPUT21), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n303), .B1(new_n304), .B2(new_n289), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n305), .B(KEYINPUT98), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n307));
  INV_X1    g106(.A(G155gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n307), .B(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n306), .B(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n296), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n294), .B(new_n295), .ZN(new_n312));
  OR2_X1    g111(.A1(new_n306), .A2(new_n309), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n306), .A2(new_n309), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  AND2_X1   g114(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n275), .A2(KEYINPUT102), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT102), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n319), .B1(new_n316), .B2(new_n274), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n285), .A2(new_n288), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n243), .B(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT10), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n289), .A2(new_n324), .ZN(new_n325));
  AOI22_X1  g124(.A1(new_n323), .A2(new_n324), .B1(new_n247), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(G230gat), .A2(G233gat), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  OR2_X1    g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  OR2_X1    g128(.A1(new_n323), .A2(new_n327), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G120gat), .B(G148gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(G176gat), .B(G204gat), .ZN(new_n333));
  XOR2_X1   g132(.A(new_n332), .B(new_n333), .Z(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n329), .A2(new_n330), .A3(new_n334), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n321), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n251), .B(new_n303), .C1(new_n255), .C2(new_n256), .ZN(new_n341));
  NAND2_X1  g140(.A1(G229gat), .A2(G233gat), .ZN(new_n342));
  OR2_X1    g141(.A1(new_n303), .A2(new_n230), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT18), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n341), .A2(KEYINPUT18), .A3(new_n342), .A4(new_n343), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n303), .B(new_n230), .ZN(new_n348));
  XOR2_X1   g147(.A(new_n342), .B(KEYINPUT13), .Z(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n346), .A2(new_n347), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT88), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G113gat), .B(G141gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(KEYINPUT87), .B(G197gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n354), .B(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT11), .B(G169gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  XOR2_X1   g157(.A(new_n358), .B(KEYINPUT12), .Z(new_n359));
  NAND2_X1  g158(.A1(new_n353), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n359), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n351), .A2(new_n352), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT84), .ZN(new_n365));
  AND2_X1   g164(.A1(G155gat), .A2(G162gat), .ZN(new_n366));
  NOR2_X1   g165(.A1(G155gat), .A2(G162gat), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G141gat), .B(G148gat), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT2), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n370), .B1(G155gat), .B2(G162gat), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n368), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(G141gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(G148gat), .ZN(new_n374));
  INV_X1    g173(.A(G148gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(G141gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G155gat), .B(G162gat), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT2), .B1(new_n308), .B2(new_n267), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n372), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(G134gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(G127gat), .ZN(new_n384));
  INV_X1    g183(.A(G127gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(G134gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G113gat), .B(G120gat), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n387), .B1(new_n388), .B2(KEYINPUT1), .ZN(new_n389));
  INV_X1    g188(.A(G120gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(G113gat), .ZN(new_n391));
  INV_X1    g190(.A(G113gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(G120gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(G127gat), .B(G134gat), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT1), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  AND2_X1   g196(.A1(new_n389), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT4), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n382), .A2(new_n398), .A3(KEYINPUT78), .A4(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT78), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n372), .A2(new_n389), .A3(new_n380), .A4(new_n397), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n401), .B1(new_n402), .B2(KEYINPUT4), .ZN(new_n403));
  AND3_X1   g202(.A1(new_n402), .A2(KEYINPUT79), .A3(KEYINPUT4), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT79), .B1(new_n402), .B2(KEYINPUT4), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n400), .B(new_n403), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT5), .ZN(new_n407));
  NAND2_X1  g206(.A1(G225gat), .A2(G233gat), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n381), .A2(KEYINPUT3), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT3), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n372), .A2(new_n380), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n389), .A2(new_n397), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n409), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n406), .A2(new_n407), .A3(new_n408), .A4(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT77), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n381), .A2(new_n412), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n416), .A2(KEYINPUT76), .A3(new_n402), .ZN(new_n417));
  INV_X1    g216(.A(new_n408), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT76), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n381), .A2(new_n412), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n417), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n421), .A2(KEYINPUT5), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n399), .B1(new_n382), .B2(new_n398), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n402), .A2(KEYINPUT4), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n413), .B(new_n408), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n415), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n425), .A2(KEYINPUT5), .A3(new_n421), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n427), .A2(KEYINPUT77), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n414), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  XOR2_X1   g228(.A(G1gat), .B(G29gat), .Z(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(KEYINPUT0), .ZN(new_n431));
  XNOR2_X1  g230(.A(G57gat), .B(G85gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n429), .A2(KEYINPUT6), .A3(new_n434), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n433), .B(new_n414), .C1(new_n426), .C2(new_n428), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT6), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n433), .B(KEYINPUT81), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n422), .A2(new_n415), .A3(new_n425), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n427), .A2(KEYINPUT77), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n439), .B1(new_n442), .B2(new_n414), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n435), .B1(new_n438), .B2(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(G211gat), .B(G218gat), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT71), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n448));
  OR2_X1    g247(.A1(G197gat), .A2(G204gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(G197gat), .A2(G204gat), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n447), .B(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(G226gat), .ZN(new_n453));
  INV_X1    g252(.A(G233gat), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT25), .ZN(new_n456));
  NOR2_X1   g255(.A1(G183gat), .A2(G190gat), .ZN(new_n457));
  NAND2_X1  g256(.A1(G183gat), .A2(G190gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT24), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT24), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n460), .A2(G183gat), .A3(G190gat), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n457), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(G169gat), .ZN(new_n463));
  INV_X1    g262(.A(G176gat), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT23), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT23), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n466), .B1(G169gat), .B2(G176gat), .ZN(new_n467));
  NAND2_X1  g266(.A1(G169gat), .A2(G176gat), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n456), .B1(new_n462), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT64), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI211_X1 g271(.A(KEYINPUT64), .B(new_n456), .C1(new_n462), .C2(new_n469), .ZN(new_n473));
  XNOR2_X1  g272(.A(KEYINPUT65), .B(G183gat), .ZN(new_n474));
  INV_X1    g273(.A(G190gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n461), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n469), .A2(new_n456), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n472), .A2(new_n473), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n463), .A2(new_n464), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT26), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n458), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT26), .B1(new_n463), .B2(new_n464), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n484), .B1(new_n468), .B2(new_n485), .ZN(new_n486));
  OR2_X1    g285(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT27), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n487), .B1(new_n474), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT28), .B1(new_n489), .B2(new_n475), .ZN(new_n490));
  XOR2_X1   g289(.A(KEYINPUT27), .B(G183gat), .Z(new_n491));
  INV_X1    g290(.A(KEYINPUT28), .ZN(new_n492));
  NOR3_X1   g291(.A1(new_n491), .A2(new_n492), .A3(G190gat), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n486), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n481), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(KEYINPUT72), .B(KEYINPUT29), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n455), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AOI211_X1 g296(.A(new_n453), .B(new_n454), .C1(new_n481), .C2(new_n494), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n452), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n495), .A2(new_n455), .ZN(new_n500));
  INV_X1    g299(.A(new_n452), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT29), .B1(new_n481), .B2(new_n494), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n500), .B(new_n501), .C1(new_n455), .C2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n499), .A2(KEYINPUT37), .A3(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n501), .B1(new_n497), .B2(new_n498), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT37), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n500), .B(new_n452), .C1(new_n455), .C2(new_n502), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(G8gat), .B(G36gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(G64gat), .B(G92gat), .ZN(new_n510));
  XOR2_X1   g309(.A(new_n509), .B(new_n510), .Z(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(KEYINPUT73), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n512), .A2(KEYINPUT38), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n504), .A2(new_n508), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n505), .A2(new_n511), .A3(new_n507), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT75), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n505), .A2(KEYINPUT75), .A3(new_n511), .A4(new_n507), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n514), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n365), .B1(new_n444), .B2(new_n519), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n514), .A2(new_n517), .A3(new_n518), .ZN(new_n521));
  INV_X1    g320(.A(new_n439), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n429), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n523), .A2(new_n437), .A3(new_n436), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n521), .A2(new_n524), .A3(KEYINPUT84), .A4(new_n435), .ZN(new_n525));
  INV_X1    g324(.A(new_n505), .ZN(new_n526));
  INV_X1    g325(.A(new_n507), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT37), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n511), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(new_n529), .A3(new_n508), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT38), .ZN(new_n531));
  AND3_X1   g330(.A1(new_n520), .A2(new_n525), .A3(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G78gat), .B(G106gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(new_n204), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(G22gat), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n452), .B1(new_n411), .B2(new_n496), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n537), .B1(G228gat), .B2(G233gat), .ZN(new_n538));
  AND2_X1   g337(.A1(new_n452), .A2(new_n496), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n381), .B1(new_n539), .B2(KEYINPUT3), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT29), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n452), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n382), .B1(new_n543), .B2(new_n410), .ZN(new_n544));
  OAI211_X1 g343(.A(G228gat), .B(G233gat), .C1(new_n544), .C2(new_n537), .ZN(new_n545));
  XNOR2_X1  g344(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n541), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n547), .B1(new_n541), .B2(new_n545), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n536), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n550), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n552), .A2(new_n535), .A3(new_n548), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  AOI211_X1 g354(.A(KEYINPUT39), .B(new_n408), .C1(new_n406), .C2(new_n413), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT82), .B1(new_n556), .B2(new_n522), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n408), .B1(new_n406), .B2(new_n413), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT39), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT82), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n560), .A2(new_n561), .A3(new_n439), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n557), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n558), .A2(new_n559), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n418), .B1(new_n417), .B2(new_n420), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT83), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT40), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI22_X1  g369(.A1(new_n557), .A2(new_n562), .B1(new_n566), .B2(new_n564), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(KEYINPUT40), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n570), .A2(new_n523), .A3(new_n572), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n505), .A2(KEYINPUT30), .A3(new_n511), .A4(new_n507), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT74), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT30), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n517), .A2(new_n577), .A3(new_n518), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n526), .A2(new_n527), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n579), .A2(new_n512), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n576), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n555), .B1(new_n573), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(KEYINPUT85), .B1(new_n532), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT70), .ZN(new_n585));
  AND3_X1   g384(.A1(new_n481), .A2(new_n398), .A3(new_n494), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n398), .B1(new_n481), .B2(new_n494), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT67), .ZN(new_n589));
  NAND2_X1  g388(.A1(G227gat), .A2(G233gat), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n495), .A2(new_n412), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n481), .A2(new_n398), .A3(new_n494), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n592), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(KEYINPUT67), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT34), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT34), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n591), .A2(new_n595), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n590), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n601), .B1(new_n586), .B2(new_n587), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT32), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT33), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G71gat), .B(G99gat), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT66), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(G15gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n606), .B(KEYINPUT66), .ZN(new_n610));
  INV_X1    g409(.A(G15gat), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AND3_X1   g411(.A1(new_n609), .A2(new_n612), .A3(G43gat), .ZN(new_n613));
  AOI21_X1  g412(.A(G43gat), .B1(new_n609), .B2(new_n612), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n603), .A2(new_n605), .A3(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT68), .ZN(new_n617));
  INV_X1    g416(.A(new_n615), .ZN(new_n618));
  OAI211_X1 g417(.A(new_n602), .B(KEYINPUT32), .C1(new_n618), .C2(new_n604), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n616), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n600), .A2(new_n620), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n616), .A2(new_n617), .A3(new_n619), .ZN(new_n622));
  AND3_X1   g421(.A1(new_n591), .A2(new_n595), .A3(new_n598), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n598), .B1(new_n591), .B2(new_n595), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n590), .B1(new_n592), .B2(new_n593), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n615), .B1(new_n627), .B2(KEYINPUT33), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT32), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n619), .ZN(new_n632));
  OAI21_X1  g431(.A(KEYINPUT68), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n621), .B1(new_n626), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT36), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n585), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n633), .A2(new_n620), .A3(new_n600), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n625), .ZN(new_n638));
  AND4_X1   g437(.A1(new_n585), .A2(new_n637), .A3(new_n635), .A4(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT69), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n637), .A2(new_n638), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n640), .B1(new_n641), .B2(KEYINPUT36), .ZN(new_n642));
  AOI211_X1 g441(.A(KEYINPUT69), .B(new_n635), .C1(new_n637), .C2(new_n638), .ZN(new_n643));
  OAI22_X1  g442(.A1(new_n636), .A2(new_n639), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n433), .B1(new_n442), .B2(new_n414), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n435), .B1(new_n438), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n582), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n554), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n523), .B1(new_n571), .B2(KEYINPUT40), .ZN(new_n649));
  AND3_X1   g448(.A1(new_n563), .A2(KEYINPUT40), .A3(new_n567), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n554), .B1(new_n651), .B2(new_n581), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT85), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n520), .A2(new_n525), .A3(new_n531), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n584), .A2(new_n644), .A3(new_n648), .A4(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT86), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n555), .A2(new_n641), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n658), .A2(new_n581), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT35), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n659), .A2(new_n660), .A3(new_n444), .ZN(new_n661));
  OAI21_X1  g460(.A(KEYINPUT35), .B1(new_n658), .B2(new_n647), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AND3_X1   g462(.A1(new_n656), .A2(new_n657), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n657), .B1(new_n656), .B2(new_n663), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n364), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT95), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI211_X1 g467(.A(KEYINPUT95), .B(new_n364), .C1(new_n664), .C2(new_n665), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n340), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n646), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(G1gat), .ZN(G1324gat));
  INV_X1    g472(.A(KEYINPUT103), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n670), .A2(new_n581), .ZN(new_n675));
  XNOR2_X1  g474(.A(KEYINPUT16), .B(G8gat), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n674), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n677), .A2(KEYINPUT42), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n675), .A2(G8gat), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n677), .A2(KEYINPUT42), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(G1325gat));
  INV_X1    g480(.A(new_n644), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n670), .A2(G15gat), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n656), .A2(new_n663), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT86), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n656), .A2(new_n657), .A3(new_n663), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(KEYINPUT95), .B1(new_n687), .B2(new_n364), .ZN(new_n688));
  INV_X1    g487(.A(new_n669), .ZN(new_n689));
  OAI211_X1 g488(.A(new_n641), .B(new_n339), .C1(new_n688), .C2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT104), .ZN(new_n691));
  AND3_X1   g490(.A1(new_n690), .A2(new_n691), .A3(new_n611), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n691), .B1(new_n690), .B2(new_n611), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n683), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(KEYINPUT105), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n696), .B(new_n683), .C1(new_n692), .C2(new_n693), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(G1326gat));
  XNOR2_X1  g497(.A(KEYINPUT43), .B(G22gat), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  OAI211_X1 g499(.A(new_n554), .B(new_n339), .C1(new_n688), .C2(new_n689), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(KEYINPUT106), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT107), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n670), .A2(new_n704), .A3(new_n554), .ZN(new_n705));
  AND3_X1   g504(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n703), .B1(new_n702), .B2(new_n705), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n700), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n701), .A2(KEYINPUT106), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n704), .B1(new_n670), .B2(new_n554), .ZN(new_n710));
  OAI21_X1  g509(.A(KEYINPUT107), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n711), .A2(new_n699), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n708), .A2(new_n713), .ZN(G1327gat));
  NOR2_X1   g513(.A1(new_n317), .A2(new_n338), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n716), .A2(new_n275), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n718), .B1(new_n668), .B2(new_n669), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n719), .A2(new_n223), .A3(new_n671), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT45), .ZN(new_n721));
  OAI211_X1 g520(.A(KEYINPUT44), .B(new_n274), .C1(new_n664), .C2(new_n665), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n656), .A2(new_n663), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n723), .B1(new_n724), .B2(new_n275), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n716), .A2(new_n363), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(G29gat), .B1(new_n728), .B2(new_n646), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n721), .A2(new_n729), .ZN(G1328gat));
  INV_X1    g529(.A(KEYINPUT46), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n719), .A2(new_n211), .A3(new_n581), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(KEYINPUT108), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n732), .A2(KEYINPUT108), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n731), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n732), .A2(KEYINPUT108), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n737), .A2(KEYINPUT46), .A3(new_n733), .ZN(new_n738));
  OAI21_X1  g537(.A(G36gat), .B1(new_n728), .B2(new_n582), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n736), .A2(new_n738), .A3(new_n739), .ZN(G1329gat));
  AND2_X1   g539(.A1(new_n719), .A2(new_n641), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n741), .A2(new_n220), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n682), .A2(new_n220), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n728), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT47), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT47), .ZN(new_n746));
  OAI221_X1 g545(.A(new_n746), .B1(new_n728), .B2(new_n743), .C1(new_n741), .C2(new_n220), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(G1330gat));
  NAND4_X1  g547(.A1(new_n722), .A2(new_n554), .A3(new_n725), .A4(new_n727), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n749), .A2(G50gat), .ZN(new_n750));
  OR2_X1    g549(.A1(new_n719), .A2(KEYINPUT109), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n554), .A2(new_n204), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n752), .B1(new_n719), .B2(KEYINPUT109), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n750), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g554(.A(new_n338), .ZN(new_n756));
  NOR4_X1   g555(.A1(new_n724), .A2(new_n364), .A3(new_n321), .A4(new_n756), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT110), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n671), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n581), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n762), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n763));
  XOR2_X1   g562(.A(KEYINPUT49), .B(G64gat), .Z(new_n764));
  OAI21_X1  g563(.A(new_n763), .B1(new_n762), .B2(new_n764), .ZN(G1333gat));
  NOR2_X1   g564(.A1(new_n634), .A2(G71gat), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n759), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(G71gat), .B1(new_n758), .B2(new_n644), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT50), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n769), .B(new_n770), .ZN(G1334gat));
  NAND2_X1  g570(.A1(new_n759), .A2(new_n554), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g572(.A1(new_n364), .A2(new_n317), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n338), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n726), .A2(new_n776), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n777), .A2(new_n671), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n724), .A2(new_n275), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n774), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT51), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n782), .A2(KEYINPUT111), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n779), .A2(KEYINPUT51), .A3(new_n774), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n782), .A2(KEYINPUT111), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n671), .A2(new_n235), .A3(new_n338), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT112), .ZN(new_n788));
  OAI22_X1  g587(.A1(new_n778), .A2(new_n235), .B1(new_n786), .B2(new_n788), .ZN(G1336gat));
  NAND2_X1  g588(.A1(new_n777), .A2(new_n581), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(G92gat), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n582), .A2(G92gat), .A3(new_n756), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n785), .A2(new_n783), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n782), .A2(new_n784), .ZN(new_n796));
  AOI22_X1  g595(.A1(new_n790), .A2(G92gat), .B1(new_n796), .B2(new_n794), .ZN(new_n797));
  OAI22_X1  g596(.A1(new_n793), .A2(new_n795), .B1(new_n797), .B2(new_n792), .ZN(G1337gat));
  AND2_X1   g597(.A1(new_n777), .A2(new_n682), .ZN(new_n799));
  INV_X1    g598(.A(G99gat), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n641), .A2(new_n800), .A3(new_n338), .ZN(new_n801));
  OAI22_X1  g600(.A1(new_n799), .A2(new_n800), .B1(new_n786), .B2(new_n801), .ZN(G1338gat));
  NAND3_X1  g601(.A1(new_n726), .A2(new_n554), .A3(new_n776), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n803), .A2(G106gat), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n555), .A2(G106gat), .A3(new_n756), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n796), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT53), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT53), .B1(new_n803), .B2(G106gat), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n783), .A2(new_n785), .A3(new_n805), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT113), .ZN(new_n810));
  AND3_X1   g609(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n810), .B1(new_n808), .B2(new_n809), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n807), .B1(new_n811), .B2(new_n812), .ZN(G1339gat));
  AND3_X1   g612(.A1(new_n326), .A2(KEYINPUT114), .A3(new_n328), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT114), .B1(new_n326), .B2(new_n328), .ZN(new_n815));
  OAI211_X1 g614(.A(KEYINPUT54), .B(new_n329), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n326), .A2(new_n328), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n334), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n816), .A2(KEYINPUT55), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n337), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n816), .A2(new_n819), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n824), .A2(new_n360), .A3(new_n362), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n342), .B1(new_n341), .B2(new_n343), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n348), .A2(new_n349), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n358), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n828), .B1(new_n351), .B2(new_n359), .ZN(new_n829));
  OR2_X1    g628(.A1(new_n829), .A2(new_n756), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n274), .B1(new_n825), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n824), .A2(new_n274), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n832), .A2(new_n829), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n316), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n318), .A2(new_n363), .A3(new_n320), .A4(new_n756), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n646), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n836), .A2(new_n659), .ZN(new_n837));
  AOI21_X1  g636(.A(G113gat), .B1(new_n837), .B2(new_n364), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n554), .B1(new_n834), .B2(new_n835), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n581), .A2(new_n646), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(new_n634), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n363), .A2(new_n392), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n838), .B1(new_n843), .B2(new_n844), .ZN(G1340gat));
  AOI21_X1  g644(.A(new_n390), .B1(new_n843), .B2(new_n338), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n756), .A2(G120gat), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n846), .B1(new_n837), .B2(new_n847), .ZN(new_n848));
  XOR2_X1   g647(.A(new_n848), .B(KEYINPUT115), .Z(G1341gat));
  INV_X1    g648(.A(new_n843), .ZN(new_n850));
  OAI21_X1  g649(.A(G127gat), .B1(new_n850), .B2(new_n316), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n837), .A2(new_n385), .A3(new_n317), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(G1342gat));
  NAND3_X1  g652(.A1(new_n837), .A2(new_n383), .A3(new_n274), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n854), .A2(KEYINPUT56), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(KEYINPUT116), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n383), .B1(new_n843), .B2(new_n274), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n857), .B1(KEYINPUT56), .B2(new_n854), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT117), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n856), .A2(new_n861), .A3(new_n858), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(new_n862), .ZN(G1343gat));
  NAND2_X1  g662(.A1(new_n834), .A2(new_n835), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n555), .A2(KEYINPUT57), .ZN(new_n865));
  AOI211_X1 g664(.A(new_n682), .B(new_n841), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT55), .B1(new_n823), .B2(KEYINPUT118), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n816), .A2(new_n868), .A3(new_n819), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n821), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n870), .A2(new_n360), .A3(new_n362), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n274), .B1(new_n871), .B2(new_n830), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n316), .B1(new_n872), .B2(new_n833), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n555), .B1(new_n873), .B2(new_n835), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT57), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n866), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n364), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT58), .B1(new_n878), .B2(G141gat), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n364), .A2(new_n373), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n836), .A2(new_n554), .A3(new_n644), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n881), .A2(KEYINPUT120), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(KEYINPUT120), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n882), .A2(new_n582), .A3(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n879), .B1(new_n880), .B2(new_n884), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n878), .A2(KEYINPUT119), .A3(G141gat), .ZN(new_n886));
  AOI21_X1  g685(.A(KEYINPUT119), .B1(new_n878), .B2(G141gat), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n881), .A2(new_n581), .A3(new_n880), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT58), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n885), .B1(new_n889), .B2(new_n890), .ZN(G1344gat));
  NAND2_X1  g690(.A1(new_n877), .A2(new_n338), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(new_n893), .A3(G148gat), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT124), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n644), .A2(KEYINPUT121), .A3(new_n840), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT121), .B1(new_n644), .B2(new_n840), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n896), .A2(new_n897), .A3(new_n756), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT122), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n554), .A2(KEYINPUT57), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n900), .B1(new_n834), .B2(new_n835), .ZN(new_n901));
  OAI22_X1  g700(.A1(new_n899), .A2(new_n901), .B1(new_n874), .B2(KEYINPUT57), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n901), .A2(new_n899), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n898), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(G148gat), .B1(new_n904), .B2(KEYINPUT123), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT123), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n901), .A2(new_n899), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n874), .A2(KEYINPUT57), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n901), .A2(new_n899), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n906), .B1(new_n910), .B2(new_n898), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n895), .B(KEYINPUT59), .C1(new_n905), .C2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n910), .A2(new_n906), .A3(new_n898), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n904), .A2(KEYINPUT123), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n914), .A2(new_n915), .A3(G148gat), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n895), .B1(new_n916), .B2(KEYINPUT59), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n894), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(new_n884), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n375), .A3(new_n338), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(G1345gat));
  NAND3_X1  g720(.A1(new_n919), .A2(new_n308), .A3(new_n317), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n877), .A2(new_n317), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n308), .B2(new_n923), .ZN(G1346gat));
  AOI21_X1  g723(.A(G162gat), .B1(new_n919), .B2(new_n274), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n275), .A2(new_n267), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n925), .B1(new_n877), .B2(new_n926), .ZN(G1347gat));
  NOR2_X1   g726(.A1(new_n582), .A2(new_n671), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n929), .A2(new_n634), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n839), .A2(new_n930), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n931), .A2(new_n463), .A3(new_n363), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n671), .B1(new_n834), .B2(new_n835), .ZN(new_n933));
  AND4_X1   g732(.A1(new_n581), .A2(new_n933), .A3(new_n555), .A4(new_n641), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(new_n364), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n932), .B1(new_n935), .B2(new_n463), .ZN(G1348gat));
  NAND3_X1  g735(.A1(new_n934), .A2(new_n464), .A3(new_n338), .ZN(new_n937));
  OAI21_X1  g736(.A(G176gat), .B1(new_n931), .B2(new_n756), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(G1349gat));
  INV_X1    g738(.A(new_n931), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n474), .B1(new_n940), .B2(new_n317), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n316), .A2(new_n491), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n941), .B1(new_n934), .B2(new_n942), .ZN(new_n943));
  XOR2_X1   g742(.A(new_n943), .B(KEYINPUT60), .Z(G1350gat));
  OAI21_X1  g743(.A(G190gat), .B1(new_n931), .B2(new_n275), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT61), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n934), .A2(new_n475), .A3(new_n274), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(G1351gat));
  XNOR2_X1  g747(.A(KEYINPUT125), .B(G197gat), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n682), .A2(new_n929), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n910), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n949), .B1(new_n951), .B2(new_n363), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n933), .A2(new_n581), .A3(new_n554), .A4(new_n644), .ZN(new_n953));
  OR2_X1    g752(.A1(new_n363), .A2(new_n949), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(G1352gat));
  NOR3_X1   g754(.A1(new_n953), .A2(G204gat), .A3(new_n756), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n956), .B(KEYINPUT62), .ZN(new_n957));
  OAI21_X1  g756(.A(G204gat), .B1(new_n951), .B2(new_n756), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1353gat));
  OR3_X1    g758(.A1(new_n953), .A2(G211gat), .A3(new_n316), .ZN(new_n960));
  OAI211_X1 g759(.A(new_n317), .B(new_n950), .C1(new_n902), .C2(new_n903), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n961), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n962));
  AOI21_X1  g761(.A(KEYINPUT63), .B1(new_n961), .B2(G211gat), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n960), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT126), .ZN(G1354gat));
  OAI21_X1  g764(.A(G218gat), .B1(new_n951), .B2(new_n275), .ZN(new_n966));
  OR3_X1    g765(.A1(new_n953), .A2(G218gat), .A3(new_n275), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  XOR2_X1   g767(.A(new_n968), .B(KEYINPUT127), .Z(G1355gat));
endmodule


