//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 1 1 1 1 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 1 0 1 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 1 0 0 0 1 1 0 0 1 1 0 1 0 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n790, new_n791, new_n792,
    new_n794, new_n795, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891;
  INV_X1    g000(.A(G155gat), .ZN(new_n202));
  INV_X1    g001(.A(G162gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT80), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(G155gat), .B2(G162gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT80), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n204), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT81), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n209), .ZN(new_n211));
  XOR2_X1   g010(.A(G141gat), .B(G148gat), .Z(new_n212));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n212), .B1(new_n213), .B2(new_n204), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n210), .A2(new_n211), .A3(new_n214), .ZN(new_n215));
  NOR3_X1   g014(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n204), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT82), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n217), .B1(new_n218), .B2(new_n212), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(new_n218), .B2(new_n212), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G113gat), .B(G120gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  XOR2_X1   g022(.A(G127gat), .B(G134gat), .Z(new_n224));
  XNOR2_X1  g023(.A(new_n223), .B(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  OR3_X1    g025(.A1(new_n221), .A2(KEYINPUT4), .A3(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT4), .B1(new_n221), .B2(new_n226), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n215), .A2(new_n220), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT3), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n221), .A2(KEYINPUT3), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n232), .A2(new_n226), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT5), .ZN(new_n235));
  NAND2_X1  g034(.A1(G225gat), .A2(G233gat), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n229), .A2(new_n234), .A3(new_n235), .A4(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n229), .A2(new_n236), .A3(new_n234), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n221), .B(new_n226), .ZN(new_n239));
  INV_X1    g038(.A(new_n236), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n235), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  AOI22_X1  g040(.A1(KEYINPUT83), .A2(new_n237), .B1(new_n238), .B2(new_n241), .ZN(new_n242));
  AND2_X1   g041(.A1(new_n229), .A2(new_n234), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT83), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n243), .A2(new_n244), .A3(new_n235), .A4(new_n236), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n242), .A2(new_n245), .ZN(new_n246));
  XOR2_X1   g045(.A(G1gat), .B(G29gat), .Z(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(G85gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT0), .B(G57gat), .ZN(new_n249));
  XOR2_X1   g048(.A(new_n248), .B(new_n249), .Z(new_n250));
  NAND2_X1  g049(.A1(new_n246), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT6), .ZN(new_n252));
  INV_X1    g051(.A(new_n250), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n242), .A2(new_n253), .A3(new_n245), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n251), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n246), .A2(KEYINPUT6), .A3(new_n250), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT77), .ZN(new_n259));
  NAND2_X1  g058(.A1(G226gat), .A2(G233gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(G183gat), .A2(G190gat), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n263), .B1(KEYINPUT67), .B2(KEYINPUT24), .ZN(new_n264));
  NAND2_X1  g063(.A1(G183gat), .A2(G190gat), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n262), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n263), .A2(KEYINPUT24), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n264), .B1(new_n268), .B2(new_n265), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT25), .ZN(new_n271));
  NOR2_X1   g070(.A1(G169gat), .A2(G176gat), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n272), .A2(KEYINPUT23), .ZN(new_n273));
  AOI211_X1 g072(.A(new_n271), .B(new_n273), .C1(G169gat), .C2(G176gat), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT23), .ZN(new_n275));
  OR2_X1    g074(.A1(G169gat), .A2(G176gat), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n270), .B(new_n274), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279));
  XOR2_X1   g078(.A(KEYINPUT64), .B(G176gat), .Z(new_n280));
  INV_X1    g079(.A(G169gat), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n280), .A2(KEYINPUT23), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT65), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n279), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n265), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n261), .B1(new_n285), .B2(KEYINPUT24), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n286), .B1(KEYINPUT24), .B2(new_n285), .ZN(new_n287));
  XNOR2_X1  g086(.A(KEYINPUT64), .B(G176gat), .ZN(new_n288));
  NOR3_X1   g087(.A1(new_n288), .A2(new_n275), .A3(G169gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n283), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n287), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n271), .B1(new_n284), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT66), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n282), .B1(new_n283), .B2(new_n273), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n289), .A2(KEYINPUT65), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n294), .A2(new_n295), .A3(new_n279), .A4(new_n287), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT66), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n296), .A2(new_n297), .A3(new_n271), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n278), .B1(new_n293), .B2(new_n298), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n276), .A2(KEYINPUT26), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT26), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n279), .B1(new_n272), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n265), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n303), .B(KEYINPUT72), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT69), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT27), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n307), .B1(new_n308), .B2(G183gat), .ZN(new_n309));
  AOI21_X1  g108(.A(G190gat), .B1(new_n308), .B2(G183gat), .ZN(new_n310));
  INV_X1    g109(.A(G183gat), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n311), .A2(KEYINPUT69), .A3(KEYINPUT27), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n309), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT28), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT70), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT70), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n313), .A2(new_n317), .A3(new_n314), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n311), .A2(KEYINPUT27), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n310), .A2(KEYINPUT28), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n306), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n313), .A2(new_n317), .A3(new_n314), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n317), .B1(new_n313), .B2(new_n314), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n306), .B(new_n321), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n305), .B1(new_n322), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT73), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n321), .B1(new_n323), .B2(new_n324), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT71), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(new_n325), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT73), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n331), .A2(new_n332), .A3(new_n305), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n299), .B1(new_n328), .B2(new_n333), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n259), .B(new_n260), .C1(new_n334), .C2(KEYINPUT29), .ZN(new_n335));
  XNOR2_X1  g134(.A(G197gat), .B(G204gat), .ZN(new_n336));
  AND2_X1   g135(.A1(G211gat), .A2(G218gat), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n336), .B1(KEYINPUT22), .B2(new_n337), .ZN(new_n338));
  NOR2_X1   g137(.A1(G211gat), .A2(G218gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  XOR2_X1   g139(.A(new_n338), .B(new_n340), .Z(new_n341));
  NOR2_X1   g140(.A1(new_n292), .A2(KEYINPUT66), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n297), .B1(new_n296), .B2(new_n271), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n277), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n327), .ZN(new_n345));
  INV_X1    g144(.A(new_n260), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT77), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n332), .B1(new_n331), .B2(new_n305), .ZN(new_n349));
  AOI211_X1 g148(.A(KEYINPUT73), .B(new_n304), .C1(new_n330), .C2(new_n325), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n344), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT29), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n346), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n335), .B(new_n341), .C1(new_n348), .C2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n334), .A2(new_n346), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n345), .A2(new_n352), .A3(new_n260), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n341), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G8gat), .B(G36gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(G92gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(KEYINPUT78), .B(G64gat), .ZN(new_n362));
  XOR2_X1   g161(.A(new_n361), .B(new_n362), .Z(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n354), .A2(new_n359), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT38), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT37), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n354), .A2(new_n368), .A3(new_n359), .ZN(new_n369));
  AND2_X1   g168(.A1(new_n369), .A2(new_n363), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT90), .B1(new_n357), .B2(new_n358), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT90), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n355), .A2(new_n356), .A3(new_n372), .A4(new_n341), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n260), .B1(new_n334), .B2(KEYINPUT29), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n375), .A2(KEYINPUT77), .A3(new_n347), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n341), .B1(new_n376), .B2(new_n335), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT37), .B1(new_n374), .B2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n367), .B1(new_n370), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n369), .A2(new_n363), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n368), .B1(new_n354), .B2(new_n359), .ZN(new_n381));
  NOR3_X1   g180(.A1(new_n380), .A2(new_n366), .A3(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n258), .B1(new_n379), .B2(new_n382), .ZN(new_n383));
  AND3_X1   g182(.A1(new_n354), .A2(new_n359), .A3(new_n364), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT79), .B1(new_n384), .B2(KEYINPUT30), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n364), .B1(new_n354), .B2(new_n359), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n386), .B1(new_n384), .B2(KEYINPUT30), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT79), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT30), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n365), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n385), .A2(new_n387), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT40), .ZN(new_n392));
  AOI211_X1 g191(.A(KEYINPUT39), .B(new_n236), .C1(new_n229), .C2(new_n234), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT88), .B1(new_n393), .B2(new_n250), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT88), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n229), .A2(new_n234), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(new_n240), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n395), .B(new_n253), .C1(new_n397), .C2(KEYINPUT39), .ZN(new_n398));
  AND2_X1   g197(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  OR2_X1    g198(.A1(new_n239), .A2(new_n240), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n400), .A2(KEYINPUT39), .ZN(new_n401));
  AND2_X1   g200(.A1(new_n401), .A2(new_n397), .ZN(new_n402));
  OAI211_X1 g201(.A(KEYINPUT89), .B(new_n392), .C1(new_n399), .C2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT89), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n394), .A2(new_n398), .B1(new_n397), .B2(new_n401), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n404), .B1(new_n405), .B2(KEYINPUT40), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n253), .B1(new_n242), .B2(new_n245), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n407), .B1(new_n405), .B2(KEYINPUT40), .ZN(new_n408));
  AND3_X1   g207(.A1(new_n403), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n391), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n341), .A2(KEYINPUT85), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n338), .A2(new_n340), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n411), .B(new_n352), .C1(KEYINPUT85), .C2(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n230), .B1(new_n413), .B2(new_n231), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n358), .B1(new_n232), .B2(new_n352), .ZN(new_n415));
  INV_X1    g214(.A(G228gat), .ZN(new_n416));
  INV_X1    g215(.A(G233gat), .ZN(new_n417));
  OAI22_X1  g216(.A1(new_n414), .A2(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT86), .ZN(new_n419));
  AND2_X1   g218(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n231), .B1(new_n341), .B2(KEYINPUT29), .ZN(new_n421));
  AOI211_X1 g220(.A(new_n416), .B(new_n417), .C1(new_n421), .C2(new_n221), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n422), .B1(new_n415), .B2(new_n419), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n418), .B1(new_n420), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(G22gat), .ZN(new_n425));
  INV_X1    g224(.A(G22gat), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n418), .B(new_n426), .C1(new_n420), .C2(new_n423), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT87), .B1(new_n424), .B2(G22gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(G50gat), .ZN(new_n431));
  XOR2_X1   g230(.A(G78gat), .B(G106gat), .Z(new_n432));
  XOR2_X1   g231(.A(new_n431), .B(new_n432), .Z(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n428), .B1(new_n429), .B2(new_n434), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n425), .A2(KEYINPUT87), .A3(new_n427), .A4(new_n433), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n383), .A2(new_n410), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT36), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n351), .A2(new_n226), .ZN(new_n440));
  NAND2_X1  g239(.A1(G227gat), .A2(G233gat), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n225), .B(new_n344), .C1(new_n349), .C2(new_n350), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT76), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT34), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n445), .B1(new_n443), .B2(new_n444), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  XOR2_X1   g247(.A(G71gat), .B(G99gat), .Z(new_n449));
  XNOR2_X1  g248(.A(new_n449), .B(KEYINPUT75), .ZN(new_n450));
  XNOR2_X1  g249(.A(G15gat), .B(G43gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n450), .B(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n441), .B1(new_n440), .B2(new_n442), .ZN(new_n453));
  OAI211_X1 g252(.A(KEYINPUT74), .B(new_n452), .C1(new_n453), .C2(KEYINPUT33), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT32), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n452), .A2(KEYINPUT33), .ZN(new_n456));
  NOR3_X1   g255(.A1(new_n453), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT74), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n459), .B(new_n452), .C1(new_n453), .C2(KEYINPUT33), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n440), .A2(new_n442), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT32), .B1(new_n461), .B2(new_n441), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n448), .A2(new_n458), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n448), .B1(new_n463), .B2(new_n458), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n439), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n458), .A2(new_n463), .ZN(new_n468));
  INV_X1    g267(.A(new_n448), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n470), .A2(KEYINPUT36), .A3(new_n464), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n385), .A2(new_n387), .A3(new_n257), .A4(new_n390), .ZN(new_n472));
  INV_X1    g271(.A(new_n437), .ZN(new_n473));
  AOI22_X1  g272(.A1(new_n467), .A2(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n438), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT35), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n470), .A2(KEYINPUT91), .A3(new_n437), .A4(new_n464), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n476), .B1(new_n477), .B2(new_n472), .ZN(new_n478));
  AND4_X1   g277(.A1(KEYINPUT91), .A2(new_n470), .A3(new_n437), .A4(new_n464), .ZN(new_n479));
  INV_X1    g278(.A(new_n472), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n479), .A2(KEYINPUT35), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n475), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(G57gat), .B(G64gat), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT9), .ZN(new_n484));
  NAND2_X1  g283(.A1(G71gat), .A2(G78gat), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n485), .ZN(new_n487));
  NOR2_X1   g286(.A1(G71gat), .A2(G78gat), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n485), .A2(KEYINPUT96), .ZN(new_n490));
  OR3_X1    g289(.A1(new_n486), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n489), .B1(new_n486), .B2(new_n490), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(KEYINPUT97), .B(KEYINPUT21), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n496), .B(G127gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n497), .B(G155gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(G183gat), .B(G211gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n499), .B(KEYINPUT100), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(KEYINPUT19), .ZN(new_n501));
  XOR2_X1   g300(.A(new_n501), .B(KEYINPUT20), .Z(new_n502));
  XNOR2_X1  g301(.A(new_n498), .B(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G15gat), .B(G22gat), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT16), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n504), .B1(new_n505), .B2(G1gat), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n506), .B1(G1gat), .B2(new_n504), .ZN(new_n507));
  INV_X1    g306(.A(G8gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n507), .B(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n493), .B(KEYINPUT99), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n510), .B1(new_n511), .B2(KEYINPUT21), .ZN(new_n512));
  NAND2_X1  g311(.A1(G231gat), .A2(G233gat), .ZN(new_n513));
  XOR2_X1   g312(.A(new_n513), .B(KEYINPUT98), .Z(new_n514));
  XNOR2_X1  g313(.A(new_n512), .B(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n503), .B(new_n515), .ZN(new_n516));
  AND2_X1   g315(.A1(G232gat), .A2(G233gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT41), .ZN(new_n518));
  NOR2_X1   g317(.A1(G29gat), .A2(G36gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(KEYINPUT14), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT92), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n521), .B1(G29gat), .B2(G36gat), .ZN(new_n522));
  INV_X1    g321(.A(G29gat), .ZN(new_n523));
  INV_X1    g322(.A(G36gat), .ZN(new_n524));
  NOR3_X1   g323(.A1(new_n523), .A2(new_n524), .A3(KEYINPUT92), .ZN(new_n525));
  NOR3_X1   g324(.A1(new_n520), .A2(new_n522), .A3(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(G43gat), .B(G50gat), .ZN(new_n527));
  AOI22_X1  g326(.A1(new_n526), .A2(KEYINPUT93), .B1(KEYINPUT15), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n526), .B1(KEYINPUT15), .B2(new_n527), .ZN(new_n529));
  OR2_X1    g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n529), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G85gat), .A2(G92gat), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT102), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(KEYINPUT102), .A2(G85gat), .A3(G92gat), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n537), .A2(KEYINPUT7), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n535), .B1(new_n539), .B2(KEYINPUT103), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n540), .B1(KEYINPUT103), .B2(new_n539), .ZN(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT104), .B(G85gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(KEYINPUT105), .B(G92gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(G99gat), .A2(G106gat), .ZN(new_n544));
  AOI22_X1  g343(.A1(new_n542), .A2(new_n543), .B1(KEYINPUT8), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  XOR2_X1   g345(.A(G99gat), .B(G106gat), .Z(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n546), .A2(new_n547), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT106), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT17), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n533), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n530), .A2(new_n554), .A3(new_n531), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n551), .B1(new_n556), .B2(new_n552), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n518), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n517), .A2(KEYINPUT41), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(G162gat), .ZN(new_n560));
  AND2_X1   g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n560), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n562), .B(new_n518), .C1(new_n555), .C2(new_n557), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G190gat), .B(G218gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT107), .ZN(new_n566));
  XOR2_X1   g365(.A(KEYINPUT101), .B(G134gat), .Z(new_n567));
  XOR2_X1   g366(.A(new_n566), .B(new_n567), .Z(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  OR3_X1    g368(.A1(new_n561), .A2(new_n564), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n569), .B1(new_n561), .B2(new_n564), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n551), .A2(new_n493), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n494), .B1(new_n549), .B2(new_n550), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G230gat), .A2(G233gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(KEYINPUT108), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G120gat), .B(G148gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(G176gat), .B(G204gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT10), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n573), .A2(new_n574), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n511), .A2(new_n551), .A3(KEYINPUT10), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n577), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(KEYINPUT109), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT109), .B1(new_n586), .B2(new_n587), .ZN(new_n590));
  OAI211_X1 g389(.A(new_n578), .B(new_n582), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n578), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n577), .B(KEYINPUT110), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n594), .B1(new_n584), .B2(new_n585), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n581), .B1(new_n592), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  NOR3_X1   g396(.A1(new_n516), .A2(new_n572), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n532), .A2(KEYINPUT17), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n599), .A2(new_n509), .A3(new_n556), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n530), .A2(new_n531), .A3(new_n510), .ZN(new_n601));
  NAND2_X1  g400(.A1(G229gat), .A2(G233gat), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n600), .A2(KEYINPUT18), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n532), .A2(new_n509), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(new_n601), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n602), .B(KEYINPUT13), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n603), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n510), .B1(new_n532), .B2(KEYINPUT17), .ZN(new_n610));
  AOI22_X1  g409(.A1(new_n610), .A2(new_n556), .B1(new_n533), .B2(new_n510), .ZN(new_n611));
  AOI21_X1  g410(.A(KEYINPUT18), .B1(new_n611), .B2(new_n602), .ZN(new_n612));
  XNOR2_X1  g411(.A(G113gat), .B(G141gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(G197gat), .ZN(new_n614));
  XOR2_X1   g413(.A(KEYINPUT11), .B(G169gat), .Z(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT12), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NOR3_X1   g417(.A1(new_n609), .A2(new_n612), .A3(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT94), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT18), .ZN(new_n622));
  AND3_X1   g421(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n621), .B1(new_n620), .B2(new_n622), .ZN(new_n624));
  NOR3_X1   g423(.A1(new_n623), .A2(new_n624), .A3(new_n609), .ZN(new_n625));
  OAI21_X1  g424(.A(KEYINPUT95), .B1(new_n625), .B2(new_n617), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT95), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n624), .A2(new_n609), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n627), .B(new_n618), .C1(new_n628), .C2(new_n623), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n619), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n598), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n482), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(new_n258), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(G1gat), .ZN(G1324gat));
  INV_X1    g435(.A(new_n391), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(KEYINPUT42), .B1(new_n638), .B2(new_n508), .ZN(new_n639));
  NAND2_X1  g438(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n505), .A2(new_n508), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n638), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  MUX2_X1   g441(.A(KEYINPUT42), .B(new_n639), .S(new_n642), .Z(G1325gat));
  NAND2_X1  g442(.A1(new_n467), .A2(new_n471), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  AND3_X1   g444(.A1(new_n634), .A2(G15gat), .A3(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n465), .A2(new_n466), .ZN(new_n647));
  AOI21_X1  g446(.A(G15gat), .B1(new_n634), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n646), .A2(new_n648), .ZN(G1326gat));
  NOR2_X1   g448(.A1(new_n633), .A2(new_n437), .ZN(new_n650));
  XOR2_X1   g449(.A(KEYINPUT43), .B(G22gat), .Z(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(G1327gat));
  INV_X1    g451(.A(new_n572), .ZN(new_n653));
  AOI21_X1  g452(.A(KEYINPUT35), .B1(new_n479), .B2(new_n480), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n477), .A2(new_n472), .A3(new_n476), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n653), .B1(new_n656), .B2(new_n475), .ZN(new_n657));
  INV_X1    g456(.A(new_n516), .ZN(new_n658));
  NOR3_X1   g457(.A1(new_n658), .A2(new_n630), .A3(new_n597), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n657), .A2(new_n523), .A3(new_n258), .A4(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT111), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT45), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n438), .A2(new_n474), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n481), .A2(new_n478), .ZN(new_n665));
  OAI211_X1 g464(.A(KEYINPUT112), .B(new_n572), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n482), .A2(KEYINPUT112), .A3(KEYINPUT44), .A4(new_n572), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n668), .A2(new_n669), .A3(new_n659), .ZN(new_n670));
  OAI21_X1  g469(.A(G29gat), .B1(new_n670), .B2(new_n257), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n661), .A2(new_n662), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n663), .A2(new_n671), .A3(new_n672), .ZN(G1328gat));
  AND2_X1   g472(.A1(new_n657), .A2(new_n659), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n674), .A2(new_n524), .A3(new_n391), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n675), .B(KEYINPUT46), .Z(new_n676));
  OAI21_X1  g475(.A(G36gat), .B1(new_n670), .B2(new_n637), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(G1329gat));
  OAI21_X1  g477(.A(G43gat), .B1(new_n670), .B2(new_n644), .ZN(new_n679));
  INV_X1    g478(.A(G43gat), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n674), .A2(new_n680), .A3(new_n647), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT47), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n679), .A2(KEYINPUT47), .A3(new_n681), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(G1330gat));
  OAI21_X1  g485(.A(G50gat), .B1(new_n670), .B2(new_n437), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n437), .A2(G50gat), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT113), .Z(new_n689));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT48), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n687), .A2(new_n690), .A3(KEYINPUT48), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(G1331gat));
  NAND4_X1  g494(.A1(new_n658), .A2(new_n630), .A3(new_n653), .A4(new_n597), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n696), .B1(new_n656), .B2(new_n475), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n258), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g498(.A(new_n637), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT114), .ZN(new_n702));
  NOR2_X1   g501(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(G1333gat));
  NAND2_X1  g503(.A1(new_n697), .A2(new_n645), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n465), .A2(new_n466), .A3(G71gat), .ZN(new_n706));
  AOI22_X1  g505(.A1(new_n705), .A2(G71gat), .B1(new_n697), .B2(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g507(.A1(new_n697), .A2(new_n473), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g509(.A1(new_n631), .A2(new_n658), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n482), .A2(KEYINPUT51), .A3(new_n572), .A4(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT115), .ZN(new_n713));
  OR2_X1    g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n713), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n657), .A2(new_n711), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT51), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n714), .A2(new_n715), .A3(new_n718), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n719), .A2(new_n258), .A3(new_n542), .A4(new_n597), .ZN(new_n720));
  INV_X1    g519(.A(new_n597), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n631), .A2(new_n658), .A3(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n668), .A2(new_n669), .A3(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n723), .A2(new_n257), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n720), .B1(new_n542), .B2(new_n724), .ZN(G1336gat));
  NOR3_X1   g524(.A1(new_n637), .A2(G92gat), .A3(new_n721), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n717), .A2(KEYINPUT116), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n727), .B1(new_n657), .B2(new_n711), .ZN(new_n728));
  AND4_X1   g527(.A1(new_n482), .A2(new_n572), .A3(new_n711), .A4(new_n727), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n726), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(KEYINPUT117), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n668), .A2(new_n391), .A3(new_n669), .A4(new_n722), .ZN(new_n732));
  INV_X1    g531(.A(new_n543), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT117), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n735), .B(new_n726), .C1(new_n728), .C2(new_n729), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n731), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(KEYINPUT52), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n719), .A2(new_n726), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT52), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n739), .A2(new_n740), .A3(new_n734), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n738), .A2(new_n741), .ZN(G1337gat));
  NOR2_X1   g541(.A1(new_n721), .A2(G99gat), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n719), .A2(new_n647), .A3(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(G99gat), .B1(new_n723), .B2(new_n644), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(G1338gat));
  NOR3_X1   g545(.A1(new_n721), .A2(new_n437), .A3(G106gat), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n719), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n668), .A2(new_n473), .A3(new_n669), .A4(new_n722), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G106gat), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT53), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  OR2_X1    g551(.A1(new_n728), .A2(new_n729), .ZN(new_n753));
  AOI22_X1  g552(.A1(new_n753), .A2(new_n747), .B1(new_n749), .B2(G106gat), .ZN(new_n754));
  OAI22_X1  g553(.A1(new_n748), .A2(new_n752), .B1(new_n754), .B2(new_n751), .ZN(G1339gat));
  NAND2_X1  g554(.A1(new_n598), .A2(new_n630), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n604), .A2(new_n601), .A3(new_n606), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT118), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n611), .A2(new_n602), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n616), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT119), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OAI211_X1 g562(.A(KEYINPUT119), .B(new_n616), .C1(new_n759), .C2(new_n760), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n619), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n572), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT54), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n582), .B1(new_n595), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n589), .A2(new_n590), .ZN(new_n769));
  OAI21_X1  g568(.A(KEYINPUT54), .B1(new_n586), .B2(new_n593), .ZN(new_n770));
  OAI211_X1 g569(.A(KEYINPUT55), .B(new_n768), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT55), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n586), .A2(new_n587), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT109), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n770), .B1(new_n775), .B2(new_n588), .ZN(new_n776));
  INV_X1    g575(.A(new_n768), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n772), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n771), .A2(new_n778), .A3(new_n591), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n766), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n597), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n781), .B1(new_n630), .B2(new_n779), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n780), .B1(new_n782), .B2(new_n653), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n756), .B1(new_n783), .B2(new_n658), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n465), .A2(new_n473), .A3(new_n466), .ZN(new_n785));
  AND3_X1   g584(.A1(new_n784), .A2(new_n258), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n637), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n787), .A2(new_n630), .ZN(new_n788));
  XOR2_X1   g587(.A(new_n788), .B(G113gat), .Z(G1340gat));
  OAI21_X1  g588(.A(G120gat), .B1(new_n787), .B2(new_n721), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n721), .A2(G120gat), .ZN(new_n791));
  XOR2_X1   g590(.A(new_n791), .B(KEYINPUT120), .Z(new_n792));
  OAI21_X1  g591(.A(new_n790), .B1(new_n787), .B2(new_n792), .ZN(G1341gat));
  NOR2_X1   g592(.A1(new_n787), .A2(new_n516), .ZN(new_n794));
  XNOR2_X1  g593(.A(KEYINPUT121), .B(G127gat), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n794), .B(new_n795), .ZN(G1342gat));
  INV_X1    g595(.A(G134gat), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n637), .A2(new_n572), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(KEYINPUT122), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n786), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  XOR2_X1   g599(.A(new_n800), .B(KEYINPUT56), .Z(new_n801));
  OAI21_X1  g600(.A(G134gat), .B1(new_n787), .B2(new_n653), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(G1343gat));
  INV_X1    g602(.A(G141gat), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n645), .A2(new_n257), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n637), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n784), .A2(new_n473), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n784), .A2(KEYINPUT57), .A3(new_n473), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n806), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n804), .B1(new_n811), .B2(new_n631), .ZN(new_n812));
  NOR4_X1   g611(.A1(new_n807), .A2(new_n806), .A3(G141gat), .A4(new_n630), .ZN(new_n813));
  OR3_X1    g612(.A1(new_n812), .A2(KEYINPUT58), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(KEYINPUT58), .B1(new_n812), .B2(new_n813), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(G1344gat));
  NOR2_X1   g615(.A1(new_n807), .A2(new_n806), .ZN(new_n817));
  INV_X1    g616(.A(G148gat), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n817), .A2(new_n818), .A3(new_n597), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT59), .ZN(new_n820));
  INV_X1    g619(.A(new_n806), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT123), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n810), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n784), .A2(KEYINPUT123), .A3(KEYINPUT57), .A4(new_n473), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n516), .B1(new_n783), .B2(KEYINPUT124), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT124), .ZN(new_n827));
  AOI211_X1 g626(.A(new_n827), .B(new_n780), .C1(new_n782), .C2(new_n653), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n756), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT57), .B1(new_n829), .B2(new_n473), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n597), .B(new_n821), .C1(new_n825), .C2(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n820), .B1(new_n831), .B2(G148gat), .ZN(new_n832));
  AOI211_X1 g631(.A(KEYINPUT59), .B(new_n818), .C1(new_n811), .C2(new_n597), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n819), .B1(new_n832), .B2(new_n833), .ZN(G1345gat));
  AOI21_X1  g633(.A(G155gat), .B1(new_n817), .B2(new_n658), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n516), .A2(new_n202), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n835), .B1(new_n811), .B2(new_n836), .ZN(G1346gat));
  AND2_X1   g636(.A1(new_n811), .A2(new_n572), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n799), .A2(new_n805), .A3(new_n203), .ZN(new_n839));
  OAI22_X1  g638(.A1(new_n838), .A2(new_n203), .B1(new_n807), .B2(new_n839), .ZN(G1347gat));
  AND2_X1   g639(.A1(new_n784), .A2(new_n257), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n785), .A2(new_n391), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n843), .A2(new_n630), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n844), .B(new_n281), .ZN(G1348gat));
  AND2_X1   g644(.A1(new_n841), .A2(new_n842), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n597), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n847), .A2(G176gat), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n847), .A2(new_n288), .ZN(new_n849));
  OAI21_X1  g648(.A(KEYINPUT125), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n847), .A2(G176gat), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT125), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n851), .B(new_n852), .C1(new_n288), .C2(new_n847), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n850), .A2(new_n853), .ZN(G1349gat));
  INV_X1    g653(.A(new_n320), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n311), .A2(KEYINPUT27), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n846), .B(new_n658), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n311), .B1(new_n843), .B2(new_n516), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT60), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n859), .B(new_n860), .ZN(G1350gat));
  NOR2_X1   g660(.A1(new_n843), .A2(new_n653), .ZN(new_n862));
  NAND2_X1  g661(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XOR2_X1   g663(.A(KEYINPUT61), .B(G190gat), .Z(new_n865));
  OAI21_X1  g664(.A(new_n864), .B1(new_n862), .B2(new_n865), .ZN(G1351gat));
  OR2_X1    g665(.A1(new_n825), .A2(new_n830), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n645), .A2(new_n258), .A3(new_n637), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(new_n631), .A3(new_n868), .ZN(new_n869));
  XOR2_X1   g668(.A(KEYINPUT127), .B(G197gat), .Z(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n645), .A2(new_n637), .A3(new_n437), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n872), .A2(KEYINPUT126), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(KEYINPUT126), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n841), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  OR3_X1    g674(.A1(new_n875), .A2(new_n630), .A3(new_n870), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n871), .A2(new_n876), .ZN(G1352gat));
  NAND3_X1  g676(.A1(new_n867), .A2(new_n597), .A3(new_n868), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(G204gat), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n875), .A2(G204gat), .A3(new_n721), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n880), .B(KEYINPUT62), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(new_n881), .ZN(G1353gat));
  OR3_X1    g681(.A1(new_n875), .A2(G211gat), .A3(new_n516), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n658), .B(new_n868), .C1(new_n825), .C2(new_n830), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n884), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n885));
  AOI21_X1  g684(.A(KEYINPUT63), .B1(new_n884), .B2(G211gat), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n883), .B1(new_n885), .B2(new_n886), .ZN(G1354gat));
  AND2_X1   g686(.A1(new_n867), .A2(new_n868), .ZN(new_n888));
  INV_X1    g687(.A(G218gat), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n653), .A2(new_n889), .ZN(new_n890));
  OR2_X1    g689(.A1(new_n875), .A2(new_n653), .ZN(new_n891));
  AOI22_X1  g690(.A1(new_n888), .A2(new_n890), .B1(new_n889), .B2(new_n891), .ZN(G1355gat));
endmodule


