

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U553 ( .A1(n647), .A2(n533), .ZN(n636) );
  INV_X1 U554 ( .A(KEYINPUT31), .ZN(n699) );
  XOR2_X1 U555 ( .A(KEYINPUT72), .B(n571), .Z(n520) );
  INV_X1 U556 ( .A(KEYINPUT99), .ZN(n691) );
  XNOR2_X1 U557 ( .A(n691), .B(KEYINPUT30), .ZN(n692) );
  XNOR2_X1 U558 ( .A(n693), .B(n692), .ZN(n694) );
  INV_X1 U559 ( .A(n688), .ZN(n715) );
  OR2_X1 U560 ( .A1(n788), .A2(n787), .ZN(n688) );
  NAND2_X1 U561 ( .A1(n688), .A2(G8), .ZN(n776) );
  AND2_X1 U562 ( .A1(n525), .A2(G2104), .ZN(n892) );
  XOR2_X1 U563 ( .A(KEYINPUT73), .B(n576), .Z(n930) );
  NOR2_X1 U564 ( .A1(G651), .A2(n647), .ZN(n642) );
  XOR2_X1 U565 ( .A(KEYINPUT17), .B(n524), .Z(n893) );
  INV_X1 U566 ( .A(G2105), .ZN(n525) );
  NAND2_X1 U567 ( .A1(G101), .A2(n892), .ZN(n521) );
  XOR2_X1 U568 ( .A(KEYINPUT23), .B(n521), .Z(n523) );
  AND2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n888) );
  NAND2_X1 U570 ( .A1(n888), .A2(G113), .ZN(n522) );
  NAND2_X1 U571 ( .A1(n523), .A2(n522), .ZN(n529) );
  NOR2_X1 U572 ( .A1(G2104), .A2(G2105), .ZN(n524) );
  NAND2_X1 U573 ( .A1(G137), .A2(n893), .ZN(n527) );
  NOR2_X1 U574 ( .A1(G2104), .A2(n525), .ZN(n889) );
  NAND2_X1 U575 ( .A1(G125), .A2(n889), .ZN(n526) );
  NAND2_X1 U576 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U577 ( .A1(n529), .A2(n528), .ZN(G160) );
  INV_X1 U578 ( .A(G96), .ZN(G221) );
  INV_X1 U579 ( .A(G651), .ZN(n533) );
  NOR2_X1 U580 ( .A1(G543), .A2(n533), .ZN(n530) );
  XOR2_X1 U581 ( .A(KEYINPUT1), .B(n530), .Z(n646) );
  NAND2_X1 U582 ( .A1(G64), .A2(n646), .ZN(n532) );
  XOR2_X1 U583 ( .A(G543), .B(KEYINPUT0), .Z(n647) );
  NAND2_X1 U584 ( .A1(G52), .A2(n642), .ZN(n531) );
  NAND2_X1 U585 ( .A1(n532), .A2(n531), .ZN(n538) );
  NOR2_X1 U586 ( .A1(G651), .A2(G543), .ZN(n633) );
  NAND2_X1 U587 ( .A1(G90), .A2(n633), .ZN(n535) );
  NAND2_X1 U588 ( .A1(G77), .A2(n636), .ZN(n534) );
  NAND2_X1 U589 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U590 ( .A(KEYINPUT9), .B(n536), .Z(n537) );
  NOR2_X1 U591 ( .A1(n538), .A2(n537), .ZN(G171) );
  INV_X1 U592 ( .A(G171), .ZN(G301) );
  AND2_X1 U593 ( .A1(G138), .A2(n893), .ZN(n543) );
  NAND2_X1 U594 ( .A1(n889), .A2(G126), .ZN(n542) );
  NAND2_X1 U595 ( .A1(G102), .A2(n892), .ZN(n540) );
  NAND2_X1 U596 ( .A1(G114), .A2(n888), .ZN(n539) );
  AND2_X1 U597 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U598 ( .A1(n542), .A2(n541), .ZN(n681) );
  NOR2_X1 U599 ( .A1(n543), .A2(n681), .ZN(G164) );
  NAND2_X1 U600 ( .A1(n633), .A2(G89), .ZN(n544) );
  XNOR2_X1 U601 ( .A(KEYINPUT4), .B(n544), .ZN(n547) );
  NAND2_X1 U602 ( .A1(n636), .A2(G76), .ZN(n545) );
  XOR2_X1 U603 ( .A(KEYINPUT75), .B(n545), .Z(n546) );
  NAND2_X1 U604 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U605 ( .A(n548), .B(KEYINPUT5), .ZN(n553) );
  NAND2_X1 U606 ( .A1(G63), .A2(n646), .ZN(n550) );
  NAND2_X1 U607 ( .A1(G51), .A2(n642), .ZN(n549) );
  NAND2_X1 U608 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U609 ( .A(KEYINPUT6), .B(n551), .Z(n552) );
  NAND2_X1 U610 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U611 ( .A(n554), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U612 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U613 ( .A1(G94), .A2(G452), .ZN(n555) );
  XOR2_X1 U614 ( .A(KEYINPUT66), .B(n555), .Z(G173) );
  NAND2_X1 U615 ( .A1(G7), .A2(G661), .ZN(n556) );
  XNOR2_X1 U616 ( .A(n556), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U617 ( .A(G223), .B(KEYINPUT69), .ZN(n836) );
  NAND2_X1 U618 ( .A1(n836), .A2(G567), .ZN(n557) );
  XOR2_X1 U619 ( .A(KEYINPUT11), .B(n557), .Z(G234) );
  INV_X1 U620 ( .A(G860), .ZN(n590) );
  NAND2_X1 U621 ( .A1(n633), .A2(G81), .ZN(n558) );
  XNOR2_X1 U622 ( .A(n558), .B(KEYINPUT12), .ZN(n560) );
  NAND2_X1 U623 ( .A1(G68), .A2(n636), .ZN(n559) );
  NAND2_X1 U624 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U625 ( .A(KEYINPUT13), .B(n561), .ZN(n567) );
  NAND2_X1 U626 ( .A1(G56), .A2(n646), .ZN(n562) );
  XOR2_X1 U627 ( .A(KEYINPUT14), .B(n562), .Z(n565) );
  NAND2_X1 U628 ( .A1(n642), .A2(G43), .ZN(n563) );
  XOR2_X1 U629 ( .A(KEYINPUT70), .B(n563), .Z(n564) );
  NOR2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X1 U631 ( .A1(n567), .A2(n566), .ZN(n931) );
  NOR2_X1 U632 ( .A1(n590), .A2(n931), .ZN(n568) );
  XNOR2_X1 U633 ( .A(n568), .B(KEYINPUT71), .ZN(G153) );
  NAND2_X1 U634 ( .A1(G54), .A2(n642), .ZN(n574) );
  NAND2_X1 U635 ( .A1(G92), .A2(n633), .ZN(n570) );
  NAND2_X1 U636 ( .A1(G66), .A2(n646), .ZN(n569) );
  NAND2_X1 U637 ( .A1(n570), .A2(n569), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n636), .A2(G79), .ZN(n571) );
  NOR2_X1 U639 ( .A1(n572), .A2(n520), .ZN(n573) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n575), .B(KEYINPUT15), .ZN(n576) );
  OR2_X1 U642 ( .A1(n930), .A2(G868), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n577), .B(KEYINPUT74), .ZN(n579) );
  NAND2_X1 U644 ( .A1(G868), .A2(G301), .ZN(n578) );
  NAND2_X1 U645 ( .A1(n579), .A2(n578), .ZN(G284) );
  NAND2_X1 U646 ( .A1(G78), .A2(n636), .ZN(n581) );
  NAND2_X1 U647 ( .A1(G65), .A2(n646), .ZN(n580) );
  NAND2_X1 U648 ( .A1(n581), .A2(n580), .ZN(n584) );
  NAND2_X1 U649 ( .A1(G91), .A2(n633), .ZN(n582) );
  XNOR2_X1 U650 ( .A(KEYINPUT67), .B(n582), .ZN(n583) );
  NOR2_X1 U651 ( .A1(n584), .A2(n583), .ZN(n586) );
  NAND2_X1 U652 ( .A1(n642), .A2(G53), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n586), .A2(n585), .ZN(G299) );
  INV_X1 U654 ( .A(G868), .ZN(n659) );
  NOR2_X1 U655 ( .A1(G286), .A2(n659), .ZN(n587) );
  XNOR2_X1 U656 ( .A(n587), .B(KEYINPUT76), .ZN(n589) );
  NOR2_X1 U657 ( .A1(G299), .A2(G868), .ZN(n588) );
  NOR2_X1 U658 ( .A1(n589), .A2(n588), .ZN(G297) );
  NAND2_X1 U659 ( .A1(n590), .A2(G559), .ZN(n591) );
  NAND2_X1 U660 ( .A1(n591), .A2(n930), .ZN(n592) );
  XNOR2_X1 U661 ( .A(n592), .B(KEYINPUT16), .ZN(n593) );
  XOR2_X1 U662 ( .A(KEYINPUT77), .B(n593), .Z(G148) );
  NAND2_X1 U663 ( .A1(n930), .A2(G868), .ZN(n594) );
  NOR2_X1 U664 ( .A1(G559), .A2(n594), .ZN(n595) );
  XNOR2_X1 U665 ( .A(n595), .B(KEYINPUT78), .ZN(n597) );
  NOR2_X1 U666 ( .A1(n931), .A2(G868), .ZN(n596) );
  NOR2_X1 U667 ( .A1(n597), .A2(n596), .ZN(G282) );
  NAND2_X1 U668 ( .A1(G99), .A2(n892), .ZN(n599) );
  NAND2_X1 U669 ( .A1(G111), .A2(n888), .ZN(n598) );
  NAND2_X1 U670 ( .A1(n599), .A2(n598), .ZN(n606) );
  NAND2_X1 U671 ( .A1(n893), .A2(G135), .ZN(n600) );
  XNOR2_X1 U672 ( .A(KEYINPUT79), .B(n600), .ZN(n603) );
  NAND2_X1 U673 ( .A1(n889), .A2(G123), .ZN(n601) );
  XOR2_X1 U674 ( .A(KEYINPUT18), .B(n601), .Z(n602) );
  NOR2_X1 U675 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U676 ( .A(KEYINPUT80), .B(n604), .Z(n605) );
  NOR2_X1 U677 ( .A1(n606), .A2(n605), .ZN(n607) );
  XOR2_X1 U678 ( .A(KEYINPUT81), .B(n607), .Z(n1016) );
  XNOR2_X1 U679 ( .A(n1016), .B(G2096), .ZN(n608) );
  XNOR2_X1 U680 ( .A(n608), .B(KEYINPUT82), .ZN(n609) );
  INV_X1 U681 ( .A(G2100), .ZN(n842) );
  NAND2_X1 U682 ( .A1(n609), .A2(n842), .ZN(G156) );
  NAND2_X1 U683 ( .A1(G67), .A2(n646), .ZN(n611) );
  NAND2_X1 U684 ( .A1(G55), .A2(n642), .ZN(n610) );
  NAND2_X1 U685 ( .A1(n611), .A2(n610), .ZN(n615) );
  NAND2_X1 U686 ( .A1(G93), .A2(n633), .ZN(n613) );
  NAND2_X1 U687 ( .A1(G80), .A2(n636), .ZN(n612) );
  NAND2_X1 U688 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U689 ( .A1(n615), .A2(n614), .ZN(n658) );
  NAND2_X1 U690 ( .A1(G559), .A2(n930), .ZN(n616) );
  XNOR2_X1 U691 ( .A(n616), .B(n931), .ZN(n656) );
  XOR2_X1 U692 ( .A(KEYINPUT83), .B(n656), .Z(n617) );
  NOR2_X1 U693 ( .A1(G860), .A2(n617), .ZN(n618) );
  XNOR2_X1 U694 ( .A(n658), .B(n618), .ZN(G145) );
  NAND2_X1 U695 ( .A1(G88), .A2(n633), .ZN(n620) );
  NAND2_X1 U696 ( .A1(G75), .A2(n636), .ZN(n619) );
  NAND2_X1 U697 ( .A1(n620), .A2(n619), .ZN(n623) );
  NAND2_X1 U698 ( .A1(n646), .A2(G62), .ZN(n621) );
  XOR2_X1 U699 ( .A(KEYINPUT84), .B(n621), .Z(n622) );
  NOR2_X1 U700 ( .A1(n623), .A2(n622), .ZN(n625) );
  NAND2_X1 U701 ( .A1(n642), .A2(G50), .ZN(n624) );
  NAND2_X1 U702 ( .A1(n625), .A2(n624), .ZN(G303) );
  NAND2_X1 U703 ( .A1(G60), .A2(n646), .ZN(n627) );
  NAND2_X1 U704 ( .A1(G47), .A2(n642), .ZN(n626) );
  NAND2_X1 U705 ( .A1(n627), .A2(n626), .ZN(n631) );
  NAND2_X1 U706 ( .A1(G85), .A2(n633), .ZN(n629) );
  NAND2_X1 U707 ( .A1(G72), .A2(n636), .ZN(n628) );
  NAND2_X1 U708 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U709 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U710 ( .A(n632), .B(KEYINPUT65), .ZN(G290) );
  NAND2_X1 U711 ( .A1(G86), .A2(n633), .ZN(n635) );
  NAND2_X1 U712 ( .A1(G61), .A2(n646), .ZN(n634) );
  NAND2_X1 U713 ( .A1(n635), .A2(n634), .ZN(n639) );
  NAND2_X1 U714 ( .A1(n636), .A2(G73), .ZN(n637) );
  XOR2_X1 U715 ( .A(KEYINPUT2), .B(n637), .Z(n638) );
  NOR2_X1 U716 ( .A1(n639), .A2(n638), .ZN(n641) );
  NAND2_X1 U717 ( .A1(n642), .A2(G48), .ZN(n640) );
  NAND2_X1 U718 ( .A1(n641), .A2(n640), .ZN(G305) );
  NAND2_X1 U719 ( .A1(G49), .A2(n642), .ZN(n644) );
  NAND2_X1 U720 ( .A1(G74), .A2(G651), .ZN(n643) );
  NAND2_X1 U721 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U722 ( .A1(n646), .A2(n645), .ZN(n649) );
  NAND2_X1 U723 ( .A1(n647), .A2(G87), .ZN(n648) );
  NAND2_X1 U724 ( .A1(n649), .A2(n648), .ZN(G288) );
  XOR2_X1 U725 ( .A(G303), .B(G290), .Z(n650) );
  XNOR2_X1 U726 ( .A(n650), .B(G305), .ZN(n653) );
  XOR2_X1 U727 ( .A(KEYINPUT19), .B(KEYINPUT85), .Z(n651) );
  XNOR2_X1 U728 ( .A(G288), .B(n651), .ZN(n652) );
  XOR2_X1 U729 ( .A(n653), .B(n652), .Z(n655) );
  XOR2_X1 U730 ( .A(G299), .B(n658), .Z(n654) );
  XNOR2_X1 U731 ( .A(n655), .B(n654), .ZN(n906) );
  XNOR2_X1 U732 ( .A(n656), .B(n906), .ZN(n657) );
  NAND2_X1 U733 ( .A1(n657), .A2(G868), .ZN(n661) );
  NAND2_X1 U734 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U735 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U736 ( .A(KEYINPUT86), .B(n662), .Z(G295) );
  NAND2_X1 U737 ( .A1(G2078), .A2(G2084), .ZN(n663) );
  XNOR2_X1 U738 ( .A(n663), .B(KEYINPUT20), .ZN(n664) );
  XNOR2_X1 U739 ( .A(n664), .B(KEYINPUT87), .ZN(n665) );
  NAND2_X1 U740 ( .A1(n665), .A2(G2090), .ZN(n666) );
  XNOR2_X1 U741 ( .A(KEYINPUT21), .B(n666), .ZN(n667) );
  NAND2_X1 U742 ( .A1(n667), .A2(G2072), .ZN(G158) );
  XOR2_X1 U743 ( .A(KEYINPUT68), .B(G57), .Z(G237) );
  XNOR2_X1 U744 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U745 ( .A1(G108), .A2(G120), .ZN(n668) );
  NOR2_X1 U746 ( .A1(G237), .A2(n668), .ZN(n669) );
  NAND2_X1 U747 ( .A1(G69), .A2(n669), .ZN(n840) );
  NAND2_X1 U748 ( .A1(G567), .A2(n840), .ZN(n670) );
  XOR2_X1 U749 ( .A(KEYINPUT90), .B(n670), .Z(n677) );
  NAND2_X1 U750 ( .A1(G132), .A2(G82), .ZN(n671) );
  XNOR2_X1 U751 ( .A(n671), .B(KEYINPUT22), .ZN(n672) );
  XNOR2_X1 U752 ( .A(n672), .B(KEYINPUT88), .ZN(n673) );
  NOR2_X1 U753 ( .A1(G218), .A2(n673), .ZN(n674) );
  XNOR2_X1 U754 ( .A(n674), .B(KEYINPUT89), .ZN(n675) );
  OR2_X1 U755 ( .A1(G221), .A2(n675), .ZN(n841) );
  AND2_X1 U756 ( .A1(n841), .A2(G2106), .ZN(n676) );
  NOR2_X1 U757 ( .A1(n677), .A2(n676), .ZN(G319) );
  INV_X1 U758 ( .A(G319), .ZN(n679) );
  NAND2_X1 U759 ( .A1(G483), .A2(G661), .ZN(n678) );
  NOR2_X1 U760 ( .A1(n679), .A2(n678), .ZN(n839) );
  NAND2_X1 U761 ( .A1(n839), .A2(G36), .ZN(G176) );
  INV_X1 U762 ( .A(G1384), .ZN(n682) );
  AND2_X1 U763 ( .A1(G138), .A2(n682), .ZN(n680) );
  NAND2_X1 U764 ( .A1(n893), .A2(n680), .ZN(n684) );
  NAND2_X1 U765 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U766 ( .A1(n684), .A2(n683), .ZN(n686) );
  INV_X1 U767 ( .A(KEYINPUT64), .ZN(n685) );
  XNOR2_X1 U768 ( .A(n686), .B(n685), .ZN(n788) );
  NAND2_X1 U769 ( .A1(G160), .A2(G40), .ZN(n787) );
  NOR2_X1 U770 ( .A1(n776), .A2(G1966), .ZN(n687) );
  XNOR2_X1 U771 ( .A(n687), .B(KEYINPUT94), .ZN(n746) );
  INV_X1 U772 ( .A(n715), .ZN(n730) );
  NOR2_X1 U773 ( .A1(G2084), .A2(n730), .ZN(n743) );
  NOR2_X1 U774 ( .A1(n746), .A2(n743), .ZN(n689) );
  XNOR2_X1 U775 ( .A(KEYINPUT98), .B(n689), .ZN(n690) );
  NAND2_X1 U776 ( .A1(n690), .A2(G8), .ZN(n693) );
  NOR2_X1 U777 ( .A1(G168), .A2(n694), .ZN(n698) );
  INV_X1 U778 ( .A(G1961), .ZN(n936) );
  NAND2_X1 U779 ( .A1(n730), .A2(n936), .ZN(n696) );
  XNOR2_X1 U780 ( .A(KEYINPUT25), .B(G2078), .ZN(n957) );
  NAND2_X1 U781 ( .A1(n715), .A2(n957), .ZN(n695) );
  NAND2_X1 U782 ( .A1(n696), .A2(n695), .ZN(n701) );
  NOR2_X1 U783 ( .A1(G171), .A2(n701), .ZN(n697) );
  NOR2_X1 U784 ( .A1(n698), .A2(n697), .ZN(n700) );
  XNOR2_X1 U785 ( .A(n700), .B(n699), .ZN(n745) );
  NAND2_X1 U786 ( .A1(n701), .A2(G171), .ZN(n729) );
  XNOR2_X1 U787 ( .A(KEYINPUT29), .B(KEYINPUT97), .ZN(n727) );
  AND2_X1 U788 ( .A1(n715), .A2(G1996), .ZN(n702) );
  XOR2_X1 U789 ( .A(n702), .B(KEYINPUT26), .Z(n704) );
  NAND2_X1 U790 ( .A1(n730), .A2(G1341), .ZN(n703) );
  NAND2_X1 U791 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U792 ( .A1(n931), .A2(n705), .ZN(n706) );
  OR2_X1 U793 ( .A1(n930), .A2(n706), .ZN(n713) );
  NAND2_X1 U794 ( .A1(n930), .A2(n706), .ZN(n711) );
  NAND2_X1 U795 ( .A1(n730), .A2(G1348), .ZN(n707) );
  XNOR2_X1 U796 ( .A(n707), .B(KEYINPUT96), .ZN(n709) );
  NAND2_X1 U797 ( .A1(n715), .A2(G2067), .ZN(n708) );
  NAND2_X1 U798 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U799 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U800 ( .A1(n713), .A2(n712), .ZN(n720) );
  INV_X1 U801 ( .A(G299), .ZN(n722) );
  NAND2_X1 U802 ( .A1(G1956), .A2(n730), .ZN(n714) );
  XNOR2_X1 U803 ( .A(KEYINPUT95), .B(n714), .ZN(n718) );
  NAND2_X1 U804 ( .A1(n715), .A2(G2072), .ZN(n716) );
  XNOR2_X1 U805 ( .A(KEYINPUT27), .B(n716), .ZN(n717) );
  NOR2_X1 U806 ( .A1(n718), .A2(n717), .ZN(n721) );
  NAND2_X1 U807 ( .A1(n722), .A2(n721), .ZN(n719) );
  NAND2_X1 U808 ( .A1(n720), .A2(n719), .ZN(n725) );
  NOR2_X1 U809 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U810 ( .A(n723), .B(KEYINPUT28), .Z(n724) );
  NAND2_X1 U811 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U812 ( .A(n727), .B(n726), .ZN(n728) );
  NAND2_X1 U813 ( .A1(n729), .A2(n728), .ZN(n744) );
  NOR2_X1 U814 ( .A1(G1971), .A2(n776), .ZN(n732) );
  NOR2_X1 U815 ( .A1(G2090), .A2(n730), .ZN(n731) );
  NOR2_X1 U816 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U817 ( .A(n733), .B(KEYINPUT100), .ZN(n734) );
  NAND2_X1 U818 ( .A1(n734), .A2(G303), .ZN(n736) );
  AND2_X1 U819 ( .A1(n744), .A2(n736), .ZN(n735) );
  NAND2_X1 U820 ( .A1(n745), .A2(n735), .ZN(n740) );
  INV_X1 U821 ( .A(n736), .ZN(n737) );
  OR2_X1 U822 ( .A1(n737), .A2(G286), .ZN(n738) );
  AND2_X1 U823 ( .A1(n738), .A2(G8), .ZN(n739) );
  NAND2_X1 U824 ( .A1(n740), .A2(n739), .ZN(n742) );
  XOR2_X1 U825 ( .A(KEYINPUT101), .B(KEYINPUT32), .Z(n741) );
  XNOR2_X1 U826 ( .A(n742), .B(n741), .ZN(n751) );
  NAND2_X1 U827 ( .A1(G8), .A2(n743), .ZN(n749) );
  AND2_X1 U828 ( .A1(n745), .A2(n744), .ZN(n747) );
  NOR2_X1 U829 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U830 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U831 ( .A1(n751), .A2(n750), .ZN(n775) );
  NOR2_X1 U832 ( .A1(G1976), .A2(G288), .ZN(n756) );
  NOR2_X1 U833 ( .A1(G1971), .A2(G303), .ZN(n752) );
  NOR2_X1 U834 ( .A1(n756), .A2(n752), .ZN(n946) );
  NAND2_X1 U835 ( .A1(n775), .A2(n946), .ZN(n753) );
  XNOR2_X1 U836 ( .A(n753), .B(KEYINPUT102), .ZN(n754) );
  NAND2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n939) );
  NAND2_X1 U838 ( .A1(n754), .A2(n939), .ZN(n755) );
  XNOR2_X1 U839 ( .A(n755), .B(KEYINPUT103), .ZN(n763) );
  INV_X1 U840 ( .A(n776), .ZN(n759) );
  INV_X1 U841 ( .A(KEYINPUT33), .ZN(n765) );
  NAND2_X1 U842 ( .A1(n759), .A2(n756), .ZN(n757) );
  NOR2_X1 U843 ( .A1(n765), .A2(n757), .ZN(n758) );
  XOR2_X1 U844 ( .A(n758), .B(KEYINPUT104), .Z(n764) );
  AND2_X1 U845 ( .A1(n759), .A2(n764), .ZN(n761) );
  XNOR2_X1 U846 ( .A(G1981), .B(G305), .ZN(n928) );
  INV_X1 U847 ( .A(n928), .ZN(n760) );
  AND2_X1 U848 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U849 ( .A1(n763), .A2(n762), .ZN(n769) );
  INV_X1 U850 ( .A(n764), .ZN(n766) );
  OR2_X1 U851 ( .A1(n766), .A2(n765), .ZN(n767) );
  OR2_X1 U852 ( .A1(n928), .A2(n767), .ZN(n768) );
  NAND2_X1 U853 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U854 ( .A(n770), .B(KEYINPUT105), .ZN(n822) );
  NOR2_X1 U855 ( .A1(G1981), .A2(G305), .ZN(n771) );
  XOR2_X1 U856 ( .A(n771), .B(KEYINPUT24), .Z(n772) );
  OR2_X1 U857 ( .A1(n776), .A2(n772), .ZN(n779) );
  NOR2_X1 U858 ( .A1(G2090), .A2(G303), .ZN(n773) );
  NAND2_X1 U859 ( .A1(G8), .A2(n773), .ZN(n774) );
  NAND2_X1 U860 ( .A1(n775), .A2(n774), .ZN(n777) );
  NAND2_X1 U861 ( .A1(n777), .A2(n776), .ZN(n778) );
  AND2_X1 U862 ( .A1(n779), .A2(n778), .ZN(n820) );
  NAND2_X1 U863 ( .A1(G117), .A2(n888), .ZN(n781) );
  NAND2_X1 U864 ( .A1(G141), .A2(n893), .ZN(n780) );
  NAND2_X1 U865 ( .A1(n781), .A2(n780), .ZN(n784) );
  NAND2_X1 U866 ( .A1(n892), .A2(G105), .ZN(n782) );
  XOR2_X1 U867 ( .A(KEYINPUT38), .B(n782), .Z(n783) );
  NOR2_X1 U868 ( .A1(n784), .A2(n783), .ZN(n786) );
  NAND2_X1 U869 ( .A1(n889), .A2(G129), .ZN(n785) );
  NAND2_X1 U870 ( .A1(n786), .A2(n785), .ZN(n873) );
  NOR2_X1 U871 ( .A1(G1996), .A2(n873), .ZN(n1013) );
  INV_X1 U872 ( .A(n788), .ZN(n789) );
  NOR2_X1 U873 ( .A1(n787), .A2(n789), .ZN(n825) );
  NAND2_X1 U874 ( .A1(G1996), .A2(n873), .ZN(n797) );
  INV_X1 U875 ( .A(G1991), .ZN(n851) );
  NAND2_X1 U876 ( .A1(G95), .A2(n892), .ZN(n791) );
  NAND2_X1 U877 ( .A1(G107), .A2(n888), .ZN(n790) );
  NAND2_X1 U878 ( .A1(n791), .A2(n790), .ZN(n795) );
  NAND2_X1 U879 ( .A1(G131), .A2(n893), .ZN(n793) );
  NAND2_X1 U880 ( .A1(G119), .A2(n889), .ZN(n792) );
  NAND2_X1 U881 ( .A1(n793), .A2(n792), .ZN(n794) );
  NOR2_X1 U882 ( .A1(n795), .A2(n794), .ZN(n885) );
  OR2_X1 U883 ( .A1(n851), .A2(n885), .ZN(n796) );
  NAND2_X1 U884 ( .A1(n797), .A2(n796), .ZN(n1008) );
  NAND2_X1 U885 ( .A1(n825), .A2(n1008), .ZN(n824) );
  NOR2_X1 U886 ( .A1(G1986), .A2(G290), .ZN(n798) );
  XOR2_X1 U887 ( .A(n798), .B(KEYINPUT106), .Z(n799) );
  NAND2_X1 U888 ( .A1(n885), .A2(n851), .ZN(n1017) );
  NAND2_X1 U889 ( .A1(n799), .A2(n1017), .ZN(n800) );
  NAND2_X1 U890 ( .A1(n824), .A2(n800), .ZN(n801) );
  XNOR2_X1 U891 ( .A(KEYINPUT107), .B(n801), .ZN(n802) );
  NOR2_X1 U892 ( .A1(n1013), .A2(n802), .ZN(n803) );
  XNOR2_X1 U893 ( .A(KEYINPUT39), .B(n803), .ZN(n815) );
  XOR2_X1 U894 ( .A(G2067), .B(KEYINPUT37), .Z(n816) );
  NAND2_X1 U895 ( .A1(G104), .A2(n892), .ZN(n805) );
  NAND2_X1 U896 ( .A1(G140), .A2(n893), .ZN(n804) );
  NAND2_X1 U897 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U898 ( .A(KEYINPUT34), .B(n806), .ZN(n812) );
  NAND2_X1 U899 ( .A1(n889), .A2(G128), .ZN(n807) );
  XOR2_X1 U900 ( .A(KEYINPUT91), .B(n807), .Z(n809) );
  NAND2_X1 U901 ( .A1(n888), .A2(G116), .ZN(n808) );
  NAND2_X1 U902 ( .A1(n809), .A2(n808), .ZN(n810) );
  XOR2_X1 U903 ( .A(KEYINPUT35), .B(n810), .Z(n811) );
  NOR2_X1 U904 ( .A1(n812), .A2(n811), .ZN(n813) );
  XOR2_X1 U905 ( .A(KEYINPUT36), .B(n813), .Z(n903) );
  NAND2_X1 U906 ( .A1(n816), .A2(n903), .ZN(n814) );
  XOR2_X1 U907 ( .A(KEYINPUT92), .B(n814), .Z(n1020) );
  NAND2_X1 U908 ( .A1(n825), .A2(n1020), .ZN(n830) );
  NAND2_X1 U909 ( .A1(n815), .A2(n830), .ZN(n818) );
  NOR2_X1 U910 ( .A1(n816), .A2(n903), .ZN(n1009) );
  INV_X1 U911 ( .A(n1009), .ZN(n817) );
  NAND2_X1 U912 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U913 ( .A1(n819), .A2(n825), .ZN(n823) );
  AND2_X1 U914 ( .A1(n820), .A2(n823), .ZN(n821) );
  NAND2_X1 U915 ( .A1(n822), .A2(n821), .ZN(n834) );
  INV_X1 U916 ( .A(n823), .ZN(n832) );
  XNOR2_X1 U917 ( .A(KEYINPUT93), .B(n824), .ZN(n828) );
  XOR2_X1 U918 ( .A(G1986), .B(G290), .Z(n945) );
  INV_X1 U919 ( .A(n945), .ZN(n826) );
  AND2_X1 U920 ( .A1(n826), .A2(n825), .ZN(n827) );
  NOR2_X1 U921 ( .A1(n828), .A2(n827), .ZN(n829) );
  AND2_X1 U922 ( .A1(n830), .A2(n829), .ZN(n831) );
  OR2_X1 U923 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U924 ( .A1(n834), .A2(n833), .ZN(n835) );
  XNOR2_X1 U925 ( .A(n835), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U926 ( .A1(G2106), .A2(n836), .ZN(G217) );
  AND2_X1 U927 ( .A1(G15), .A2(G2), .ZN(n837) );
  NAND2_X1 U928 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U929 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U930 ( .A1(n839), .A2(n838), .ZN(G188) );
  XOR2_X1 U931 ( .A(G120), .B(KEYINPUT108), .Z(G236) );
  INV_X1 U933 ( .A(G132), .ZN(G219) );
  INV_X1 U934 ( .A(G108), .ZN(G238) );
  INV_X1 U935 ( .A(G82), .ZN(G220) );
  INV_X1 U936 ( .A(G69), .ZN(G235) );
  NOR2_X1 U937 ( .A1(n841), .A2(n840), .ZN(G325) );
  INV_X1 U938 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U939 ( .A(n842), .B(G2096), .ZN(n844) );
  XNOR2_X1 U940 ( .A(KEYINPUT42), .B(G2678), .ZN(n843) );
  XNOR2_X1 U941 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U942 ( .A(KEYINPUT43), .B(G2090), .Z(n846) );
  XNOR2_X1 U943 ( .A(G2067), .B(G2072), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U945 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U946 ( .A(G2078), .B(G2084), .ZN(n849) );
  XNOR2_X1 U947 ( .A(n850), .B(n849), .ZN(G227) );
  XOR2_X1 U948 ( .A(G1981), .B(G1956), .Z(n853) );
  XOR2_X1 U949 ( .A(n851), .B(G1966), .Z(n852) );
  XNOR2_X1 U950 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U951 ( .A(G1976), .B(G1971), .Z(n855) );
  XOR2_X1 U952 ( .A(G1986), .B(n936), .Z(n854) );
  XNOR2_X1 U953 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U954 ( .A(n857), .B(n856), .Z(n859) );
  XNOR2_X1 U955 ( .A(KEYINPUT109), .B(G2474), .ZN(n858) );
  XNOR2_X1 U956 ( .A(n859), .B(n858), .ZN(n860) );
  XNOR2_X1 U957 ( .A(KEYINPUT41), .B(n860), .ZN(n861) );
  XOR2_X1 U958 ( .A(n861), .B(G1996), .Z(G229) );
  NAND2_X1 U959 ( .A1(n889), .A2(G124), .ZN(n862) );
  XNOR2_X1 U960 ( .A(n862), .B(KEYINPUT44), .ZN(n864) );
  NAND2_X1 U961 ( .A1(G136), .A2(n893), .ZN(n863) );
  NAND2_X1 U962 ( .A1(n864), .A2(n863), .ZN(n865) );
  XNOR2_X1 U963 ( .A(KEYINPUT110), .B(n865), .ZN(n869) );
  NAND2_X1 U964 ( .A1(G100), .A2(n892), .ZN(n867) );
  NAND2_X1 U965 ( .A1(G112), .A2(n888), .ZN(n866) );
  NAND2_X1 U966 ( .A1(n867), .A2(n866), .ZN(n868) );
  NOR2_X1 U967 ( .A1(n869), .A2(n868), .ZN(G162) );
  XOR2_X1 U968 ( .A(KEYINPUT46), .B(KEYINPUT112), .Z(n871) );
  XNOR2_X1 U969 ( .A(G160), .B(KEYINPUT114), .ZN(n870) );
  XNOR2_X1 U970 ( .A(n871), .B(n870), .ZN(n872) );
  XNOR2_X1 U971 ( .A(KEYINPUT48), .B(n872), .ZN(n875) );
  XNOR2_X1 U972 ( .A(n873), .B(KEYINPUT111), .ZN(n874) );
  XNOR2_X1 U973 ( .A(n875), .B(n874), .ZN(n884) );
  NAND2_X1 U974 ( .A1(G103), .A2(n892), .ZN(n877) );
  NAND2_X1 U975 ( .A1(G139), .A2(n893), .ZN(n876) );
  NAND2_X1 U976 ( .A1(n877), .A2(n876), .ZN(n882) );
  NAND2_X1 U977 ( .A1(G115), .A2(n888), .ZN(n879) );
  NAND2_X1 U978 ( .A1(G127), .A2(n889), .ZN(n878) );
  NAND2_X1 U979 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U980 ( .A(KEYINPUT47), .B(n880), .Z(n881) );
  NOR2_X1 U981 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U982 ( .A(KEYINPUT113), .B(n883), .Z(n1004) );
  XOR2_X1 U983 ( .A(n884), .B(n1004), .Z(n887) );
  XNOR2_X1 U984 ( .A(G164), .B(n885), .ZN(n886) );
  XNOR2_X1 U985 ( .A(n887), .B(n886), .ZN(n900) );
  NAND2_X1 U986 ( .A1(G118), .A2(n888), .ZN(n891) );
  NAND2_X1 U987 ( .A1(G130), .A2(n889), .ZN(n890) );
  NAND2_X1 U988 ( .A1(n891), .A2(n890), .ZN(n898) );
  NAND2_X1 U989 ( .A1(G106), .A2(n892), .ZN(n895) );
  NAND2_X1 U990 ( .A1(G142), .A2(n893), .ZN(n894) );
  NAND2_X1 U991 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U992 ( .A(KEYINPUT45), .B(n896), .Z(n897) );
  NOR2_X1 U993 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U994 ( .A(n900), .B(n899), .Z(n902) );
  XNOR2_X1 U995 ( .A(n1016), .B(G162), .ZN(n901) );
  XNOR2_X1 U996 ( .A(n902), .B(n901), .ZN(n904) );
  XNOR2_X1 U997 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U998 ( .A1(G37), .A2(n905), .ZN(G395) );
  XNOR2_X1 U999 ( .A(G286), .B(n906), .ZN(n908) );
  XOR2_X1 U1000 ( .A(n931), .B(G301), .Z(n907) );
  XNOR2_X1 U1001 ( .A(n908), .B(n907), .ZN(n909) );
  XNOR2_X1 U1002 ( .A(n909), .B(n930), .ZN(n910) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n910), .ZN(G397) );
  XOR2_X1 U1004 ( .A(G2451), .B(G2430), .Z(n912) );
  XNOR2_X1 U1005 ( .A(G2438), .B(G2443), .ZN(n911) );
  XNOR2_X1 U1006 ( .A(n912), .B(n911), .ZN(n918) );
  XOR2_X1 U1007 ( .A(G2435), .B(G2454), .Z(n914) );
  XNOR2_X1 U1008 ( .A(G1341), .B(G1348), .ZN(n913) );
  XNOR2_X1 U1009 ( .A(n914), .B(n913), .ZN(n916) );
  XOR2_X1 U1010 ( .A(G2446), .B(G2427), .Z(n915) );
  XNOR2_X1 U1011 ( .A(n916), .B(n915), .ZN(n917) );
  XOR2_X1 U1012 ( .A(n918), .B(n917), .Z(n919) );
  NAND2_X1 U1013 ( .A1(G14), .A2(n919), .ZN(n925) );
  NAND2_X1 U1014 ( .A1(G319), .A2(n925), .ZN(n922) );
  NOR2_X1 U1015 ( .A1(G227), .A2(G229), .ZN(n920) );
  XNOR2_X1 U1016 ( .A(KEYINPUT49), .B(n920), .ZN(n921) );
  NOR2_X1 U1017 ( .A1(n922), .A2(n921), .ZN(n924) );
  NOR2_X1 U1018 ( .A1(G395), .A2(G397), .ZN(n923) );
  NAND2_X1 U1019 ( .A1(n924), .A2(n923), .ZN(G225) );
  INV_X1 U1020 ( .A(G225), .ZN(G308) );
  INV_X1 U1021 ( .A(n925), .ZN(G401) );
  XNOR2_X1 U1022 ( .A(G16), .B(KEYINPUT56), .ZN(n926) );
  XNOR2_X1 U1023 ( .A(n926), .B(KEYINPUT119), .ZN(n950) );
  XOR2_X1 U1024 ( .A(G168), .B(G1966), .Z(n927) );
  NOR2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1026 ( .A(KEYINPUT57), .B(n929), .Z(n944) );
  XNOR2_X1 U1027 ( .A(n930), .B(G1348), .ZN(n933) );
  XOR2_X1 U1028 ( .A(G1341), .B(n931), .Z(n932) );
  NAND2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n942) );
  XOR2_X1 U1030 ( .A(G299), .B(G1956), .Z(n935) );
  NAND2_X1 U1031 ( .A1(G1971), .A2(G303), .ZN(n934) );
  NAND2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n938) );
  XOR2_X1 U1033 ( .A(n936), .B(G301), .Z(n937) );
  NOR2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n940) );
  NAND2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n941) );
  NOR2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1037 ( .A1(n944), .A2(n943), .ZN(n948) );
  NAND2_X1 U1038 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1039 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1040 ( .A1(n950), .A2(n949), .ZN(n1002) );
  INV_X1 U1041 ( .A(KEYINPUT55), .ZN(n1027) );
  XOR2_X1 U1042 ( .A(G25), .B(G1991), .Z(n951) );
  NAND2_X1 U1043 ( .A1(n951), .A2(G28), .ZN(n956) );
  XNOR2_X1 U1044 ( .A(G2067), .B(G26), .ZN(n953) );
  XNOR2_X1 U1045 ( .A(G2072), .B(G33), .ZN(n952) );
  NOR2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(n954), .B(KEYINPUT117), .ZN(n955) );
  NOR2_X1 U1048 ( .A1(n956), .A2(n955), .ZN(n961) );
  XOR2_X1 U1049 ( .A(n957), .B(G27), .Z(n959) );
  XNOR2_X1 U1050 ( .A(G1996), .B(G32), .ZN(n958) );
  NOR2_X1 U1051 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1052 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1053 ( .A(n962), .B(KEYINPUT53), .ZN(n965) );
  XOR2_X1 U1054 ( .A(G2084), .B(G34), .Z(n963) );
  XNOR2_X1 U1055 ( .A(KEYINPUT54), .B(n963), .ZN(n964) );
  NAND2_X1 U1056 ( .A1(n965), .A2(n964), .ZN(n968) );
  XNOR2_X1 U1057 ( .A(KEYINPUT116), .B(G2090), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(G35), .B(n966), .ZN(n967) );
  NOR2_X1 U1059 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1060 ( .A(n1027), .B(n969), .Z(n971) );
  INV_X1 U1061 ( .A(G29), .ZN(n970) );
  NAND2_X1 U1062 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1063 ( .A1(n972), .A2(G11), .ZN(n973) );
  XOR2_X1 U1064 ( .A(KEYINPUT118), .B(n973), .Z(n1000) );
  XOR2_X1 U1065 ( .A(G16), .B(KEYINPUT120), .Z(n998) );
  XOR2_X1 U1066 ( .A(G5), .B(G1961), .Z(n993) );
  XOR2_X1 U1067 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n980) );
  XNOR2_X1 U1068 ( .A(G1971), .B(G22), .ZN(n975) );
  XNOR2_X1 U1069 ( .A(G23), .B(G1976), .ZN(n974) );
  NOR2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n978) );
  XOR2_X1 U1071 ( .A(G1986), .B(KEYINPUT122), .Z(n976) );
  XNOR2_X1 U1072 ( .A(G24), .B(n976), .ZN(n977) );
  NAND2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1074 ( .A(n980), .B(n979), .ZN(n991) );
  XNOR2_X1 U1075 ( .A(KEYINPUT59), .B(G4), .ZN(n981) );
  XNOR2_X1 U1076 ( .A(n981), .B(KEYINPUT121), .ZN(n982) );
  XNOR2_X1 U1077 ( .A(G1348), .B(n982), .ZN(n984) );
  XNOR2_X1 U1078 ( .A(G1981), .B(G6), .ZN(n983) );
  NOR2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n988) );
  XNOR2_X1 U1080 ( .A(G1341), .B(G19), .ZN(n986) );
  XNOR2_X1 U1081 ( .A(G1956), .B(G20), .ZN(n985) );
  NOR2_X1 U1082 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1083 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1084 ( .A(KEYINPUT60), .B(n989), .ZN(n990) );
  NOR2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n995) );
  XNOR2_X1 U1087 ( .A(G21), .B(G1966), .ZN(n994) );
  NOR2_X1 U1088 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1089 ( .A(n996), .B(KEYINPUT61), .ZN(n997) );
  NAND2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1093 ( .A(KEYINPUT124), .B(n1003), .ZN(n1031) );
  XOR2_X1 U1094 ( .A(G2072), .B(n1004), .Z(n1006) );
  XOR2_X1 U1095 ( .A(G164), .B(G2078), .Z(n1005) );
  NOR2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(KEYINPUT50), .B(n1007), .ZN(n1011) );
  NOR2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1025) );
  XOR2_X1 U1100 ( .A(G2090), .B(G162), .Z(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1102 ( .A(KEYINPUT51), .B(n1014), .Z(n1023) );
  XOR2_X1 U1103 ( .A(G2084), .B(G160), .Z(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1018) );
  NAND2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1107 ( .A(KEYINPUT115), .B(n1021), .Z(n1022) );
  NAND2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1109 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1110 ( .A(KEYINPUT52), .B(n1026), .ZN(n1028) );
  NAND2_X1 U1111 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1112 ( .A1(n1029), .A2(G29), .ZN(n1030) );
  NAND2_X1 U1113 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1114 ( .A(n1032), .B(KEYINPUT62), .ZN(n1033) );
  XNOR2_X1 U1115 ( .A(KEYINPUT125), .B(n1033), .ZN(G311) );
  XOR2_X1 U1116 ( .A(KEYINPUT126), .B(G311), .Z(G150) );
  INV_X1 U1117 ( .A(G303), .ZN(G166) );
endmodule

