//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 0 1 1 0 0 0 1 0 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 0 0 1 1 0 0 1 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008;
  INV_X1    g000(.A(KEYINPUT94), .ZN(new_n187));
  INV_X1    g001(.A(G469), .ZN(new_n188));
  XOR2_X1   g002(.A(KEYINPUT77), .B(G902), .Z(new_n189));
  XNOR2_X1  g003(.A(G110), .B(G140), .ZN(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  AND2_X1   g005(.A1(new_n191), .A2(G227), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n190), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G134), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT67), .B1(new_n195), .B2(G137), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT11), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT11), .ZN(new_n198));
  OAI211_X1 g012(.A(KEYINPUT67), .B(new_n198), .C1(new_n195), .C2(G137), .ZN(new_n199));
  INV_X1    g013(.A(G137), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n200), .A2(G134), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n197), .A2(new_n199), .A3(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G131), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n201), .B1(new_n196), .B2(KEYINPUT11), .ZN(new_n205));
  INV_X1    g019(.A(G131), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(new_n199), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n204), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G104), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT3), .B1(new_n209), .B2(G107), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT3), .ZN(new_n211));
  INV_X1    g025(.A(G107), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n212), .A3(G104), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n209), .A2(G107), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n210), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT80), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n210), .A2(new_n213), .A3(KEYINPUT80), .A4(new_n214), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(G101), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G101), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n210), .A2(new_n213), .A3(new_n220), .A4(new_n214), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n221), .A2(KEYINPUT4), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT4), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n217), .A2(new_n224), .A3(G101), .A4(new_n218), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT71), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT0), .B(G128), .ZN(new_n227));
  INV_X1    g041(.A(G143), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT65), .B1(new_n228), .B2(G146), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT65), .ZN(new_n230));
  INV_X1    g044(.A(G146), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n230), .A2(new_n231), .A3(G143), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n234), .B1(new_n231), .B2(G143), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n228), .A2(KEYINPUT66), .A3(G146), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n227), .B1(new_n233), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n231), .A2(G143), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n228), .A2(G146), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n239), .A2(new_n240), .A3(KEYINPUT0), .A4(G128), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n226), .B1(new_n238), .B2(new_n242), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n229), .A2(new_n232), .B1(new_n235), .B2(new_n236), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n241), .B(KEYINPUT71), .C1(new_n244), .C2(new_n227), .ZN(new_n245));
  AND4_X1   g059(.A1(new_n223), .A2(new_n225), .A3(new_n243), .A4(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT81), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n209), .A2(G107), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n212), .A2(G104), .ZN(new_n249));
  OAI21_X1  g063(.A(G101), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n247), .B1(new_n221), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G128), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n253), .A2(KEYINPUT1), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(new_n239), .A3(new_n240), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n253), .B1(new_n239), .B2(KEYINPUT1), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n255), .B1(new_n244), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n221), .A2(new_n250), .A3(new_n247), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n252), .A2(new_n257), .A3(KEYINPUT10), .A4(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n239), .A2(KEYINPUT1), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n260), .A2(G128), .B1(new_n239), .B2(new_n240), .ZN(new_n261));
  INV_X1    g075(.A(new_n255), .ZN(new_n262));
  OAI211_X1 g076(.A(new_n221), .B(new_n250), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT10), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n259), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n208), .B1(new_n246), .B2(new_n266), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n223), .A2(new_n225), .A3(new_n243), .A4(new_n245), .ZN(new_n268));
  INV_X1    g082(.A(new_n207), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n206), .B1(new_n205), .B2(new_n199), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n268), .A2(new_n271), .A3(new_n259), .A4(new_n265), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n194), .B1(new_n267), .B2(new_n272), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n221), .A2(new_n250), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n263), .B1(new_n257), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(KEYINPUT82), .B1(new_n204), .B2(new_n207), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT12), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT12), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n275), .A2(new_n279), .A3(new_n276), .ZN(new_n280));
  AND4_X1   g094(.A1(new_n272), .A2(new_n194), .A3(new_n278), .A4(new_n280), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n188), .B(new_n189), .C1(new_n273), .C2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(G469), .A2(G902), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n272), .A2(new_n278), .A3(new_n280), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n193), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n267), .A2(new_n272), .A3(new_n194), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(G469), .A3(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n282), .A2(new_n283), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT83), .ZN(new_n289));
  XNOR2_X1  g103(.A(KEYINPUT9), .B(G234), .ZN(new_n290));
  OAI21_X1  g104(.A(G221), .B1(new_n290), .B2(G902), .ZN(new_n291));
  AND3_X1   g105(.A1(new_n288), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n289), .B1(new_n288), .B2(new_n291), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G217), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n290), .A2(new_n295), .A3(G953), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT93), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT68), .ZN(new_n298));
  INV_X1    g112(.A(G116), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(KEYINPUT68), .A2(G116), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(G122), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT14), .ZN(new_n303));
  OAI21_X1  g117(.A(G107), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AND2_X1   g118(.A1(KEYINPUT68), .A2(G116), .ZN(new_n305));
  NOR2_X1   g119(.A1(KEYINPUT68), .A2(G116), .ZN(new_n306));
  INV_X1    g120(.A(G122), .ZN(new_n307));
  NOR3_X1   g121(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n299), .A2(G122), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n304), .B1(new_n303), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n228), .A2(G128), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n253), .A2(G143), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G134), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n312), .A2(new_n313), .A3(new_n195), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n309), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n302), .A2(new_n212), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n297), .B1(new_n311), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n212), .B1(new_n308), .B2(KEYINPUT14), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n302), .A2(new_n318), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n322), .B1(KEYINPUT14), .B2(new_n323), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n324), .A2(KEYINPUT93), .A3(new_n319), .A4(new_n317), .ZN(new_n325));
  INV_X1    g139(.A(new_n316), .ZN(new_n326));
  OAI21_X1  g140(.A(G107), .B1(new_n308), .B2(new_n309), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n326), .B1(new_n327), .B2(new_n319), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT90), .B(KEYINPUT13), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n313), .B1(new_n329), .B2(new_n312), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n312), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT91), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT91), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n329), .A2(new_n333), .A3(new_n312), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n330), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n328), .B1(new_n335), .B2(new_n195), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT92), .ZN(new_n337));
  AOI22_X1  g151(.A1(new_n321), .A2(new_n325), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n328), .B(KEYINPUT92), .C1(new_n335), .C2(new_n195), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n296), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n321), .A2(new_n325), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n336), .A2(new_n337), .ZN(new_n342));
  AND4_X1   g156(.A1(new_n339), .A2(new_n341), .A3(new_n342), .A4(new_n296), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n189), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(G478), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n345), .A2(KEYINPUT15), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n341), .A2(new_n342), .A3(new_n339), .ZN(new_n348));
  INV_X1    g162(.A(new_n296), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n338), .A2(new_n339), .A3(new_n296), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n346), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n352), .A2(new_n189), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n347), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G952), .ZN(new_n356));
  AOI211_X1 g170(.A(G953), .B(new_n356), .C1(G234), .C2(G237), .ZN(new_n357));
  AOI211_X1 g171(.A(new_n191), .B(new_n189), .C1(G234), .C2(G237), .ZN(new_n358));
  XNOR2_X1  g172(.A(KEYINPUT21), .B(G898), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G902), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT16), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT78), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n364), .A2(G125), .ZN(new_n365));
  INV_X1    g179(.A(G125), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n366), .A2(KEYINPUT78), .ZN(new_n367));
  OAI21_X1  g181(.A(G140), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(G125), .A2(G140), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n363), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G140), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n363), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n366), .A2(KEYINPUT78), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n364), .A2(G125), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n231), .B1(new_n371), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n372), .B1(new_n374), .B2(new_n375), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT16), .B1(new_n378), .B2(new_n369), .ZN(new_n379));
  INV_X1    g193(.A(new_n376), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(G146), .A3(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(G237), .A2(G953), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(G143), .A3(G214), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(G143), .B1(new_n382), .B2(G214), .ZN(new_n385));
  OAI21_X1  g199(.A(G131), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n385), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(new_n206), .A3(new_n383), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT17), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n386), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n387), .A2(new_n383), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(KEYINPUT17), .A3(G131), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n377), .A2(new_n381), .A3(new_n390), .A4(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(G113), .B(G122), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n394), .B(new_n209), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT89), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n391), .A2(new_n396), .A3(KEYINPUT18), .A4(G131), .ZN(new_n397));
  XNOR2_X1  g211(.A(G125), .B(G140), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(new_n231), .ZN(new_n399));
  XNOR2_X1  g213(.A(KEYINPUT78), .B(G125), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n370), .B1(new_n400), .B2(new_n372), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n399), .B1(new_n401), .B2(new_n231), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n396), .A2(KEYINPUT18), .A3(G131), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n387), .A2(new_n383), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n397), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n393), .A2(new_n395), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n395), .B1(new_n393), .B2(new_n405), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n362), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G475), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n386), .A2(new_n388), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n398), .A2(KEYINPUT19), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n412), .B1(new_n401), .B2(KEYINPUT19), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n381), .B(new_n411), .C1(G146), .C2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n405), .ZN(new_n415));
  INV_X1    g229(.A(new_n395), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n406), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT20), .ZN(new_n419));
  NOR2_X1   g233(.A1(G475), .A2(G902), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n419), .B1(new_n418), .B2(new_n420), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n361), .B(new_n410), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n355), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(G214), .B1(G237), .B2(G902), .ZN(new_n426));
  XOR2_X1   g240(.A(new_n426), .B(KEYINPUT84), .Z(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n300), .A2(G119), .A3(new_n301), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n299), .A2(G119), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n429), .A2(KEYINPUT5), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(G113), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT5), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n433), .B1(new_n430), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT86), .ZN(new_n437));
  XOR2_X1   g251(.A(KEYINPUT2), .B(G113), .Z(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(new_n429), .A3(new_n431), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n274), .A2(new_n436), .A3(new_n437), .A4(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n274), .A2(new_n436), .A3(new_n439), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT86), .ZN(new_n442));
  INV_X1    g256(.A(new_n439), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT69), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n429), .A2(new_n444), .A3(new_n431), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n444), .B1(new_n429), .B2(new_n431), .ZN(new_n446));
  OAI21_X1  g260(.A(KEYINPUT5), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n443), .B1(new_n447), .B2(new_n435), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n440), .B(new_n442), .C1(new_n448), .C2(new_n274), .ZN(new_n449));
  XNOR2_X1  g263(.A(G110), .B(G122), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n450), .B(KEYINPUT85), .ZN(new_n451));
  XOR2_X1   g265(.A(new_n451), .B(KEYINPUT8), .Z(new_n452));
  NAND2_X1  g266(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(KEYINPUT87), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT87), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n448), .A2(new_n274), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n442), .A2(new_n440), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n455), .B(new_n452), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n257), .A2(new_n400), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n374), .A2(new_n375), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n241), .B(new_n461), .C1(new_n244), .C2(new_n227), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n191), .A2(G224), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(KEYINPUT7), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(KEYINPUT7), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n460), .A2(new_n462), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(G119), .ZN(new_n469));
  NOR3_X1   g283(.A1(new_n305), .A2(new_n306), .A3(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(KEYINPUT69), .B1(new_n470), .B2(new_n430), .ZN(new_n471));
  INV_X1    g285(.A(new_n438), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n429), .A2(new_n444), .A3(new_n431), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(KEYINPUT70), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT70), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n471), .A2(new_n476), .A3(new_n472), .A4(new_n473), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n475), .A2(new_n477), .A3(new_n439), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n223), .A2(new_n225), .ZN(new_n479));
  INV_X1    g293(.A(new_n258), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n480), .A2(new_n251), .ZN(new_n481));
  AOI22_X1  g295(.A1(new_n478), .A2(new_n479), .B1(new_n481), .B2(new_n448), .ZN(new_n482));
  INV_X1    g296(.A(new_n451), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n468), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(G902), .B1(new_n459), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(G210), .B1(G237), .B2(G902), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(KEYINPUT88), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n223), .A2(new_n225), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n443), .B1(new_n474), .B2(KEYINPUT70), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n489), .B1(new_n477), .B2(new_n490), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n448), .A2(new_n481), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n451), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n448), .A2(new_n481), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n475), .A2(new_n477), .A3(new_n439), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n483), .B(new_n494), .C1(new_n495), .C2(new_n489), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n493), .A2(KEYINPUT6), .A3(new_n496), .ZN(new_n497));
  OR3_X1    g311(.A1(new_n482), .A2(KEYINPUT6), .A3(new_n483), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n463), .B(new_n464), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n485), .A2(new_n488), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n488), .B1(new_n485), .B2(new_n500), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n425), .B(new_n428), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n187), .B1(new_n294), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n189), .ZN(new_n505));
  INV_X1    g319(.A(new_n272), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n233), .A2(new_n237), .ZN(new_n507));
  INV_X1    g321(.A(new_n256), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n264), .B1(new_n509), .B2(new_n255), .ZN(new_n510));
  AOI22_X1  g324(.A1(new_n481), .A2(new_n510), .B1(new_n264), .B2(new_n263), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n271), .B1(new_n511), .B2(new_n268), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n193), .B1(new_n506), .B2(new_n512), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n272), .A2(new_n194), .A3(new_n278), .A4(new_n280), .ZN(new_n514));
  AOI211_X1 g328(.A(G469), .B(new_n505), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n287), .A2(new_n283), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n291), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT83), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n288), .A2(new_n289), .A3(new_n291), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AND3_X1   g334(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n521));
  INV_X1    g335(.A(new_n458), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n455), .B1(new_n449), .B2(new_n452), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n484), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n362), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n487), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n485), .A2(new_n488), .A3(new_n500), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n427), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n520), .A2(KEYINPUT94), .A3(new_n528), .A4(new_n425), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n530), .B(KEYINPUT22), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n531), .B(G137), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT79), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n253), .A2(G119), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT23), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n469), .A2(G128), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n253), .A2(KEYINPUT23), .A3(G119), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(G110), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n535), .A2(new_n538), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT24), .B(G110), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n544), .B1(new_n377), .B2(new_n381), .ZN(new_n545));
  INV_X1    g359(.A(G110), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n537), .A2(new_n539), .A3(new_n546), .A4(new_n538), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n542), .A2(new_n543), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n381), .A2(new_n399), .A3(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n534), .B1(new_n545), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n542), .A2(new_n543), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n552), .B1(G110), .B2(new_n540), .ZN(new_n553));
  AOI211_X1 g367(.A(new_n231), .B(new_n376), .C1(new_n401), .C2(KEYINPUT16), .ZN(new_n554));
  AOI21_X1  g368(.A(G146), .B1(new_n379), .B2(new_n380), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n549), .A2(new_n399), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n381), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n556), .A2(KEYINPUT79), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n533), .B1(new_n551), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n377), .A2(new_n381), .ZN(new_n562));
  AOI22_X1  g376(.A1(new_n562), .A2(new_n553), .B1(new_n381), .B2(new_n557), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n532), .B1(new_n563), .B2(KEYINPUT79), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n561), .A2(new_n189), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT25), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n295), .B1(new_n189), .B2(G234), .ZN(new_n568));
  NOR3_X1   g382(.A1(new_n560), .A2(new_n564), .A3(new_n505), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT25), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n567), .A2(new_n568), .A3(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n560), .A2(new_n564), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n568), .A2(G902), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n208), .A2(new_n243), .A3(new_n245), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n195), .A2(G137), .ZN(new_n579));
  OAI21_X1  g393(.A(G131), .B1(new_n579), .B2(new_n201), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n257), .A2(new_n207), .A3(new_n580), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(KEYINPUT28), .B1(new_n582), .B2(new_n495), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n382), .A2(G210), .ZN(new_n584));
  XOR2_X1   g398(.A(new_n584), .B(KEYINPUT27), .Z(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(KEYINPUT26), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(G101), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n241), .B1(new_n244), .B2(new_n227), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n581), .B1(new_n271), .B2(new_n588), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n589), .A2(new_n478), .A3(KEYINPUT75), .ZN(new_n590));
  AOI21_X1  g404(.A(KEYINPUT75), .B1(new_n589), .B2(new_n478), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n495), .A2(KEYINPUT72), .A3(new_n578), .A4(new_n581), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT72), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n578), .A2(new_n581), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n594), .B1(new_n595), .B2(new_n478), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  AOI211_X1 g412(.A(new_n583), .B(new_n587), .C1(new_n598), .C2(KEYINPUT28), .ZN(new_n599));
  XOR2_X1   g413(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n600));
  NAND2_X1  g414(.A1(new_n589), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT30), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n601), .B(new_n478), .C1(new_n602), .C2(new_n595), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n597), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n587), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT29), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n189), .B1(new_n599), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n583), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n587), .A2(new_n606), .ZN(new_n610));
  AOI22_X1  g424(.A1(new_n578), .A2(new_n581), .B1(new_n490), .B2(new_n477), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n611), .B1(new_n593), .B2(new_n596), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT28), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n609), .B(new_n610), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT76), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(G472), .B1(new_n608), .B2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(G472), .A2(G902), .ZN(new_n618));
  AOI22_X1  g432(.A1(new_n582), .A2(KEYINPUT30), .B1(new_n589), .B2(new_n600), .ZN(new_n619));
  AOI22_X1  g433(.A1(new_n619), .A2(new_n478), .B1(new_n593), .B2(new_n596), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n586), .B(new_n220), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT73), .B(KEYINPUT31), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n620), .A2(KEYINPUT74), .A3(new_n621), .A4(new_n622), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n597), .A2(new_n621), .A3(new_n603), .A4(new_n622), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT74), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n597), .A2(new_n621), .A3(new_n603), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(KEYINPUT31), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n623), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n598), .A2(KEYINPUT28), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n621), .B1(new_n630), .B2(new_n609), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n618), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT32), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OAI211_X1 g448(.A(KEYINPUT32), .B(new_n618), .C1(new_n629), .C2(new_n631), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n617), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n504), .A2(new_n529), .A3(new_n577), .A4(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G101), .ZN(G3));
  OAI21_X1  g452(.A(new_n189), .B1(new_n629), .B2(new_n631), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(G472), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n640), .A2(new_n632), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n294), .A2(new_n576), .ZN(new_n642));
  OAI211_X1 g456(.A(new_n428), .B(new_n361), .C1(new_n501), .C2(new_n502), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT33), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n644), .B1(new_n340), .B2(new_n343), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n350), .A2(new_n351), .A3(KEYINPUT33), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n505), .A2(new_n345), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n344), .A2(new_n345), .ZN(new_n649));
  INV_X1    g463(.A(new_n423), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n421), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n648), .A2(new_n649), .B1(new_n651), .B2(new_n410), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n643), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n641), .A2(new_n642), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT34), .B(G104), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT95), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n655), .B(new_n657), .ZN(G6));
  INV_X1    g472(.A(KEYINPUT96), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n410), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n409), .A2(KEYINPUT96), .A3(G475), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n355), .A2(new_n651), .A3(new_n660), .A4(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n643), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n641), .A2(new_n642), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT97), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT35), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G107), .ZN(G9));
  NOR2_X1   g481(.A1(new_n533), .A2(KEYINPUT36), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n563), .B(new_n668), .Z(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n574), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n671));
  NOR4_X1   g485(.A1(new_n560), .A2(new_n564), .A3(KEYINPUT25), .A4(new_n505), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT98), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n572), .A2(KEYINPUT98), .A3(new_n670), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n640), .A2(new_n677), .A3(new_n632), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(KEYINPUT99), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT99), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n640), .A2(new_n677), .A3(new_n680), .A4(new_n632), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n679), .A2(new_n504), .A3(new_n529), .A4(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(KEYINPUT37), .B(G110), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G12));
  AOI22_X1  g498(.A1(new_n519), .A2(new_n518), .B1(new_n675), .B2(new_n676), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n347), .A2(new_n354), .ZN(new_n686));
  INV_X1    g500(.A(G900), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n357), .B1(new_n358), .B2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n651), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n660), .A2(new_n661), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n686), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n636), .A2(new_n528), .A3(new_n685), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(KEYINPUT100), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G128), .ZN(G30));
  NAND2_X1  g509(.A1(G472), .A2(G902), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n627), .A2(G472), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n612), .A2(new_n621), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  XOR2_X1   g513(.A(new_n699), .B(KEYINPUT101), .Z(new_n700));
  NAND3_X1  g514(.A1(new_n700), .A2(new_n634), .A3(new_n635), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n501), .A2(new_n502), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(KEYINPUT38), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n651), .A2(new_n410), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(new_n355), .A3(new_n428), .ZN(new_n706));
  OR2_X1    g520(.A1(new_n677), .A2(new_n706), .ZN(new_n707));
  OR3_X1    g521(.A1(new_n702), .A2(new_n704), .A3(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(new_n688), .B(KEYINPUT39), .Z(new_n709));
  NAND2_X1  g523(.A1(new_n520), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT40), .ZN(new_n711));
  OR2_X1    g525(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G143), .ZN(G45));
  INV_X1    g527(.A(new_n528), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n652), .A2(new_n689), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(new_n636), .A3(new_n685), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G146), .ZN(G48));
  OAI21_X1  g532(.A(new_n189), .B1(new_n273), .B2(new_n281), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(G469), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n282), .ZN(new_n721));
  INV_X1    g535(.A(new_n291), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n636), .A2(new_n577), .A3(new_n654), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT41), .B(G113), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G15));
  NAND4_X1  g540(.A1(new_n636), .A2(new_n577), .A3(new_n663), .A4(new_n723), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G116), .ZN(G18));
  AND2_X1   g542(.A1(new_n677), .A2(new_n425), .ZN(new_n729));
  INV_X1    g543(.A(new_n723), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n714), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n729), .A2(new_n731), .A3(new_n636), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G119), .ZN(G21));
  NOR2_X1   g547(.A1(new_n730), .A2(new_n360), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n609), .B1(new_n612), .B2(new_n613), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n587), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n736), .A2(new_n623), .A3(new_n628), .A4(new_n626), .ZN(new_n737));
  AOI22_X1  g551(.A1(new_n639), .A2(G472), .B1(new_n618), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n703), .A2(new_n706), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n734), .A2(new_n738), .A3(new_n739), .A4(new_n577), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G122), .ZN(G24));
  INV_X1    g555(.A(KEYINPUT102), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n742), .B1(new_n652), .B2(new_n689), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n648), .A2(new_n649), .ZN(new_n744));
  AND4_X1   g558(.A1(new_n742), .A2(new_n744), .A3(new_n705), .A4(new_n689), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n731), .A2(new_n746), .A3(new_n677), .A4(new_n738), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G125), .ZN(G27));
  NOR2_X1   g562(.A1(new_n288), .A2(KEYINPUT103), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT103), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n272), .A2(new_n194), .ZN(new_n751));
  AOI22_X1  g565(.A1(new_n751), .A2(new_n267), .B1(new_n284), .B2(new_n193), .ZN(new_n752));
  OAI21_X1  g566(.A(G469), .B1(new_n752), .B2(G902), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n750), .B1(new_n753), .B2(new_n282), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n291), .B1(new_n749), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n526), .A2(new_n428), .A3(new_n527), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n757), .A2(new_n746), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n636), .A2(KEYINPUT104), .A3(new_n577), .ZN(new_n759));
  AOI21_X1  g573(.A(KEYINPUT104), .B1(new_n636), .B2(new_n577), .ZN(new_n760));
  OAI211_X1 g574(.A(KEYINPUT42), .B(new_n758), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n636), .A2(new_n757), .A3(new_n577), .A4(new_n746), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT42), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G131), .ZN(G33));
  NAND4_X1  g580(.A1(new_n636), .A2(new_n757), .A3(new_n577), .A4(new_n692), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G134), .ZN(G36));
  NAND2_X1  g582(.A1(new_n285), .A2(new_n286), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n188), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n771), .B1(new_n770), .B2(new_n769), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(KEYINPUT46), .A3(new_n283), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(KEYINPUT105), .ZN(new_n774));
  AOI21_X1  g588(.A(KEYINPUT46), .B1(new_n772), .B2(new_n283), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n775), .A2(new_n515), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n722), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n709), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT106), .ZN(new_n779));
  INV_X1    g593(.A(new_n756), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT43), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n648), .A2(new_n649), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n782), .A2(new_n705), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT107), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n781), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  OAI211_X1 g599(.A(KEYINPUT107), .B(KEYINPUT43), .C1(new_n782), .C2(new_n705), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n677), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT44), .ZN(new_n789));
  OR3_X1    g603(.A1(new_n788), .A2(new_n789), .A3(new_n641), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n789), .B1(new_n788), .B2(new_n641), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n779), .A2(new_n780), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G137), .ZN(G39));
  INV_X1    g607(.A(KEYINPUT47), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n777), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n777), .A2(new_n794), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR4_X1   g611(.A1(new_n636), .A2(new_n577), .A3(new_n715), .A4(new_n756), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G140), .ZN(G42));
  NAND2_X1  g614(.A1(new_n356), .A2(new_n191), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT120), .ZN(new_n802));
  OAI22_X1  g616(.A1(new_n795), .A2(new_n796), .B1(new_n291), .B2(new_n721), .ZN(new_n803));
  AND4_X1   g617(.A1(new_n357), .A2(new_n787), .A3(new_n577), .A4(new_n738), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n804), .A2(new_n780), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  OR2_X1    g620(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n704), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n723), .A2(new_n427), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT115), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n804), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n804), .A2(new_n811), .A3(KEYINPUT116), .A4(KEYINPUT50), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AND4_X1   g630(.A1(new_n357), .A2(new_n787), .A3(new_n723), .A4(new_n780), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n817), .A2(new_n677), .A3(new_n738), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n780), .A2(new_n357), .A3(new_n577), .A4(new_n723), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n820));
  OR3_X1    g634(.A1(new_n701), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n820), .B1(new_n701), .B2(new_n819), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n744), .A2(new_n705), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n806), .A2(new_n816), .A3(new_n818), .A4(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT51), .ZN(new_n826));
  OR2_X1    g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n825), .A2(KEYINPUT118), .A3(new_n826), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT118), .B1(new_n825), .B2(new_n826), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n821), .A2(new_n822), .A3(new_n652), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n804), .A2(new_n731), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n831), .A2(G952), .A3(new_n191), .A4(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n817), .B1(new_n759), .B2(new_n760), .ZN(new_n834));
  OR2_X1    g648(.A1(new_n834), .A2(KEYINPUT48), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(KEYINPUT48), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n833), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  XOR2_X1   g651(.A(new_n837), .B(KEYINPUT119), .Z(new_n838));
  OAI21_X1  g652(.A(new_n802), .B1(new_n830), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n825), .A2(new_n826), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT118), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n825), .A2(KEYINPUT118), .A3(new_n826), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n837), .B(KEYINPUT119), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n844), .A2(KEYINPUT120), .A3(new_n845), .A4(new_n827), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n839), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n757), .A2(new_n746), .A3(new_n677), .A4(new_n738), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n767), .A2(new_n848), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n690), .A2(new_n355), .A3(new_n691), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n703), .A2(new_n850), .A3(KEYINPUT110), .A4(new_n428), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT110), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n688), .B1(new_n650), .B2(new_n421), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n686), .A2(new_n660), .A3(new_n661), .A4(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n852), .B1(new_n756), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n856), .A2(new_n636), .A3(new_n685), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(KEYINPUT111), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT111), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n856), .A2(new_n859), .A3(new_n636), .A4(new_n685), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n849), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT109), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n355), .A2(new_n410), .A3(new_n651), .ZN(new_n863));
  OR3_X1    g677(.A1(new_n643), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n862), .B1(new_n643), .B2(new_n863), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n864), .A2(new_n641), .A3(new_n642), .A4(new_n865), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n682), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n637), .A2(KEYINPUT108), .A3(new_n655), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n637), .A2(new_n655), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT108), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n861), .A2(new_n867), .A3(new_n868), .A4(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT114), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n755), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n673), .A2(new_n688), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n701), .A2(new_n739), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n877), .A2(new_n693), .A3(new_n747), .A4(new_n717), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT52), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n879), .A2(KEYINPUT112), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n879), .A2(KEYINPUT112), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n878), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n882), .B1(new_n879), .B2(new_n878), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n682), .A2(new_n866), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT108), .B1(new_n637), .B2(new_n655), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n886), .A2(KEYINPUT114), .A3(new_n868), .A4(new_n861), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT53), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n724), .A2(new_n727), .A3(new_n732), .A4(new_n740), .ZN(new_n889));
  AOI211_X1 g703(.A(new_n888), .B(new_n889), .C1(new_n761), .C2(new_n764), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n874), .A2(new_n883), .A3(new_n887), .A4(new_n890), .ZN(new_n891));
  XNOR2_X1  g705(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n889), .B1(new_n761), .B2(new_n764), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n893), .A2(new_n886), .A3(new_n868), .A4(new_n861), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n878), .B(KEYINPUT52), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n892), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT54), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n891), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n894), .A2(new_n895), .A3(new_n892), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n886), .A2(new_n868), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n900), .A2(new_n883), .A3(new_n893), .A4(new_n861), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n899), .B1(new_n888), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n898), .B1(new_n902), .B2(new_n897), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n801), .B1(new_n847), .B2(new_n903), .ZN(new_n904));
  AND4_X1   g718(.A1(new_n291), .A2(new_n577), .A3(new_n783), .A4(new_n428), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n721), .B(KEYINPUT49), .Z(new_n906));
  NAND4_X1  g720(.A1(new_n702), .A2(new_n704), .A3(new_n905), .A4(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n904), .A2(new_n907), .ZN(G75));
  NAND2_X1  g722(.A1(new_n891), .A2(new_n896), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n505), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n910), .A2(new_n488), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n911), .A2(KEYINPUT56), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n497), .A2(new_n498), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(new_n499), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT55), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n191), .A2(G952), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  XOR2_X1   g732(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n919));
  NAND2_X1  g733(.A1(new_n915), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n918), .B1(new_n911), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n916), .A2(new_n921), .ZN(G51));
  NAND2_X1  g736(.A1(new_n909), .A2(KEYINPUT54), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n898), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n283), .B(KEYINPUT57), .Z(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n926), .B1(new_n273), .B2(new_n281), .ZN(new_n927));
  OR2_X1    g741(.A1(new_n910), .A2(new_n772), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n917), .B1(new_n927), .B2(new_n928), .ZN(G54));
  AND4_X1   g743(.A1(KEYINPUT58), .A2(new_n909), .A3(G475), .A4(new_n505), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n918), .B1(new_n930), .B2(new_n418), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n931), .B1(new_n418), .B2(new_n930), .ZN(G60));
  AND2_X1   g746(.A1(new_n645), .A2(new_n646), .ZN(new_n933));
  NAND2_X1  g747(.A1(G478), .A2(G902), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT59), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n924), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n933), .B1(new_n903), .B2(new_n935), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n936), .A2(new_n937), .A3(new_n917), .ZN(G63));
  INV_X1    g752(.A(KEYINPUT61), .ZN(new_n939));
  NAND2_X1  g753(.A1(G217), .A2(G902), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT60), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(new_n891), .B2(new_n896), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n669), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n918), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n942), .A2(new_n573), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n939), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n941), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n909), .A2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n573), .ZN(new_n949));
  AOI21_X1  g763(.A(KEYINPUT122), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT122), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n942), .A2(new_n951), .A3(new_n573), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n943), .A2(KEYINPUT61), .A3(new_n918), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(KEYINPUT123), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n948), .A2(KEYINPUT122), .A3(new_n949), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n951), .B1(new_n942), .B2(new_n573), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT123), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n959), .A2(new_n960), .A3(new_n954), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n946), .B1(new_n956), .B2(new_n961), .ZN(G66));
  INV_X1    g776(.A(new_n889), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n900), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(G224), .A2(G953), .ZN(new_n965));
  OAI22_X1  g779(.A1(new_n964), .A2(G953), .B1(new_n359), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n913), .B1(G898), .B2(new_n191), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n966), .B(new_n967), .Z(G69));
  NAND3_X1  g782(.A1(new_n747), .A2(new_n693), .A3(new_n717), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n712), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n971), .A2(KEYINPUT62), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT124), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n971), .A2(KEYINPUT62), .ZN(new_n974));
  INV_X1    g788(.A(new_n710), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n756), .B1(new_n653), .B2(new_n863), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n975), .A2(new_n577), .A3(new_n636), .A4(new_n976), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n974), .A2(new_n792), .A3(new_n799), .A4(new_n977), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n973), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(new_n191), .ZN(new_n980));
  NAND3_X1  g794(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n619), .B(new_n413), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n792), .A2(new_n767), .A3(new_n799), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n759), .A2(new_n760), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n985), .A2(new_n703), .A3(new_n706), .ZN(new_n986));
  AOI22_X1  g800(.A1(new_n779), .A2(new_n986), .B1(new_n761), .B2(new_n764), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n984), .A2(new_n970), .A3(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT125), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n984), .A2(new_n987), .A3(KEYINPUT125), .A4(new_n970), .ZN(new_n991));
  AOI21_X1  g805(.A(G953), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n687), .A2(new_n191), .A3(G227), .ZN(new_n993));
  OR2_X1    g807(.A1(new_n982), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n983), .B1(new_n992), .B2(new_n994), .ZN(G72));
  XOR2_X1   g809(.A(new_n696), .B(KEYINPUT63), .Z(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(new_n964), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n997), .B1(new_n979), .B2(new_n998), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n620), .B(KEYINPUT126), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(new_n621), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n918), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  OR2_X1    g816(.A1(new_n1000), .A2(new_n621), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n990), .A2(new_n998), .A3(new_n991), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1003), .B1(new_n1004), .B2(new_n996), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n997), .B1(new_n605), .B2(new_n627), .ZN(new_n1006));
  XOR2_X1   g820(.A(new_n1006), .B(KEYINPUT127), .Z(new_n1007));
  NOR2_X1   g821(.A1(new_n902), .A2(new_n1007), .ZN(new_n1008));
  NOR3_X1   g822(.A1(new_n1002), .A2(new_n1005), .A3(new_n1008), .ZN(G57));
endmodule


