//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 0 1 0 1 0 0 0 1 1 0 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 1 1 0 1 0 0 0 0 0 0 0 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1282, new_n1283, new_n1284, new_n1285,
    new_n1286, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI211_X1 g0005(.A(G50), .B(G77), .C1(new_n204), .C2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n204), .A2(new_n205), .ZN(new_n215));
  INV_X1    g0015(.A(G50), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n209), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AND2_X1   g0020(.A1(KEYINPUT65), .A2(G77), .ZN(new_n221));
  NOR2_X1   g0021(.A1(KEYINPUT65), .A2(G77), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  AND2_X1   g0024(.A1(new_n224), .A2(G244), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G58), .A2(G232), .ZN(new_n229));
  NAND4_X1  g0029(.A1(new_n226), .A2(new_n227), .A3(new_n228), .A4(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n211), .B1(new_n225), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n214), .B(new_n220), .C1(KEYINPUT1), .C2(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XNOR2_X1  g0042(.A(G68), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n202), .ZN(new_n244));
  XOR2_X1   g0044(.A(KEYINPUT66), .B(G50), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  XNOR2_X1  g0050(.A(KEYINPUT3), .B(G33), .ZN(new_n251));
  INV_X1    g0051(.A(G1698), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n251), .A2(G222), .A3(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n251), .A2(G223), .A3(G1698), .ZN(new_n254));
  OAI211_X1 g0054(.A(new_n253), .B(new_n254), .C1(new_n223), .C2(new_n251), .ZN(new_n255));
  AND2_X1   g0055(.A1(G33), .A2(G41), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n256), .A2(new_n218), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(G274), .B1(new_n256), .B2(new_n218), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AND2_X1   g0061(.A1(G1), .A2(G13), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G33), .A2(G41), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n260), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n261), .B1(G226), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n258), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT67), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n258), .A2(KEYINPUT67), .A3(new_n267), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n270), .A2(G200), .A3(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n218), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n209), .B1(new_n215), .B2(new_n216), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT8), .B(G58), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n209), .A2(G33), .ZN(new_n277));
  INV_X1    g0077(.A(G150), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G20), .A2(G33), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  OAI22_X1  g0080(.A1(new_n276), .A2(new_n277), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n274), .B1(new_n275), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n284), .A2(new_n274), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n216), .B1(new_n208), .B2(G20), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n285), .A2(new_n286), .B1(new_n216), .B2(new_n284), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n282), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g0088(.A(new_n288), .B(KEYINPUT9), .ZN(new_n289));
  AND2_X1   g0089(.A1(new_n272), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT69), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n270), .A2(new_n271), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G190), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n290), .A2(new_n291), .A3(KEYINPUT10), .A4(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n271), .ZN(new_n295));
  AOI21_X1  g0095(.A(KEYINPUT67), .B1(new_n258), .B2(new_n267), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G190), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n272), .B(new_n289), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n291), .A2(KEYINPUT10), .ZN(new_n300));
  OR2_X1    g0100(.A1(new_n291), .A2(KEYINPUT10), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G179), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n292), .A2(new_n303), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n304), .B(new_n288), .C1(G169), .C2(new_n292), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n294), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n284), .A2(new_n203), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n307), .B(KEYINPUT12), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n279), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n309));
  INV_X1    g0109(.A(G77), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n309), .B1(new_n310), .B2(new_n277), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n311), .A2(KEYINPUT11), .A3(new_n274), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n208), .A2(G20), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n285), .A2(G68), .A3(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n308), .A2(new_n312), .A3(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(KEYINPUT11), .B1(new_n311), .B2(new_n274), .ZN(new_n316));
  OR2_X1    g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT14), .ZN(new_n318));
  INV_X1    g0118(.A(G33), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT3), .ZN(new_n320));
  INV_X1    g0120(.A(G226), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n252), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT3), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G33), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n235), .A2(G1698), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n320), .A2(new_n322), .A3(new_n324), .A4(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(G33), .A2(G97), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT70), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT70), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n326), .A2(new_n330), .A3(new_n327), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n329), .A2(new_n257), .A3(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT13), .ZN(new_n333));
  INV_X1    g0133(.A(G274), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n334), .B1(new_n262), .B2(new_n263), .ZN(new_n335));
  INV_X1    g0135(.A(new_n260), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G238), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n337), .B1(new_n265), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  AND3_X1   g0140(.A1(new_n332), .A2(new_n333), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n333), .B1(new_n332), .B2(new_n340), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n318), .B(G169), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  AND3_X1   g0143(.A1(new_n326), .A2(new_n330), .A3(new_n327), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n330), .B1(new_n326), .B2(new_n327), .ZN(new_n345));
  NOR3_X1   g0145(.A1(new_n344), .A2(new_n345), .A3(new_n264), .ZN(new_n346));
  OAI21_X1  g0146(.A(KEYINPUT13), .B1(new_n346), .B2(new_n339), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n332), .A2(new_n333), .A3(new_n340), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n347), .A2(new_n348), .A3(G179), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n343), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n347), .A2(new_n348), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n318), .B1(new_n351), .B2(G169), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n317), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n341), .A2(new_n342), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n317), .B1(new_n354), .B2(G190), .ZN(new_n355));
  INV_X1    g0155(.A(G200), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n355), .B1(new_n356), .B2(new_n354), .ZN(new_n357));
  XNOR2_X1  g0157(.A(KEYINPUT15), .B(G87), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n358), .A2(new_n277), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n359), .B1(G20), .B2(new_n224), .ZN(new_n360));
  INV_X1    g0160(.A(new_n276), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n279), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n360), .A2(new_n362), .B1(new_n218), .B2(new_n273), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n285), .A2(G77), .A3(new_n313), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(new_n224), .B2(new_n283), .ZN(new_n365));
  OR2_X1    g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n251), .A2(G238), .A3(G1698), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n251), .A2(G232), .A3(new_n252), .ZN(new_n368));
  INV_X1    g0168(.A(G107), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n367), .B(new_n368), .C1(new_n369), .C2(new_n251), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n257), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n261), .B1(G244), .B2(new_n266), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G169), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n366), .B(new_n375), .C1(G179), .C2(new_n373), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n373), .A2(G200), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT68), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n371), .A2(G190), .A3(new_n372), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n363), .A2(new_n365), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT68), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n381), .B1(new_n379), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n353), .A2(new_n357), .A3(new_n376), .A4(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT16), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT73), .B1(new_n319), .B2(KEYINPUT3), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT72), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n323), .B2(G33), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT73), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n391), .A2(new_n323), .A3(G33), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n319), .A2(KEYINPUT72), .A3(KEYINPUT3), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n388), .A2(new_n390), .A3(new_n392), .A4(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT7), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n395), .A2(G20), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n395), .B1(new_n251), .B2(G20), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n203), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(G58), .A2(G68), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n204), .A2(new_n205), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(G20), .ZN(new_n402));
  INV_X1    g0202(.A(G159), .ZN(new_n403));
  NOR3_X1   g0203(.A1(new_n403), .A2(G20), .A3(G33), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n387), .B1(new_n399), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n320), .A2(new_n324), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT7), .B1(new_n408), .B2(new_n209), .ZN(new_n409));
  AOI211_X1 g0209(.A(new_n395), .B(G20), .C1(new_n320), .C2(new_n324), .ZN(new_n410));
  OAI21_X1  g0210(.A(G68), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(KEYINPUT71), .B1(new_n402), .B2(new_n405), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT71), .ZN(new_n413));
  AOI211_X1 g0213(.A(new_n413), .B(new_n404), .C1(new_n401), .C2(G20), .ZN(new_n414));
  OAI211_X1 g0214(.A(KEYINPUT16), .B(new_n411), .C1(new_n412), .C2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n407), .A2(new_n415), .A3(new_n274), .ZN(new_n416));
  INV_X1    g0216(.A(new_n285), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n361), .A2(new_n313), .ZN(new_n418));
  OAI22_X1  g0218(.A1(new_n417), .A2(new_n418), .B1(new_n283), .B2(new_n361), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n416), .A2(new_n420), .ZN(new_n421));
  OR2_X1    g0221(.A1(G223), .A2(G1698), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n321), .A2(G1698), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n251), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(G33), .A2(G87), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n264), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n337), .B1(new_n235), .B2(new_n265), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n374), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  NOR3_X1   g0230(.A1(new_n426), .A2(new_n428), .A3(new_n303), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n421), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT18), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n432), .B1(new_n416), .B2(new_n420), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT18), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n427), .A2(new_n429), .A3(new_n298), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n356), .B1(new_n426), .B2(new_n428), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n416), .A2(new_n420), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT17), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n416), .A2(KEYINPUT17), .A3(new_n420), .A4(new_n441), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n435), .A2(new_n438), .A3(new_n444), .A4(new_n445), .ZN(new_n446));
  NOR3_X1   g0246(.A1(new_n306), .A2(new_n386), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(G33), .A2(G283), .ZN(new_n449));
  INV_X1    g0249(.A(G97), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n449), .B(new_n209), .C1(G33), .C2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(G116), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(G20), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n451), .A2(new_n274), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT20), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n451), .A2(KEYINPUT20), .A3(new_n274), .A4(new_n453), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n283), .A2(new_n452), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n208), .A2(G33), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n283), .A2(new_n460), .A3(new_n218), .A4(new_n273), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n459), .B1(new_n462), .B2(new_n452), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n374), .B1(new_n458), .B2(new_n463), .ZN(new_n464));
  XNOR2_X1  g0264(.A(KEYINPUT77), .B(G303), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n408), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G264), .A2(G1698), .ZN(new_n467));
  INV_X1    g0267(.A(G257), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n467), .B1(new_n468), .B2(G1698), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n251), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT78), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n466), .A2(new_n470), .A3(KEYINPUT78), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n264), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(G45), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(G1), .ZN(new_n477));
  NAND2_X1  g0277(.A1(KEYINPUT5), .A2(G41), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(KEYINPUT5), .A2(G41), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(KEYINPUT74), .B1(new_n481), .B2(new_n259), .ZN(new_n482));
  XNOR2_X1  g0282(.A(KEYINPUT5), .B(G41), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT74), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n335), .A2(new_n483), .A3(new_n484), .A4(new_n477), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n257), .B1(new_n477), .B2(new_n483), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G270), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n464), .B(KEYINPUT21), .C1(new_n475), .C2(new_n489), .ZN(new_n490));
  AND3_X1   g0290(.A1(new_n466), .A2(new_n470), .A3(KEYINPUT78), .ZN(new_n491));
  AOI21_X1  g0291(.A(KEYINPUT78), .B1(new_n466), .B2(new_n470), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n257), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n458), .A2(new_n463), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n482), .A2(new_n485), .B1(new_n487), .B2(G270), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n493), .A2(new_n494), .A3(G179), .A4(new_n495), .ZN(new_n496));
  AND2_X1   g0296(.A1(new_n490), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n493), .A2(new_n495), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n464), .ZN(new_n499));
  XOR2_X1   g0299(.A(KEYINPUT79), .B(KEYINPUT21), .Z(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n498), .A2(G200), .ZN(new_n502));
  INV_X1    g0302(.A(new_n494), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n493), .A2(G190), .A3(new_n495), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n497), .A2(new_n501), .A3(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n283), .A2(G97), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n507), .B1(new_n462), .B2(G97), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT6), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n450), .A2(new_n369), .ZN(new_n511));
  NOR2_X1   g0311(.A1(G97), .A2(G107), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR3_X1   g0313(.A1(new_n510), .A2(new_n450), .A3(G107), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n516), .A2(G20), .B1(G77), .B2(new_n279), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n409), .B1(new_n394), .B2(new_n396), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n517), .B1(new_n518), .B2(new_n369), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n509), .B1(new_n519), .B2(new_n274), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n320), .A2(new_n324), .A3(G244), .A4(new_n252), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT4), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n251), .A2(G250), .A3(G1698), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n523), .A2(new_n449), .A3(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n521), .A2(new_n522), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n257), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n482), .A2(new_n485), .B1(new_n487), .B2(G257), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n527), .A2(new_n298), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(G200), .B1(new_n527), .B2(new_n528), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n520), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n527), .A2(new_n528), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n374), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n369), .B1(new_n397), .B2(new_n398), .ZN(new_n534));
  XNOR2_X1  g0334(.A(G97), .B(G107), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n514), .B1(new_n510), .B2(new_n535), .ZN(new_n536));
  OAI22_X1  g0336(.A1(new_n536), .A2(new_n209), .B1(new_n310), .B2(new_n280), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n274), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n508), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n527), .A2(new_n303), .A3(new_n528), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n533), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n531), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n320), .A2(new_n324), .A3(G244), .A4(G1698), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n320), .A2(new_n324), .A3(G238), .A4(new_n252), .ZN(new_n544));
  NAND2_X1  g0344(.A1(G33), .A2(G116), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(G250), .ZN(new_n547));
  OAI22_X1  g0347(.A1(KEYINPUT75), .A2(new_n547), .B1(new_n476), .B2(G1), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n548), .A2(new_n264), .ZN(new_n549));
  NAND2_X1  g0349(.A1(KEYINPUT75), .A2(G250), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n477), .A2(new_n334), .A3(new_n550), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n546), .A2(new_n257), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n303), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT19), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n209), .B1(new_n327), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(G87), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n512), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n320), .A2(new_n324), .A3(new_n209), .A4(G68), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n554), .B1(new_n277), .B2(new_n450), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n274), .ZN(new_n562));
  INV_X1    g0362(.A(new_n358), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(KEYINPUT76), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT76), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n358), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n462), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n358), .A2(new_n284), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n562), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n553), .B(new_n569), .C1(G169), .C2(new_n552), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n546), .A2(new_n257), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n549), .A2(new_n551), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(G200), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n462), .A2(G87), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n562), .A2(new_n575), .A3(new_n568), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n552), .A2(G190), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n570), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n468), .A2(G1698), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(G250), .B2(G1698), .ZN(new_n581));
  INV_X1    g0381(.A(G294), .ZN(new_n582));
  OAI22_X1  g0382(.A1(new_n581), .A2(new_n408), .B1(new_n319), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n257), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n487), .A2(G264), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n486), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n586), .A2(KEYINPUT81), .A3(new_n356), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n486), .A2(new_n584), .A3(new_n585), .A4(new_n298), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n588), .A2(KEYINPUT81), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n257), .A2(new_n583), .B1(new_n487), .B2(G264), .ZN(new_n590));
  AOI21_X1  g0390(.A(G200), .B1(new_n590), .B2(new_n486), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n587), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n320), .A2(new_n324), .A3(new_n209), .A4(G87), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(KEYINPUT22), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT22), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n251), .A2(new_n595), .A3(new_n209), .A4(G87), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(KEYINPUT23), .B1(new_n209), .B2(G107), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT23), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n599), .A2(new_n369), .A3(G20), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n209), .A2(G33), .A3(G116), .ZN(new_n601));
  NAND2_X1  g0401(.A1(KEYINPUT80), .A2(KEYINPUT24), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n598), .A2(new_n600), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT80), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT24), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n597), .A2(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n606), .ZN(new_n608));
  AOI211_X1 g0408(.A(new_n608), .B(new_n603), .C1(new_n594), .C2(new_n596), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n274), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n284), .A2(KEYINPUT25), .A3(new_n369), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT25), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n612), .B1(new_n283), .B2(G107), .ZN(new_n613));
  AOI22_X1  g0413(.A1(G107), .A2(new_n462), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n579), .B1(new_n592), .B2(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n586), .A2(G179), .ZN(new_n618));
  AOI21_X1  g0418(.A(G169), .B1(new_n590), .B2(new_n486), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n615), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n506), .A2(new_n542), .A3(new_n617), .A4(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n448), .A2(new_n622), .ZN(G372));
  NAND2_X1  g0423(.A1(new_n444), .A2(new_n445), .ZN(new_n624));
  INV_X1    g0424(.A(new_n376), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n357), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n624), .B1(new_n626), .B2(new_n353), .ZN(new_n627));
  XNOR2_X1  g0427(.A(new_n436), .B(KEYINPUT18), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n302), .B(new_n294), .C1(new_n627), .C2(new_n629), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n630), .A2(new_n305), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n497), .A2(new_n621), .A3(new_n501), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n632), .A2(new_n542), .A3(new_n617), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n533), .A2(new_n539), .A3(new_n540), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n570), .A2(new_n578), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n634), .A2(new_n635), .A3(KEYINPUT26), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT26), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n637), .B1(new_n541), .B2(new_n579), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n633), .A2(new_n570), .A3(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n631), .B1(new_n448), .B2(new_n641), .ZN(G369));
  NAND2_X1  g0442(.A1(new_n497), .A2(new_n501), .ZN(new_n643));
  INV_X1    g0443(.A(G13), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n644), .A2(G1), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n209), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT27), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n645), .A2(new_n648), .A3(new_n209), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n647), .A2(G213), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g0450(.A(new_n650), .B(KEYINPUT82), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(G343), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n652), .A2(new_n503), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n643), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n497), .A2(new_n501), .A3(new_n505), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n654), .B1(new_n655), .B2(new_n653), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(G330), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n652), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n621), .A2(new_n660), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n588), .A2(KEYINPUT81), .B1(new_n586), .B2(new_n356), .ZN(new_n662));
  INV_X1    g0462(.A(new_n587), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n610), .B(new_n614), .C1(new_n662), .C2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n616), .B2(new_n652), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n661), .B1(new_n665), .B2(new_n621), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n659), .A2(new_n666), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n499), .A2(new_n500), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n490), .A2(new_n496), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n652), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT83), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n643), .A2(KEYINPUT83), .A3(new_n652), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n661), .B1(new_n674), .B2(new_n666), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n667), .A2(new_n675), .ZN(G399));
  INV_X1    g0476(.A(new_n212), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(G41), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n217), .ZN(new_n679));
  INV_X1    g0479(.A(new_n678), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n557), .A2(G116), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(G1), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n679), .B1(new_n682), .B2(KEYINPUT84), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n683), .B1(KEYINPUT84), .B2(new_n682), .ZN(new_n684));
  XOR2_X1   g0484(.A(new_n684), .B(KEYINPUT28), .Z(new_n685));
  NAND3_X1  g0485(.A1(new_n493), .A2(G179), .A3(new_n495), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT85), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n532), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n493), .A2(KEYINPUT85), .A3(G179), .A4(new_n495), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n590), .A2(new_n552), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n688), .A2(new_n689), .A3(new_n690), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g0492(.A(KEYINPUT86), .B(KEYINPUT30), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n527), .A2(KEYINPUT30), .A3(new_n528), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n688), .A2(new_n690), .A3(new_n691), .A4(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(G179), .B1(new_n590), .B2(new_n486), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n498), .A2(new_n532), .A3(new_n697), .A4(new_n573), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  OAI211_X1 g0499(.A(KEYINPUT31), .B(new_n660), .C1(new_n694), .C2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n622), .B2(new_n660), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n696), .A2(new_n698), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n692), .A2(new_n693), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n652), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(KEYINPUT31), .ZN(new_n705));
  OAI21_X1  g0505(.A(G330), .B1(new_n701), .B2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT88), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT87), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n709), .B1(new_n640), .B2(new_n652), .ZN(new_n710));
  AOI21_X1  g0510(.A(KEYINPUT88), .B1(new_n640), .B2(new_n652), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT29), .ZN(new_n712));
  OAI22_X1  g0512(.A1(new_n708), .A2(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n640), .A2(new_n652), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(KEYINPUT87), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n715), .A2(KEYINPUT88), .A3(KEYINPUT29), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n707), .B1(new_n713), .B2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n685), .B1(new_n717), .B2(G1), .ZN(G364));
  NOR2_X1   g0518(.A1(new_n644), .A2(G20), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n208), .B1(new_n719), .B2(G45), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n678), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n659), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(G330), .B2(new_n656), .ZN(new_n724));
  NOR2_X1   g0524(.A1(G13), .A2(G33), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G20), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n218), .B1(G20), .B2(new_n374), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n677), .A2(new_n251), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n732), .B1(new_n217), .B2(new_n476), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(KEYINPUT89), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n734), .B1(G45), .B2(new_n246), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n733), .A2(KEYINPUT89), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n677), .A2(new_n408), .ZN(new_n738));
  AOI22_X1  g0538(.A1(new_n738), .A2(G355), .B1(new_n452), .B2(new_n677), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n730), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n728), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G179), .A2(G200), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n209), .B1(new_n742), .B2(G190), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n298), .A2(new_n356), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n209), .A2(G179), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(G303), .ZN(new_n747));
  OAI221_X1 g0547(.A(new_n408), .B1(new_n743), .B2(new_n582), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n209), .A2(new_n303), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n750), .A2(new_n298), .A3(G200), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(G322), .ZN(new_n753));
  INV_X1    g0553(.A(G329), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n742), .A2(G20), .A3(new_n298), .ZN(new_n755));
  OAI22_X1  g0555(.A1(new_n752), .A2(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NOR3_X1   g0556(.A1(new_n750), .A2(G190), .A3(G200), .ZN(new_n757));
  AOI211_X1 g0557(.A(new_n748), .B(new_n756), .C1(G311), .C2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT91), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n356), .A2(G190), .ZN(new_n760));
  AND3_X1   g0560(.A1(new_n749), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n759), .B1(new_n749), .B2(new_n760), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  XNOR2_X1  g0564(.A(KEYINPUT33), .B(G317), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n745), .A2(new_n760), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n767), .A2(KEYINPUT90), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(KEYINPUT90), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G283), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n749), .A2(new_n744), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT92), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G326), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n758), .A2(new_n766), .A3(new_n772), .A4(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n757), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n778), .A2(new_n223), .B1(new_n746), .B2(new_n556), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(G58), .B2(new_n751), .ZN(new_n780));
  INV_X1    g0580(.A(new_n755), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G159), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT32), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n743), .A2(new_n450), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n251), .B1(new_n773), .B2(new_n216), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n764), .A2(G68), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n770), .A2(new_n369), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n780), .A2(new_n786), .A3(new_n787), .A4(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n741), .B1(new_n777), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n722), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n740), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n727), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n793), .B1(new_n656), .B2(new_n794), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n724), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(G396));
  NAND2_X1  g0597(.A1(new_n660), .A2(new_n366), .ZN(new_n798));
  INV_X1    g0598(.A(new_n379), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n799), .B1(new_n377), .B2(KEYINPUT68), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n376), .B(new_n798), .C1(new_n800), .C2(new_n383), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT93), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n385), .A2(KEYINPUT93), .A3(new_n376), .A4(new_n798), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n625), .A2(new_n660), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT94), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n714), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n803), .A2(new_n804), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n640), .A2(new_n652), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n722), .B1(new_n812), .B2(new_n706), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n706), .B2(new_n812), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n728), .A2(new_n725), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n722), .B1(G77), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n773), .A2(new_n747), .ZN(new_n818));
  INV_X1    g0618(.A(G311), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n746), .A2(new_n369), .B1(new_n755), .B2(new_n819), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n818), .B(new_n820), .C1(G116), .C2(new_n757), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n771), .A2(G87), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n251), .B(new_n784), .C1(new_n751), .C2(G294), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n764), .A2(G283), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n821), .A2(new_n822), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n773), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n757), .A2(G159), .B1(new_n826), .B2(G137), .ZN(new_n827));
  INV_X1    g0627(.A(G143), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n827), .B1(new_n828), .B2(new_n752), .C1(new_n763), .C2(new_n278), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT34), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G132), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n251), .B1(new_n755), .B2(new_n832), .C1(new_n746), .C2(new_n216), .ZN(new_n833));
  INV_X1    g0633(.A(new_n743), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n833), .B1(G58), .B2(new_n834), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n831), .B(new_n835), .C1(new_n203), .C2(new_n770), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n829), .A2(new_n830), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n825), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n817), .B1(new_n838), .B2(new_n728), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n806), .B2(new_n726), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n814), .A2(new_n840), .ZN(G384));
  OR2_X1    g0641(.A1(new_n516), .A2(KEYINPUT35), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n516), .A2(KEYINPUT35), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n842), .A2(G116), .A3(new_n219), .A4(new_n843), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT36), .Z(new_n845));
  NAND3_X1  g0645(.A1(new_n217), .A2(new_n224), .A3(new_n400), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n216), .A2(G68), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n208), .B(G13), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n421), .A2(new_n651), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT37), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n434), .A2(new_n850), .A3(new_n851), .A4(new_n442), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n411), .B1(new_n412), .B2(new_n414), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n387), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n854), .A2(new_n274), .A3(new_n415), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n432), .B1(new_n855), .B2(new_n420), .ZN(new_n856));
  INV_X1    g0656(.A(new_n651), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n857), .B1(new_n855), .B2(new_n420), .ZN(new_n858));
  AND3_X1   g0658(.A1(new_n416), .A2(new_n420), .A3(new_n441), .ZN(new_n859));
  NOR3_X1   g0659(.A1(new_n856), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n852), .B1(new_n860), .B2(new_n851), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n446), .A2(new_n858), .ZN(new_n862));
  AND3_X1   g0662(.A1(new_n861), .A2(new_n862), .A3(KEYINPUT38), .ZN(new_n863));
  AOI21_X1  g0663(.A(KEYINPUT38), .B1(new_n861), .B2(new_n862), .ZN(new_n864));
  OAI21_X1  g0664(.A(KEYINPUT95), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT38), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n858), .A2(new_n859), .ZN(new_n867));
  INV_X1    g0667(.A(new_n856), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n851), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n852), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n858), .ZN(new_n872));
  INV_X1    g0672(.A(new_n624), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n872), .B1(new_n628), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n866), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT95), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n861), .A2(new_n862), .A3(KEYINPUT38), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n865), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n660), .A2(new_n317), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n353), .A2(new_n357), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n880), .B1(new_n353), .B2(new_n357), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n806), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT97), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n704), .B2(KEYINPUT31), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n660), .B1(new_n694), .B2(new_n699), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT31), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n886), .A2(KEYINPUT97), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n664), .A2(new_n635), .A3(new_n531), .A4(new_n541), .ZN(new_n890));
  INV_X1    g0690(.A(new_n621), .ZN(new_n891));
  NOR3_X1   g0691(.A1(new_n890), .A2(new_n655), .A3(new_n891), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n892), .A2(new_n652), .B1(new_n704), .B2(KEYINPUT31), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n883), .B1(new_n889), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT40), .B1(new_n879), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n434), .A2(new_n850), .A3(new_n442), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(KEYINPUT37), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n897), .A2(KEYINPUT96), .A3(new_n852), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n857), .B1(new_n416), .B2(new_n420), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n446), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT96), .B1(new_n897), .B2(new_n852), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n866), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n877), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT97), .B1(new_n886), .B2(new_n887), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n703), .A2(new_n696), .A3(new_n698), .ZN(new_n906));
  AOI211_X1 g0706(.A(new_n884), .B(KEYINPUT31), .C1(new_n906), .C2(new_n660), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n893), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n883), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n908), .A2(new_n909), .A3(KEYINPUT40), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n895), .B1(new_n904), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n908), .A2(new_n447), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n658), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n912), .B2(new_n914), .ZN(new_n916));
  OR2_X1    g0716(.A1(new_n353), .A2(new_n660), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n415), .A2(new_n274), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n419), .B1(new_n918), .B2(new_n854), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n442), .B1(new_n919), .B2(new_n857), .ZN(new_n920));
  OAI21_X1  g0720(.A(KEYINPUT37), .B1(new_n920), .B2(new_n856), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n852), .A2(new_n921), .B1(new_n446), .B2(new_n858), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT39), .B1(new_n922), .B2(KEYINPUT38), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n903), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT39), .B1(new_n863), .B2(new_n864), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n917), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n625), .A2(new_n652), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n811), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n881), .A2(new_n882), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(new_n865), .B2(new_n878), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n628), .A2(new_n651), .ZN(new_n933));
  NOR3_X1   g0733(.A1(new_n926), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n713), .A2(new_n716), .A3(new_n447), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n631), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n934), .B(new_n936), .Z(new_n937));
  NAND2_X1  g0737(.A1(new_n916), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n208), .B2(new_n719), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n916), .A2(new_n937), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n849), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n941), .B(KEYINPUT98), .Z(G367));
  OAI211_X1 g0742(.A(new_n531), .B(new_n541), .C1(new_n520), .C2(new_n652), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n943), .A2(new_n621), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n660), .B1(new_n944), .B2(new_n541), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n674), .A2(new_n666), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n634), .A2(new_n660), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n943), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(KEYINPUT100), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT100), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n674), .A2(new_n666), .A3(new_n952), .A4(new_n949), .ZN(new_n953));
  AND3_X1   g0753(.A1(new_n951), .A2(KEYINPUT42), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(KEYINPUT42), .B1(new_n951), .B2(new_n953), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n946), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n652), .A2(new_n576), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n579), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n570), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(KEYINPUT99), .B(KEYINPUT43), .Z(new_n962));
  NOR2_X1   g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(KEYINPUT43), .B2(new_n961), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n956), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n951), .A2(new_n953), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT42), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n951), .A2(KEYINPUT42), .A3(new_n953), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n945), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(KEYINPUT101), .B1(new_n970), .B2(new_n963), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n963), .B(new_n946), .C1(new_n954), .C2(new_n955), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT101), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n965), .B1(new_n971), .B2(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n667), .A2(new_n950), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n976), .B(new_n965), .C1(new_n971), .C2(new_n974), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n678), .B(KEYINPUT41), .Z(new_n980));
  INV_X1    g0780(.A(KEYINPUT45), .ZN(new_n981));
  INV_X1    g0781(.A(new_n661), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n947), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n981), .B1(new_n983), .B2(new_n950), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n675), .A2(KEYINPUT45), .A3(new_n949), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n983), .A2(KEYINPUT44), .A3(new_n950), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT44), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n675), .B2(new_n949), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n986), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n667), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n674), .A2(new_n666), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n947), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(new_n659), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n986), .A2(new_n990), .A3(new_n667), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n993), .A2(new_n717), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n980), .B1(new_n998), .B2(new_n717), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n978), .B(new_n979), .C1(new_n721), .C2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(G137), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n746), .A2(new_n202), .B1(new_n755), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n834), .A2(G68), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n251), .B(new_n1003), .C1(new_n778), .C2(new_n216), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n1002), .B(new_n1004), .C1(G150), .C2(new_n751), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n771), .A2(new_n224), .B1(G159), .B2(new_n764), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1005), .B(new_n1006), .C1(new_n828), .C2(new_n774), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n775), .A2(G311), .B1(new_n465), .B2(new_n751), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT102), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n251), .B1(new_n781), .B2(G317), .ZN(new_n1010));
  INV_X1    g0810(.A(G283), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1010), .B1(new_n369), .B2(new_n743), .C1(new_n778), .C2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n746), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(G116), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT46), .Z(new_n1015));
  NOR2_X1   g0815(.A1(new_n770), .A2(new_n450), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n763), .A2(new_n582), .ZN(new_n1017));
  OR4_X1    g0817(.A1(new_n1012), .A2(new_n1015), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1007), .B1(new_n1009), .B2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT47), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n728), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n958), .A2(new_n727), .A3(new_n960), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n731), .A2(new_n241), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n730), .B1(new_n677), .B2(new_n563), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n792), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1021), .A2(new_n1022), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1000), .A2(new_n1026), .ZN(G387));
  INV_X1    g0827(.A(new_n681), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n738), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(G107), .B2(new_n212), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n238), .A2(new_n476), .ZN(new_n1031));
  AOI211_X1 g0831(.A(G45), .B(new_n1028), .C1(G68), .C2(G77), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n276), .A2(G50), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT50), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n732), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1030), .B1(new_n1031), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n722), .B1(new_n1036), .B2(new_n730), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT103), .Z(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n666), .B2(new_n794), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT104), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n773), .A2(new_n403), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n251), .B1(new_n1040), .B2(new_n1041), .C1(new_n778), .C2(new_n203), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1013), .A2(new_n224), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n278), .B2(new_n755), .C1(new_n752), .C2(new_n216), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1045), .A2(new_n1016), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n764), .A2(new_n361), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n564), .A2(new_n566), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n834), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1043), .A2(new_n1046), .A3(new_n1047), .A4(new_n1049), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n465), .A2(new_n757), .B1(new_n751), .B2(G317), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n819), .B2(new_n763), .C1(new_n774), .C2(new_n753), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT105), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT48), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n746), .A2(new_n582), .B1(new_n743), .B2(new_n1011), .ZN(new_n1057));
  NOR3_X1   g0857(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(KEYINPUT49), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n251), .B1(new_n781), .B2(G326), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1059), .B(new_n1060), .C1(new_n452), .C2(new_n770), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1058), .A2(KEYINPUT49), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1050), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1039), .B1(new_n1063), .B2(new_n728), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(new_n996), .B2(new_n721), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n717), .A2(new_n996), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n678), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n717), .A2(new_n996), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1065), .B1(new_n1067), .B2(new_n1068), .ZN(G393));
  INV_X1    g0869(.A(new_n997), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n667), .B1(new_n986), .B2(new_n990), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1066), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1072), .A2(new_n998), .A3(new_n678), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n950), .A2(new_n727), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n729), .B1(new_n450), .B2(new_n212), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n731), .B2(new_n249), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n778), .A2(new_n582), .B1(new_n743), .B2(new_n452), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n764), .B2(new_n465), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT106), .Z(new_n1080));
  AOI22_X1  g0880(.A1(new_n751), .A2(G311), .B1(new_n826), .B2(G317), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT52), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n408), .B1(new_n755), .B2(new_n753), .C1(new_n746), .C2(new_n1011), .ZN(new_n1083));
  NOR4_X1   g0883(.A1(new_n1080), .A2(new_n788), .A3(new_n1082), .A4(new_n1083), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n1084), .A2(KEYINPUT107), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(KEYINPUT107), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n751), .A2(G159), .B1(new_n826), .B2(G150), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT51), .Z(new_n1088));
  OAI21_X1  g0888(.A(new_n251), .B1(new_n778), .B2(new_n276), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n746), .A2(new_n203), .B1(new_n755), .B2(new_n828), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n743), .A2(new_n310), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n764), .A2(G50), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1088), .A2(new_n822), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1085), .A2(new_n1086), .A3(new_n1094), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n792), .B(new_n1077), .C1(new_n1095), .C2(new_n728), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n1074), .A2(new_n721), .B1(new_n1075), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT108), .ZN(new_n1098));
  AND3_X1   g0898(.A1(new_n1073), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1098), .B1(new_n1073), .B2(new_n1097), .ZN(new_n1100));
  OR2_X1    g0900(.A1(new_n1099), .A2(new_n1100), .ZN(G390));
  AOI21_X1  g0901(.A(new_n792), .B1(new_n276), .B2(new_n815), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n770), .A2(new_n203), .B1(new_n369), .B2(new_n763), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n251), .B(new_n1091), .C1(G87), .C2(new_n1013), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n751), .A2(G116), .B1(G294), .B2(new_n781), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n757), .A2(G97), .B1(new_n826), .B2(G283), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1103), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(G128), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n752), .A2(new_n832), .B1(new_n773), .B2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(KEYINPUT54), .B(G143), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n778), .A2(new_n1111), .B1(new_n743), .B2(new_n403), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(new_n764), .B2(G137), .ZN(new_n1113));
  XOR2_X1   g0913(.A(new_n1113), .B(KEYINPUT112), .Z(new_n1114));
  INV_X1    g0914(.A(KEYINPUT53), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n746), .B2(new_n278), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1013), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n1110), .B(new_n1114), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(G125), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n251), .B1(new_n1119), .B2(new_n755), .C1(new_n770), .C2(new_n216), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT113), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1108), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n924), .A2(new_n925), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n1102), .B1(new_n741), .B2(new_n1122), .C1(new_n1123), .C2(new_n726), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n917), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(new_n928), .B2(new_n930), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n904), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n908), .A2(new_n909), .A3(G330), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  OAI211_X1 g0931(.A(G330), .B(new_n806), .C1(new_n701), .C2(new_n705), .ZN(new_n1132));
  OR2_X1    g0932(.A1(new_n1132), .A2(new_n929), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1127), .B(new_n1133), .C1(new_n1123), .C2(new_n1126), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1124), .B1(new_n1135), .B2(new_n720), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n658), .B1(new_n889), .B2(new_n893), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n807), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n929), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n928), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1140), .A2(new_n1141), .A3(new_n1133), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT110), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1132), .A2(new_n929), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1129), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1143), .B1(new_n1145), .B2(new_n928), .ZN(new_n1146));
  AOI211_X1 g0946(.A(KEYINPUT110), .B(new_n1141), .C1(new_n1129), .C2(new_n1144), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1142), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT109), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(new_n1138), .B2(new_n447), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1138), .A2(new_n1149), .A3(new_n447), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n936), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1148), .A2(new_n1131), .A3(new_n1134), .A4(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1154), .A2(KEYINPUT111), .A3(new_n678), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1148), .A2(new_n1153), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n1135), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(KEYINPUT111), .B1(new_n1154), .B2(new_n678), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1137), .B1(new_n1158), .B2(new_n1159), .ZN(G378));
  INV_X1    g0960(.A(new_n934), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n651), .A2(new_n288), .ZN(new_n1162));
  XOR2_X1   g0962(.A(new_n306), .B(new_n1162), .Z(new_n1163));
  XNOR2_X1  g0963(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1164));
  XOR2_X1   g0964(.A(new_n1163), .B(new_n1164), .Z(new_n1165));
  NOR3_X1   g0965(.A1(new_n863), .A2(new_n864), .A3(KEYINPUT95), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n876), .B1(new_n875), .B2(new_n877), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n894), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT40), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n658), .B1(new_n911), .B2(new_n904), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1165), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT96), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n859), .A2(new_n436), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n851), .B1(new_n1174), .B2(new_n850), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1173), .B1(new_n1175), .B2(new_n870), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1176), .A2(new_n900), .A3(new_n898), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n863), .B1(new_n866), .B2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(G330), .B1(new_n910), .B2(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1163), .B(new_n1164), .ZN(new_n1180));
  NOR3_X1   g0980(.A1(new_n895), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1161), .B1(new_n1172), .B2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1170), .A2(new_n1171), .A3(new_n1165), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1180), .B1(new_n895), .B2(new_n1179), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1183), .A2(new_n1184), .A3(new_n934), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1182), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(new_n721), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n771), .A2(G58), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1048), .A2(new_n757), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1188), .B(new_n1189), .C1(new_n450), .C2(new_n763), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n751), .A2(G107), .B1(G283), .B2(new_n781), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n452), .B2(new_n773), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n251), .A2(G41), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1044), .A2(new_n1003), .A3(new_n1193), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n1190), .A2(new_n1192), .A3(new_n1194), .ZN(new_n1195));
  XOR2_X1   g0995(.A(new_n1195), .B(KEYINPUT114), .Z(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(KEYINPUT58), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(G33), .A2(G41), .ZN(new_n1198));
  NOR3_X1   g0998(.A1(new_n1193), .A2(G50), .A3(new_n1198), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n752), .A2(new_n1109), .B1(new_n746), .B2(new_n1111), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n778), .A2(new_n1001), .B1(new_n773), .B2(new_n1119), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1200), .B(new_n1201), .C1(G150), .C2(new_n834), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n832), .B2(new_n763), .ZN(new_n1203));
  OR2_X1    g1003(.A1(new_n1203), .A2(KEYINPUT59), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n781), .A2(G124), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1198), .B(new_n1205), .C1(new_n770), .C2(new_n403), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(new_n1203), .B2(KEYINPUT59), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1199), .B1(new_n1204), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1197), .A2(new_n1208), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1196), .A2(KEYINPUT58), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n728), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n792), .B1(new_n216), .B2(new_n815), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1211), .B(new_n1212), .C1(new_n1165), .C2(new_n726), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1187), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1141), .B1(new_n1132), .B2(new_n929), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n929), .B2(new_n1139), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n894), .A2(G330), .B1(new_n929), .B2(new_n1132), .ZN(new_n1218));
  OAI21_X1  g1018(.A(KEYINPUT110), .B1(new_n1218), .B2(new_n1141), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1145), .A2(new_n1143), .A3(new_n928), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1217), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1153), .B1(new_n1135), .B2(new_n1221), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n1183), .A2(new_n1184), .A3(new_n934), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n934), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1222), .B(KEYINPUT57), .C1(new_n1223), .C2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(KEYINPUT57), .B1(new_n1186), .B2(new_n1222), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT115), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n678), .B(new_n1225), .C1(new_n1226), .C2(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1222), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT57), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1229), .A2(new_n1227), .A3(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1215), .B1(new_n1228), .B2(new_n1232), .ZN(G375));
  OAI21_X1  g1033(.A(KEYINPUT116), .B1(new_n1148), .B2(new_n1153), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n980), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT116), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1152), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n631), .B(new_n935), .C1(new_n1237), .C2(new_n1150), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1221), .A2(new_n1236), .A3(new_n1238), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1234), .A2(new_n1235), .A3(new_n1239), .A4(new_n1156), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n722), .B1(G68), .B2(new_n816), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n752), .A2(new_n1011), .B1(new_n778), .B2(new_n369), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(G97), .B2(new_n1013), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n826), .A2(G294), .B1(G303), .B2(new_n781), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n764), .A2(G116), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1243), .A2(new_n1049), .A3(new_n1244), .A4(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n408), .B1(new_n770), .B2(new_n310), .ZN(new_n1247));
  XOR2_X1   g1047(.A(new_n1247), .B(KEYINPUT117), .Z(new_n1248));
  NOR2_X1   g1048(.A1(new_n1246), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  OR2_X1    g1050(.A1(new_n1250), .A2(KEYINPUT118), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1188), .A2(new_n251), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(new_n1252), .B(KEYINPUT119), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n752), .A2(new_n1001), .B1(new_n746), .B2(new_n403), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n826), .A2(G132), .B1(G128), .B2(new_n781), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n216), .B2(new_n743), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1254), .B(new_n1256), .C1(G150), .C2(new_n757), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1253), .B(new_n1257), .C1(new_n763), .C2(new_n1111), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1250), .A2(KEYINPUT118), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1251), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1241), .B1(new_n1260), .B2(new_n728), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n929), .A2(new_n725), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1263), .B1(new_n1221), .B2(new_n720), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1240), .A2(new_n1265), .ZN(G381));
  AOI21_X1  g1066(.A(new_n1227), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1225), .A2(new_n678), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1214), .B1(new_n1269), .B2(new_n1231), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1159), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1136), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1270), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(new_n1026), .A3(new_n1000), .ZN(new_n1277));
  OR2_X1    g1077(.A1(G393), .A2(G396), .ZN(new_n1278));
  NOR4_X1   g1078(.A1(new_n1277), .A2(G384), .A3(G381), .A4(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1275), .A2(new_n1279), .ZN(new_n1280));
  XOR2_X1   g1080(.A(new_n1280), .B(KEYINPUT120), .Z(G407));
  INV_X1    g1081(.A(G213), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1282), .A2(G343), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1274), .A2(new_n1284), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1285), .B(KEYINPUT121), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(G407), .A2(G213), .A3(new_n1286), .ZN(G409));
  NAND3_X1  g1087(.A1(new_n1186), .A2(new_n1235), .A3(new_n1222), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1288), .A2(new_n1187), .A3(new_n1213), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1283), .B1(new_n1273), .B2(new_n1290), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1291), .B1(new_n1270), .B2(new_n1273), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1283), .A2(G2897), .ZN(new_n1293));
  OAI21_X1  g1093(.A(KEYINPUT60), .B1(new_n1221), .B2(new_n1238), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1234), .A2(new_n1294), .A3(new_n1239), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1296), .A2(KEYINPUT60), .A3(new_n1238), .A4(new_n1142), .ZN(new_n1297));
  AND2_X1   g1097(.A1(new_n1297), .A2(new_n678), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1295), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n1265), .ZN(new_n1300));
  INV_X1    g1100(.A(G384), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1299), .A2(G384), .A3(new_n1265), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1293), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(G384), .B1(new_n1299), .B2(new_n1265), .ZN(new_n1305));
  AOI211_X1 g1105(.A(new_n1301), .B(new_n1264), .C1(new_n1295), .C2(new_n1298), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1293), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(new_n1305), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1304), .A2(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(KEYINPUT61), .B1(new_n1292), .B2(new_n1309), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1284), .B1(G378), .B2(new_n1289), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1311), .B1(G375), .B2(G378), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1313));
  AOI21_X1  g1113(.A(KEYINPUT62), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1314));
  AOI22_X1  g1114(.A1(new_n1153), .A2(new_n1154), .B1(new_n1182), .B2(new_n1185), .ZN(new_n1315));
  OAI21_X1  g1115(.A(KEYINPUT115), .B1(new_n1315), .B2(KEYINPUT57), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n680), .B1(new_n1315), .B2(KEYINPUT57), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1316), .A2(new_n1317), .A3(new_n1231), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1273), .B1(new_n1318), .B2(new_n1215), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT62), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1321));
  NOR4_X1   g1121(.A1(new_n1319), .A2(new_n1320), .A3(new_n1321), .A4(new_n1311), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1310), .B1(new_n1314), .B2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(KEYINPUT126), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(G390), .A2(G387), .ZN(new_n1325));
  XNOR2_X1  g1125(.A(G393), .B(new_n796), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1325), .A2(new_n1277), .A3(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1326), .ZN(new_n1329));
  AOI21_X1  g1129(.A(KEYINPUT123), .B1(new_n1000), .B2(new_n1026), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1329), .B1(new_n1330), .B2(new_n1276), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT123), .ZN(new_n1332));
  AND3_X1   g1132(.A1(G387), .A2(new_n1276), .A3(new_n1332), .ZN(new_n1333));
  OAI21_X1  g1133(.A(KEYINPUT124), .B1(new_n1331), .B2(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(G387), .A2(new_n1332), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1335), .A2(G390), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT124), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1330), .A2(new_n1276), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1336), .A2(new_n1337), .A3(new_n1338), .A4(new_n1329), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1328), .B1(new_n1334), .B2(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT126), .ZN(new_n1341));
  OAI211_X1 g1141(.A(new_n1310), .B(new_n1341), .C1(new_n1314), .C2(new_n1322), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1324), .A2(new_n1340), .A3(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT125), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1334), .A2(new_n1339), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1345), .A2(new_n1327), .ZN(new_n1346));
  NOR3_X1   g1146(.A1(new_n1319), .A2(new_n1321), .A3(new_n1311), .ZN(new_n1347));
  XOR2_X1   g1147(.A(KEYINPUT122), .B(KEYINPUT63), .Z(new_n1348));
  INV_X1    g1148(.A(new_n1348), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1346), .B1(new_n1347), .B2(new_n1349), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(G375), .A2(G378), .ZN(new_n1351));
  NAND4_X1  g1151(.A1(new_n1351), .A2(KEYINPUT63), .A3(new_n1313), .A4(new_n1291), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1313), .A2(new_n1293), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1321), .A2(new_n1307), .ZN(new_n1354));
  OAI211_X1 g1154(.A(new_n1353), .B(new_n1354), .C1(new_n1319), .C2(new_n1311), .ZN(new_n1355));
  INV_X1    g1155(.A(KEYINPUT61), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1352), .A2(new_n1355), .A3(new_n1356), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1344), .B1(new_n1350), .B2(new_n1357), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1359));
  AOI21_X1  g1159(.A(new_n1340), .B1(new_n1359), .B2(new_n1348), .ZN(new_n1360));
  NAND4_X1  g1160(.A1(new_n1360), .A2(KEYINPUT125), .A3(new_n1310), .A4(new_n1352), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1358), .A2(new_n1361), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1343), .A2(new_n1362), .ZN(G405));
  OAI21_X1  g1163(.A(new_n1321), .B1(new_n1275), .B2(new_n1319), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1274), .A2(new_n1351), .A3(new_n1313), .ZN(new_n1365));
  INV_X1    g1165(.A(KEYINPUT127), .ZN(new_n1366));
  AOI22_X1  g1166(.A1(new_n1364), .A2(new_n1365), .B1(new_n1366), .B2(new_n1340), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1346), .A2(KEYINPUT127), .ZN(new_n1368));
  XNOR2_X1  g1168(.A(new_n1367), .B(new_n1368), .ZN(G402));
endmodule


