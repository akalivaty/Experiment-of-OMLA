//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 0 1 1 0 1 0 0 1 0 0 1 0 1 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 0 1 0 1 1 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 0 1 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017;
  NOR2_X1   g000(.A1(G475), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G140), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G125), .ZN(new_n189));
  OR2_X1    g003(.A1(new_n189), .A2(KEYINPUT72), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G140), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n192), .A3(KEYINPUT72), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(KEYINPUT16), .A3(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT16), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n189), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G146), .ZN(new_n198));
  NOR2_X1   g012(.A1(G237), .A2(G953), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G214), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n199), .A2(G143), .A3(G214), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G131), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT17), .ZN(new_n206));
  INV_X1    g020(.A(G131), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n202), .A2(new_n207), .A3(new_n203), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n205), .A2(new_n206), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n194), .A2(new_n210), .A3(new_n196), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n204), .A2(KEYINPUT17), .A3(G131), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n198), .A2(new_n209), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(KEYINPUT18), .A2(G131), .ZN(new_n214));
  XNOR2_X1  g028(.A(new_n204), .B(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n190), .A2(G146), .A3(new_n193), .ZN(new_n216));
  AND2_X1   g030(.A1(new_n189), .A2(new_n192), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(new_n210), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(G113), .B(G122), .ZN(new_n221));
  INV_X1    g035(.A(G104), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n221), .B(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(new_n223), .B(KEYINPUT89), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n213), .A2(new_n220), .A3(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n205), .A2(new_n208), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n217), .A2(KEYINPUT19), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n190), .A2(new_n193), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n228), .B1(new_n229), .B2(KEYINPUT19), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n198), .B(new_n227), .C1(G146), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n223), .B1(new_n231), .B2(new_n220), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n187), .B1(new_n226), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT20), .ZN(new_n234));
  AND2_X1   g048(.A1(new_n231), .A2(new_n220), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n225), .B1(new_n235), .B2(new_n223), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT20), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(new_n237), .A3(new_n187), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n213), .A2(new_n220), .ZN(new_n240));
  INV_X1    g054(.A(new_n223), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(G902), .B1(new_n242), .B2(new_n225), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G475), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n239), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT15), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G478), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT91), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n250), .B1(new_n201), .B2(G128), .ZN(new_n251));
  INV_X1    g065(.A(G128), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(KEYINPUT91), .A3(G143), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n201), .A2(G128), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G134), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n254), .A2(G134), .A3(new_n255), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT13), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n254), .A2(new_n260), .A3(G134), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n258), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n254), .A2(new_n260), .A3(G134), .A4(new_n255), .ZN(new_n263));
  INV_X1    g077(.A(G107), .ZN(new_n264));
  INV_X1    g078(.A(G116), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(G122), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(KEYINPUT66), .B(G116), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT90), .B1(new_n268), .B2(G122), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n265), .A2(KEYINPUT66), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT66), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G116), .ZN(new_n272));
  AND4_X1   g086(.A1(KEYINPUT90), .A2(new_n270), .A3(new_n272), .A4(G122), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n264), .B(new_n267), .C1(new_n269), .C2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n270), .A2(new_n272), .A3(G122), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT90), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n268), .A2(KEYINPUT90), .A3(G122), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n264), .B1(new_n280), .B2(new_n267), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n262), .B(new_n263), .C1(new_n275), .C2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n266), .B1(new_n280), .B2(KEYINPUT14), .ZN(new_n283));
  OR3_X1    g097(.A1(new_n269), .A2(new_n273), .A3(KEYINPUT14), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n264), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n274), .A2(new_n258), .A3(new_n259), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n282), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(KEYINPUT9), .B(G234), .ZN(new_n288));
  INV_X1    g102(.A(G217), .ZN(new_n289));
  NOR3_X1   g103(.A1(new_n288), .A2(new_n289), .A3(G953), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n282), .B(new_n290), .C1(new_n285), .C2(new_n286), .ZN(new_n293));
  AOI21_X1  g107(.A(G902), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT92), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI211_X1 g110(.A(KEYINPUT92), .B(G902), .C1(new_n292), .C2(new_n293), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n249), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  OR2_X1    g112(.A1(new_n297), .A2(new_n249), .ZN(new_n299));
  NOR2_X1   g113(.A1(KEYINPUT93), .A2(G952), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(KEYINPUT93), .A2(G952), .ZN(new_n302));
  AOI21_X1  g116(.A(G953), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(G234), .A2(G237), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT21), .B(G898), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n306), .A2(G902), .A3(G953), .A4(new_n304), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n247), .A2(new_n298), .A3(new_n299), .A4(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(G214), .B1(G237), .B2(G902), .ZN(new_n311));
  XOR2_X1   g125(.A(new_n311), .B(KEYINPUT83), .Z(new_n312));
  NAND3_X1  g126(.A1(new_n270), .A2(new_n272), .A3(G119), .ZN(new_n313));
  INV_X1    g127(.A(G119), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G116), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n313), .A2(KEYINPUT5), .A3(new_n315), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n316), .B(G113), .C1(KEYINPUT5), .C2(new_n315), .ZN(new_n317));
  XOR2_X1   g131(.A(KEYINPUT2), .B(G113), .Z(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(new_n313), .A3(new_n315), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT77), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(new_n264), .A3(G104), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT77), .B1(new_n222), .B2(G107), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n264), .A2(G104), .ZN(new_n324));
  OAI211_X1 g138(.A(G101), .B(new_n322), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT3), .B1(new_n222), .B2(G107), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n327), .A2(new_n264), .A3(G104), .ZN(new_n328));
  INV_X1    g142(.A(G101), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n222), .A2(G107), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n326), .A2(new_n328), .A3(new_n329), .A4(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n325), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT78), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n325), .A2(new_n331), .A3(KEYINPUT78), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OR2_X1    g150(.A1(new_n320), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n326), .A2(new_n328), .A3(new_n330), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G101), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(KEYINPUT4), .A3(new_n331), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT76), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n339), .A2(KEYINPUT76), .A3(KEYINPUT4), .A4(new_n331), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  OR2_X1    g159(.A1(new_n339), .A2(KEYINPUT4), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n313), .A2(new_n315), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT2), .B(G113), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n319), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n337), .B1(new_n345), .B2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(G110), .B(G122), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n337), .B(new_n353), .C1(new_n345), .C2(new_n351), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n355), .A2(KEYINPUT6), .A3(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT6), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n352), .A2(new_n358), .A3(new_n354), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n210), .A2(G143), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n201), .A2(G146), .ZN(new_n361));
  AND2_X1   g175(.A1(KEYINPUT0), .A2(G128), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  XNOR2_X1  g177(.A(G143), .B(G146), .ZN(new_n364));
  XNOR2_X1  g178(.A(KEYINPUT0), .B(G128), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G125), .ZN(new_n367));
  OR2_X1    g181(.A1(new_n367), .A2(KEYINPUT84), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n360), .A2(new_n361), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n360), .A2(KEYINPUT1), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n370), .A3(G128), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n360), .B(new_n361), .C1(KEYINPUT1), .C2(new_n252), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n191), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n367), .A2(KEYINPUT84), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n368), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G224), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n377), .A2(G953), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n376), .B(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n357), .A2(new_n359), .A3(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(KEYINPUT7), .B1(new_n377), .B2(G953), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n374), .A2(KEYINPUT86), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n367), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n374), .A2(KEYINPUT86), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n381), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n385), .B1(new_n376), .B2(new_n381), .ZN(new_n386));
  XNOR2_X1  g200(.A(KEYINPUT85), .B(KEYINPUT8), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n353), .B(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n320), .A2(new_n332), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n388), .B1(new_n337), .B2(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(G902), .B1(new_n391), .B2(new_n356), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n380), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(G210), .B1(G237), .B2(G902), .ZN(new_n394));
  XOR2_X1   g208(.A(new_n394), .B(KEYINPUT87), .Z(new_n395));
  XOR2_X1   g209(.A(new_n395), .B(KEYINPUT88), .Z(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n395), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n380), .A2(new_n392), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n312), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n310), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(G110), .B(G140), .ZN(new_n403));
  INV_X1    g217(.A(G953), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n404), .A2(G227), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n403), .B(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT12), .ZN(new_n407));
  INV_X1    g221(.A(new_n335), .ZN(new_n408));
  AOI21_X1  g222(.A(KEYINPUT78), .B1(new_n325), .B2(new_n331), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n373), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n373), .A2(new_n332), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT64), .ZN(new_n414));
  INV_X1    g228(.A(G137), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AND2_X1   g230(.A1(KEYINPUT11), .A2(G134), .ZN(new_n417));
  NAND2_X1  g231(.A1(KEYINPUT64), .A2(G137), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(KEYINPUT11), .A2(G134), .ZN(new_n420));
  NOR2_X1   g234(.A1(KEYINPUT11), .A2(G134), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n420), .B1(new_n421), .B2(G137), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G131), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n419), .A2(new_n422), .A3(new_n207), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n407), .B1(new_n413), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n411), .B1(new_n336), .B2(new_n373), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n407), .A2(KEYINPUT80), .ZN(new_n429));
  OR2_X1    g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n419), .A2(new_n207), .A3(new_n422), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n207), .B1(new_n419), .B2(new_n422), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT67), .ZN(new_n433));
  NOR3_X1   g247(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(KEYINPUT67), .B1(new_n424), .B2(new_n425), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n436), .B1(new_n428), .B2(KEYINPUT80), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n427), .B1(new_n430), .B2(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n411), .A2(KEYINPUT10), .ZN(new_n439));
  INV_X1    g253(.A(new_n366), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n346), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n439), .B1(new_n441), .B2(new_n344), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n371), .A2(KEYINPUT10), .A3(new_n372), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n334), .A2(new_n443), .A3(new_n335), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT79), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n334), .A2(new_n443), .A3(KEYINPUT79), .A4(new_n335), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n442), .A2(new_n448), .A3(new_n436), .ZN(new_n449));
  AOI21_X1  g263(.A(KEYINPUT81), .B1(new_n438), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n427), .ZN(new_n451));
  INV_X1    g265(.A(new_n436), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n410), .A2(KEYINPUT80), .A3(new_n412), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n452), .B(new_n453), .C1(new_n428), .C2(new_n429), .ZN(new_n454));
  AND4_X1   g268(.A1(KEYINPUT81), .A2(new_n449), .A3(new_n451), .A4(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n406), .B1(new_n450), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n442), .A2(new_n448), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n452), .ZN(new_n458));
  INV_X1    g272(.A(new_n406), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(new_n459), .A3(new_n449), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n456), .A2(G469), .A3(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(G469), .ZN(new_n462));
  INV_X1    g276(.A(G902), .ZN(new_n463));
  INV_X1    g277(.A(new_n449), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n436), .B1(new_n442), .B2(new_n448), .ZN(new_n465));
  OAI211_X1 g279(.A(KEYINPUT82), .B(new_n406), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n438), .A2(new_n459), .A3(new_n449), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n458), .A2(new_n449), .ZN(new_n469));
  AOI21_X1  g283(.A(KEYINPUT82), .B1(new_n469), .B2(new_n406), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n462), .B(new_n463), .C1(new_n468), .C2(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n462), .A2(new_n463), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n461), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(G221), .B1(new_n288), .B2(G902), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT94), .B1(new_n402), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n312), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n380), .A2(new_n392), .A3(new_n399), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n396), .B1(new_n380), .B2(new_n392), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n481), .A2(new_n309), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT94), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n482), .A2(new_n483), .A3(new_n475), .A4(new_n474), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n477), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT71), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n440), .B1(new_n434), .B2(new_n435), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n425), .A2(new_n371), .A3(new_n372), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT65), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n416), .A2(new_n257), .A3(new_n418), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n207), .B1(G134), .B2(G137), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n491), .A2(new_n490), .A3(new_n492), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n350), .B1(new_n489), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n487), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n199), .A2(G210), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n499), .B(KEYINPUT27), .ZN(new_n500));
  XNOR2_X1  g314(.A(KEYINPUT26), .B(G101), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n500), .B(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  AOI22_X1  g318(.A1(new_n489), .A2(new_n496), .B1(new_n426), .B2(new_n440), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n433), .B1(new_n431), .B2(new_n432), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n424), .A2(KEYINPUT67), .A3(new_n425), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n366), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n491), .A2(new_n490), .A3(new_n492), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n509), .A2(new_n493), .ZN(new_n510));
  OAI21_X1  g324(.A(KEYINPUT30), .B1(new_n510), .B2(new_n488), .ZN(new_n511));
  OAI22_X1  g325(.A1(new_n505), .A2(KEYINPUT30), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT68), .ZN(new_n513));
  INV_X1    g327(.A(new_n319), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n318), .B1(new_n315), .B2(new_n313), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n512), .A2(new_n513), .A3(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT30), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n518), .B1(new_n489), .B2(new_n496), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n440), .B1(new_n431), .B2(new_n432), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n520), .B1(new_n510), .B2(new_n488), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n487), .A2(new_n519), .B1(new_n521), .B2(new_n518), .ZN(new_n522));
  AOI21_X1  g336(.A(KEYINPUT68), .B1(new_n522), .B2(new_n350), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n504), .B1(new_n517), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT31), .ZN(new_n525));
  AOI21_X1  g339(.A(KEYINPUT28), .B1(new_n487), .B2(new_n497), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n516), .B1(new_n510), .B2(new_n488), .ZN(new_n527));
  OAI22_X1  g341(.A1(new_n516), .A2(new_n505), .B1(new_n508), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n526), .B1(new_n528), .B2(KEYINPUT28), .ZN(new_n529));
  OAI21_X1  g343(.A(KEYINPUT69), .B1(new_n529), .B2(new_n502), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT28), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n531), .B1(new_n508), .B2(new_n527), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n487), .A2(new_n497), .B1(new_n521), .B2(new_n350), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n532), .B1(new_n533), .B2(new_n531), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT69), .ZN(new_n535));
  INV_X1    g349(.A(new_n502), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n530), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n513), .B1(new_n512), .B2(new_n516), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n522), .A2(KEYINPUT68), .A3(new_n350), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n503), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT31), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n525), .A2(new_n538), .A3(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT32), .ZN(new_n545));
  NOR2_X1   g359(.A1(G472), .A2(G902), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n545), .B1(new_n544), .B2(new_n546), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(G472), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n498), .B1(new_n517), .B2(new_n523), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT70), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n552), .A3(new_n536), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n508), .A2(new_n527), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n554), .B1(new_n539), .B2(new_n540), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT70), .B1(new_n555), .B2(new_n502), .ZN(new_n556));
  AOI21_X1  g370(.A(KEYINPUT29), .B1(new_n529), .B2(new_n502), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n553), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n489), .A2(new_n496), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n350), .B1(new_n560), .B2(new_n508), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n531), .B1(new_n561), .B2(new_n498), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n562), .A2(new_n526), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n502), .A2(KEYINPUT29), .ZN(new_n564));
  AOI21_X1  g378(.A(G902), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n550), .B1(new_n558), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n486), .B1(new_n549), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n404), .A2(G221), .A3(G234), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(KEYINPUT74), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT22), .B(G137), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n569), .B(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n198), .A2(new_n211), .ZN(new_n572));
  XOR2_X1   g386(.A(G119), .B(G128), .Z(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT24), .B(G110), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT23), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n576), .B1(new_n314), .B2(G128), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n252), .A2(KEYINPUT23), .A3(G119), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n577), .B(new_n578), .C1(G119), .C2(new_n252), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n575), .B1(G110), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n572), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT73), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n572), .A2(KEYINPUT73), .A3(new_n580), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n573), .A2(new_n574), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n586), .B1(new_n579), .B2(G110), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n198), .A2(new_n218), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n571), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n588), .ZN(new_n590));
  INV_X1    g404(.A(new_n571), .ZN(new_n591));
  AOI211_X1 g405(.A(new_n590), .B(new_n591), .C1(new_n583), .C2(new_n584), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n593), .A2(KEYINPUT25), .A3(new_n463), .ZN(new_n594));
  INV_X1    g408(.A(new_n584), .ZN(new_n595));
  AOI21_X1  g409(.A(KEYINPUT73), .B1(new_n572), .B2(new_n580), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n588), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n591), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n585), .A2(new_n588), .A3(new_n571), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n598), .A2(new_n463), .A3(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT25), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n594), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n289), .B1(G234), .B2(new_n463), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n604), .A2(G902), .ZN(new_n605));
  OAI21_X1  g419(.A(KEYINPUT75), .B1(new_n589), .B2(new_n592), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT75), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n598), .A2(new_n607), .A3(new_n599), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  AOI22_X1  g423(.A1(new_n603), .A2(new_n604), .B1(new_n605), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n516), .B1(new_n559), .B2(new_n520), .ZN(new_n611));
  OAI21_X1  g425(.A(KEYINPUT28), .B1(new_n554), .B2(new_n611), .ZN(new_n612));
  AOI211_X1 g426(.A(KEYINPUT69), .B(new_n502), .C1(new_n612), .C2(new_n532), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n535), .B1(new_n534), .B2(new_n536), .ZN(new_n614));
  OAI22_X1  g428(.A1(new_n613), .A2(new_n614), .B1(new_n541), .B2(new_n542), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n524), .A2(KEYINPUT31), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n546), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(KEYINPUT32), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n566), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n620), .A2(KEYINPUT71), .A3(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n567), .A2(new_n610), .A3(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n485), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(new_n329), .ZN(G3));
  NAND2_X1  g439(.A1(new_n544), .A2(new_n463), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(G472), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n617), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n476), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n629), .A2(new_n630), .A3(new_n610), .ZN(new_n631));
  INV_X1    g445(.A(new_n311), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n393), .A2(new_n395), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n632), .B1(new_n633), .B2(new_n400), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n292), .A2(new_n293), .ZN(new_n635));
  OR2_X1    g449(.A1(new_n635), .A2(KEYINPUT33), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(KEYINPUT33), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n636), .A2(G478), .A3(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(G478), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n463), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n640), .B1(new_n294), .B2(new_n639), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n642), .A2(new_n247), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n634), .A2(new_n643), .A3(new_n308), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n631), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(KEYINPUT34), .B(G104), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G6));
  NAND2_X1  g461(.A1(new_n298), .A2(new_n299), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n308), .B(KEYINPUT96), .Z(new_n649));
  NAND3_X1  g463(.A1(new_n634), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n244), .A2(KEYINPUT95), .A3(G475), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT95), .ZN(new_n652));
  INV_X1    g466(.A(G475), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n652), .B1(new_n243), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n239), .A2(new_n651), .A3(new_n654), .ZN(new_n655));
  OR2_X1    g469(.A1(new_n650), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n631), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT35), .B(G107), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G9));
  INV_X1    g473(.A(KEYINPUT97), .ZN(new_n660));
  AOI21_X1  g474(.A(KEYINPUT25), .B1(new_n593), .B2(new_n463), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n600), .A2(new_n601), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n604), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n591), .A2(KEYINPUT36), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n597), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n605), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n660), .B1(new_n628), .B2(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n627), .A2(new_n667), .A3(KEYINPUT97), .A4(new_n617), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n477), .A2(new_n669), .A3(new_n484), .A4(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT37), .B(G110), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G12));
  INV_X1    g487(.A(KEYINPUT98), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n298), .A2(new_n299), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n304), .A2(G902), .A3(G953), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n305), .B1(G900), .B2(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n239), .A2(new_n651), .A3(new_n654), .A4(new_n677), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n674), .B1(new_n675), .B2(new_n678), .ZN(new_n679));
  AND4_X1   g493(.A1(new_n239), .A2(new_n651), .A3(new_n654), .A4(new_n677), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n648), .A2(new_n680), .A3(KEYINPUT98), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n679), .A2(new_n634), .A3(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n476), .A2(new_n668), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n682), .A2(new_n567), .A3(new_n622), .A4(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G128), .ZN(G30));
  NOR2_X1   g499(.A1(new_n555), .A2(new_n536), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n561), .A2(new_n498), .A3(new_n536), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n463), .ZN(new_n688));
  OAI21_X1  g502(.A(G472), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n620), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g504(.A(new_n690), .B(KEYINPUT99), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n677), .B(KEYINPUT39), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n630), .A2(new_n692), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n693), .A2(KEYINPUT40), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n693), .A2(KEYINPUT40), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n479), .A2(new_n480), .ZN(new_n696));
  XOR2_X1   g510(.A(new_n696), .B(KEYINPUT38), .Z(new_n697));
  NOR3_X1   g511(.A1(new_n675), .A2(new_n247), .A3(new_n632), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n697), .A2(new_n668), .A3(new_n698), .ZN(new_n699));
  NOR4_X1   g513(.A1(new_n691), .A2(new_n694), .A3(new_n695), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(new_n201), .ZN(G45));
  NAND4_X1  g515(.A1(new_n638), .A2(new_n246), .A3(new_n641), .A4(new_n677), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT100), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n634), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n399), .B1(new_n380), .B2(new_n392), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n311), .B1(new_n479), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g521(.A(KEYINPUT100), .B1(new_n707), .B2(new_n702), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n567), .A2(new_n709), .A3(new_n622), .A4(new_n683), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G146), .ZN(G48));
  INV_X1    g525(.A(new_n475), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n463), .B1(new_n468), .B2(new_n470), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(G469), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(KEYINPUT101), .A3(new_n471), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT101), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n713), .A2(new_n716), .A3(G469), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n712), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n567), .A2(new_n610), .A3(new_n622), .A4(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT102), .ZN(new_n721));
  INV_X1    g535(.A(new_n644), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g537(.A(KEYINPUT102), .B1(new_n719), .B2(new_n644), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(KEYINPUT41), .B(G113), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(G15));
  NOR2_X1   g541(.A1(new_n719), .A2(new_n656), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(new_n265), .ZN(G18));
  NAND4_X1  g543(.A1(new_n567), .A2(new_n622), .A3(new_n310), .A4(new_n667), .ZN(new_n730));
  AOI211_X1 g544(.A(new_n712), .B(new_n707), .C1(new_n715), .C2(new_n717), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(new_n314), .ZN(G21));
  NOR2_X1   g548(.A1(new_n650), .A2(new_n247), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n536), .B1(new_n562), .B2(new_n526), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n736), .B1(new_n541), .B2(new_n542), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(KEYINPUT103), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT103), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n739), .B(new_n736), .C1(new_n541), .C2(new_n542), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n738), .A2(new_n543), .A3(new_n740), .ZN(new_n741));
  AOI22_X1  g555(.A1(new_n546), .A2(new_n741), .B1(new_n626), .B2(G472), .ZN(new_n742));
  AOI21_X1  g556(.A(KEYINPUT104), .B1(new_n742), .B2(new_n610), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n739), .B1(new_n525), .B2(new_n736), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n740), .A2(new_n543), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n546), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  AND4_X1   g560(.A1(KEYINPUT104), .A2(new_n627), .A3(new_n746), .A4(new_n610), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n718), .B(new_n735), .C1(new_n743), .C2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G122), .ZN(G24));
  INV_X1    g563(.A(KEYINPUT105), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n750), .B1(new_n742), .B2(new_n667), .ZN(new_n751));
  AND4_X1   g565(.A1(new_n750), .A2(new_n627), .A3(new_n667), .A4(new_n746), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n731), .B(new_n703), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G125), .ZN(G27));
  INV_X1    g568(.A(KEYINPUT108), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT42), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n696), .A2(new_n475), .A3(new_n311), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT106), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n456), .A2(new_n758), .A3(G469), .A4(new_n460), .ZN(new_n759));
  AND3_X1   g573(.A1(new_n759), .A2(new_n471), .A3(new_n473), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n461), .A2(KEYINPUT106), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n757), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n567), .A2(new_n762), .A3(new_n610), .A4(new_n622), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n756), .B1(new_n763), .B2(new_n702), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT107), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OAI211_X1 g580(.A(KEYINPUT107), .B(new_n756), .C1(new_n763), .C2(new_n702), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n762), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n620), .A2(new_n621), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n610), .ZN(new_n771));
  NOR4_X1   g585(.A1(new_n769), .A2(new_n771), .A3(new_n756), .A4(new_n702), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n755), .B1(new_n768), .B2(new_n773), .ZN(new_n774));
  AOI211_X1 g588(.A(KEYINPUT108), .B(new_n772), .C1(new_n766), .C2(new_n767), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G131), .ZN(G33));
  NAND2_X1  g591(.A1(new_n679), .A2(new_n681), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n763), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G134), .ZN(G36));
  AND2_X1   g594(.A1(new_n456), .A2(new_n460), .ZN(new_n781));
  OAI21_X1  g595(.A(G469), .B1(new_n781), .B2(KEYINPUT45), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n782), .A2(KEYINPUT109), .ZN(new_n783));
  AOI22_X1  g597(.A1(new_n782), .A2(KEYINPUT109), .B1(KEYINPUT45), .B2(new_n781), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n472), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n785), .A2(KEYINPUT46), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n471), .B1(new_n785), .B2(KEYINPUT46), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AND2_X1   g602(.A1(KEYINPUT110), .A2(KEYINPUT43), .ZN(new_n789));
  NOR2_X1   g603(.A1(KEYINPUT110), .A2(KEYINPUT43), .ZN(new_n790));
  OAI22_X1  g604(.A1(new_n642), .A2(new_n246), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n642), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n247), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n791), .B1(new_n793), .B2(new_n790), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n794), .A2(new_n628), .A3(new_n667), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT44), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n479), .A2(new_n480), .A3(new_n632), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n797), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n788), .A2(new_n475), .A3(new_n692), .A4(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G137), .ZN(G39));
  AND3_X1   g617(.A1(new_n620), .A2(KEYINPUT71), .A3(new_n621), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT71), .B1(new_n620), .B2(new_n621), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n610), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n807), .A2(new_n703), .A3(new_n799), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n788), .A2(KEYINPUT47), .A3(new_n475), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n475), .B1(new_n786), .B2(new_n787), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT47), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI211_X1 g626(.A(new_n806), .B(new_n808), .C1(new_n809), .C2(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(new_n188), .ZN(G42));
  AND2_X1   g628(.A1(new_n715), .A2(new_n717), .ZN(new_n815));
  XOR2_X1   g629(.A(new_n815), .B(KEYINPUT49), .Z(new_n816));
  NAND2_X1  g630(.A1(new_n478), .A2(new_n475), .ZN(new_n817));
  NOR4_X1   g631(.A1(new_n697), .A2(new_n807), .A3(new_n793), .A4(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n816), .A2(new_n691), .A3(new_n818), .ZN(new_n819));
  XOR2_X1   g633(.A(new_n819), .B(KEYINPUT111), .Z(new_n820));
  OAI211_X1 g634(.A(new_n809), .B(new_n812), .C1(new_n475), .C2(new_n815), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n743), .A2(new_n747), .ZN(new_n822));
  INV_X1    g636(.A(new_n305), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n822), .A2(new_n823), .A3(new_n794), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n821), .A2(new_n799), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n697), .A2(new_n311), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n825), .A2(new_n718), .A3(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n751), .A2(new_n752), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n815), .A2(new_n305), .A3(new_n757), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(new_n794), .ZN(new_n831));
  OAI22_X1  g645(.A1(new_n828), .A2(KEYINPUT50), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n832), .B1(KEYINPUT50), .B2(new_n828), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n691), .A2(new_n830), .A3(new_n610), .ZN(new_n834));
  OR2_X1    g648(.A1(new_n834), .A2(KEYINPUT119), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(KEYINPUT119), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n792), .A2(new_n246), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n838), .A2(KEYINPUT120), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT120), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n834), .B(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n840), .B1(new_n842), .B2(new_n837), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n826), .B(new_n833), .C1(new_n839), .C2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT118), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT51), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT51), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n844), .A2(new_n845), .A3(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n303), .B1(new_n824), .B2(new_n732), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n831), .A2(new_n771), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT48), .ZN(new_n852));
  AOI211_X1 g666(.A(new_n850), .B(new_n852), .C1(new_n643), .C2(new_n842), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n847), .A2(new_n849), .A3(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n748), .B1(new_n719), .B2(new_n656), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n855), .A2(new_n733), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n643), .B1(new_n648), .B2(new_n247), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n401), .A2(new_n649), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n859), .A2(new_n610), .A3(new_n630), .A4(new_n629), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n671), .B(new_n860), .C1(new_n623), .C2(new_n485), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n703), .B(new_n762), .C1(new_n751), .C2(new_n752), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT112), .B1(new_n648), .B2(new_n678), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT112), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n680), .A2(new_n865), .A3(new_n298), .A4(new_n299), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n864), .A2(new_n866), .A3(new_n799), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n867), .A2(new_n476), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n868), .A2(new_n567), .A3(new_n622), .A4(new_n667), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n863), .B(new_n869), .C1(new_n763), .C2(new_n778), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n725), .A2(new_n856), .A3(new_n862), .A4(new_n871), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n774), .A2(new_n775), .A3(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT53), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n684), .A2(new_n710), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT115), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n633), .A2(new_n400), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n698), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n677), .A2(KEYINPUT113), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n677), .A2(KEYINPUT113), .ZN(new_n880));
  NOR4_X1   g694(.A1(new_n667), .A2(new_n712), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n760), .A2(new_n761), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n878), .A2(new_n881), .A3(new_n690), .A4(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n875), .A2(new_n876), .A3(new_n753), .A4(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n753), .A2(new_n684), .A3(new_n710), .A4(new_n883), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT115), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT52), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n884), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  OR3_X1    g702(.A1(new_n885), .A2(KEYINPUT114), .A3(new_n887), .ZN(new_n889));
  OAI21_X1  g703(.A(KEYINPUT114), .B1(new_n885), .B2(new_n887), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n873), .A2(new_n874), .A3(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n806), .A2(new_n610), .A3(new_n703), .A4(new_n762), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT107), .B1(new_n893), .B2(new_n756), .ZN(new_n894));
  INV_X1    g708(.A(new_n767), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n773), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(KEYINPUT108), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n768), .A2(new_n755), .A3(new_n773), .ZN(new_n898));
  AND4_X1   g712(.A1(new_n725), .A2(new_n856), .A3(new_n862), .A4(new_n871), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n884), .A2(new_n886), .A3(new_n887), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n887), .B1(new_n884), .B2(new_n886), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(KEYINPUT53), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n892), .A2(new_n904), .A3(KEYINPUT54), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n874), .B1(new_n900), .B2(new_n903), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT54), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n861), .A2(new_n870), .A3(new_n874), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n896), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT116), .B1(new_n725), .B2(new_n856), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n725), .A2(new_n856), .A3(KEYINPUT116), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n909), .B(new_n891), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n906), .A2(new_n907), .A3(new_n912), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n905), .A2(new_n913), .A3(KEYINPUT117), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT117), .B1(new_n905), .B2(new_n913), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n854), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(G952), .A2(G953), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n820), .B1(new_n916), .B2(new_n917), .ZN(G75));
  OR2_X1    g732(.A1(new_n901), .A2(new_n902), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT53), .B1(new_n873), .B2(new_n919), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n896), .B(new_n908), .C1(new_n911), .C2(new_n910), .ZN(new_n921));
  INV_X1    g735(.A(new_n891), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(G902), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(KEYINPUT56), .B1(new_n925), .B2(new_n395), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n357), .A2(new_n359), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(new_n379), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT55), .Z(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n404), .A2(G952), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n924), .A2(new_n396), .ZN(new_n934));
  AOI21_X1  g748(.A(KEYINPUT56), .B1(new_n930), .B2(KEYINPUT121), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n935), .B1(KEYINPUT121), .B2(new_n930), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n933), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n931), .A2(new_n937), .ZN(G51));
  INV_X1    g752(.A(KEYINPUT123), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n783), .A2(new_n784), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT122), .Z(new_n941));
  AOI211_X1 g755(.A(new_n463), .B(new_n941), .C1(new_n906), .C2(new_n912), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n472), .B(KEYINPUT57), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n906), .A2(new_n907), .A3(new_n912), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n907), .B1(new_n906), .B2(new_n912), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n468), .A2(new_n470), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n942), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n939), .B1(new_n949), .B2(new_n932), .ZN(new_n950));
  OAI21_X1  g764(.A(KEYINPUT54), .B1(new_n920), .B2(new_n923), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n913), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n947), .B1(new_n952), .B2(new_n943), .ZN(new_n953));
  OAI211_X1 g767(.A(KEYINPUT123), .B(new_n933), .C1(new_n953), .C2(new_n942), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n950), .A2(new_n954), .ZN(G54));
  NAND2_X1  g769(.A1(KEYINPUT58), .A2(G475), .ZN(new_n956));
  OAI221_X1 g770(.A(new_n225), .B1(new_n223), .B2(new_n235), .C1(new_n924), .C2(new_n956), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n925), .A2(KEYINPUT58), .A3(G475), .A4(new_n236), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n957), .A2(new_n958), .A3(new_n933), .ZN(G60));
  NAND2_X1  g773(.A1(new_n636), .A2(new_n637), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n640), .B(KEYINPUT59), .ZN(new_n962));
  AOI211_X1 g776(.A(new_n961), .B(new_n962), .C1(new_n951), .C2(new_n913), .ZN(new_n963));
  INV_X1    g777(.A(new_n962), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n964), .B1(new_n914), .B2(new_n915), .ZN(new_n965));
  AOI211_X1 g779(.A(new_n932), .B(new_n963), .C1(new_n965), .C2(new_n961), .ZN(G63));
  NAND2_X1  g780(.A1(G217), .A2(G902), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT60), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n968), .B1(new_n906), .B2(new_n912), .ZN(new_n969));
  OR2_X1    g783(.A1(new_n969), .A2(new_n609), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n665), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n970), .A2(new_n933), .A3(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT61), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n972), .B(new_n973), .ZN(G66));
  OAI21_X1  g788(.A(G953), .B1(new_n306), .B2(new_n377), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n725), .A2(new_n856), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n976), .A2(new_n861), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n975), .B1(new_n977), .B2(G953), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n927), .B1(G898), .B2(new_n404), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT124), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n978), .B(new_n980), .ZN(G69));
  AOI21_X1  g795(.A(new_n404), .B1(G227), .B2(G900), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n982), .A2(KEYINPUT127), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n875), .A2(new_n753), .ZN(new_n984));
  OR3_X1    g798(.A1(new_n700), .A2(new_n984), .A3(KEYINPUT62), .ZN(new_n985));
  OAI21_X1  g799(.A(KEYINPUT62), .B1(new_n700), .B2(new_n984), .ZN(new_n986));
  NOR4_X1   g800(.A1(new_n623), .A2(new_n693), .A3(new_n800), .A4(new_n857), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT125), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n985), .A2(new_n802), .A3(new_n986), .A4(new_n988), .ZN(new_n989));
  OR3_X1    g803(.A1(new_n989), .A2(new_n813), .A3(KEYINPUT126), .ZN(new_n990));
  OAI21_X1  g804(.A(KEYINPUT126), .B1(new_n989), .B2(new_n813), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n522), .B(new_n230), .ZN(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n994), .A2(G953), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n983), .B1(new_n992), .B2(new_n995), .ZN(new_n996));
  AND3_X1   g810(.A1(new_n878), .A2(new_n610), .A3(new_n770), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n788), .A2(new_n475), .A3(new_n692), .A4(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(new_n984), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n802), .A2(new_n998), .A3(new_n779), .A4(new_n999), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n813), .A2(new_n1000), .ZN(new_n1001));
  AND3_X1   g815(.A1(new_n1001), .A2(new_n404), .A3(new_n776), .ZN(new_n1002));
  AND2_X1   g816(.A1(G900), .A2(G953), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n994), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n996), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n982), .A2(KEYINPUT127), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1005), .B(new_n1006), .ZN(G72));
  NAND2_X1  g821(.A1(new_n892), .A2(new_n904), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n553), .A2(new_n556), .A3(new_n524), .ZN(new_n1009));
  NAND2_X1  g823(.A1(G472), .A2(G902), .ZN(new_n1010));
  XOR2_X1   g824(.A(new_n1010), .B(KEYINPUT63), .Z(new_n1011));
  NAND2_X1  g825(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n933), .B1(new_n1008), .B2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1001), .A2(new_n776), .A3(new_n977), .ZN(new_n1014));
  AOI211_X1 g828(.A(new_n551), .B(new_n502), .C1(new_n1014), .C2(new_n1011), .ZN(new_n1015));
  INV_X1    g829(.A(new_n977), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1011), .B1(new_n992), .B2(new_n1016), .ZN(new_n1017));
  AOI211_X1 g831(.A(new_n1013), .B(new_n1015), .C1(new_n686), .C2(new_n1017), .ZN(G57));
endmodule


