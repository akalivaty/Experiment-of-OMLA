

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580;

  AND2_X1 U320 ( .A1(n496), .A2(n454), .ZN(n288) );
  AND2_X1 U321 ( .A1(n496), .A2(n454), .ZN(n559) );
  NOR2_X1 U322 ( .A1(n394), .A2(n393), .ZN(n396) );
  XNOR2_X1 U323 ( .A(n326), .B(n325), .ZN(n329) );
  AND2_X1 U324 ( .A1(G231GAT), .A2(G233GAT), .ZN(n289) );
  XOR2_X1 U325 ( .A(G1GAT), .B(KEYINPUT72), .Z(n290) );
  XNOR2_X1 U326 ( .A(n447), .B(n289), .ZN(n309) );
  XNOR2_X1 U327 ( .A(n354), .B(n309), .ZN(n316) );
  XNOR2_X1 U328 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U329 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U330 ( .A(n458), .B(n457), .ZN(G1349GAT) );
  XOR2_X1 U331 ( .A(G71GAT), .B(G190GAT), .Z(n292) );
  XNOR2_X1 U332 ( .A(G43GAT), .B(G99GAT), .ZN(n291) );
  XNOR2_X1 U333 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U334 ( .A(G176GAT), .B(n293), .Z(n295) );
  NAND2_X1 U335 ( .A1(G227GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U336 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U337 ( .A(KEYINPUT20), .B(KEYINPUT90), .Z(n297) );
  XNOR2_X1 U338 ( .A(G15GAT), .B(KEYINPUT66), .ZN(n296) );
  XNOR2_X1 U339 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U340 ( .A(n299), .B(n298), .Z(n307) );
  XOR2_X1 U341 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n301) );
  XNOR2_X1 U342 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n300) );
  XNOR2_X1 U343 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U344 ( .A(G169GAT), .B(n302), .Z(n412) );
  XOR2_X1 U345 ( .A(G127GAT), .B(G134GAT), .Z(n304) );
  XNOR2_X1 U346 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n303) );
  XNOR2_X1 U347 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U348 ( .A(G113GAT), .B(n305), .Z(n432) );
  XNOR2_X1 U349 ( .A(n412), .B(n432), .ZN(n306) );
  XNOR2_X1 U350 ( .A(n307), .B(n306), .ZN(n524) );
  INV_X1 U351 ( .A(n524), .ZN(n496) );
  XOR2_X1 U352 ( .A(KEYINPUT115), .B(KEYINPUT47), .Z(n385) );
  XNOR2_X1 U353 ( .A(G15GAT), .B(KEYINPUT73), .ZN(n308) );
  XNOR2_X1 U354 ( .A(n290), .B(n308), .ZN(n354) );
  XOR2_X1 U355 ( .A(G22GAT), .B(G155GAT), .Z(n447) );
  XOR2_X1 U356 ( .A(KEYINPUT85), .B(G64GAT), .Z(n311) );
  XNOR2_X1 U357 ( .A(G211GAT), .B(G78GAT), .ZN(n310) );
  XNOR2_X1 U358 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U359 ( .A(G8GAT), .B(KEYINPUT80), .Z(n397) );
  XOR2_X1 U360 ( .A(n312), .B(n397), .Z(n314) );
  XNOR2_X1 U361 ( .A(G183GAT), .B(G127GAT), .ZN(n313) );
  XNOR2_X1 U362 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U363 ( .A(n316), .B(n315), .ZN(n326) );
  XOR2_X1 U364 ( .A(KEYINPUT15), .B(KEYINPUT86), .Z(n318) );
  XNOR2_X1 U365 ( .A(KEYINPUT88), .B(KEYINPUT84), .ZN(n317) );
  XNOR2_X1 U366 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U367 ( .A(KEYINPUT12), .B(KEYINPUT81), .Z(n320) );
  XNOR2_X1 U368 ( .A(KEYINPUT87), .B(KEYINPUT82), .ZN(n319) );
  XNOR2_X1 U369 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U370 ( .A(n322), .B(n321), .Z(n324) );
  INV_X1 U371 ( .A(KEYINPUT83), .ZN(n323) );
  XNOR2_X1 U372 ( .A(G71GAT), .B(G57GAT), .ZN(n327) );
  XNOR2_X1 U373 ( .A(n327), .B(KEYINPUT13), .ZN(n337) );
  XNOR2_X1 U374 ( .A(n337), .B(KEYINPUT14), .ZN(n328) );
  XNOR2_X1 U375 ( .A(n329), .B(n328), .ZN(n556) );
  INV_X1 U376 ( .A(KEYINPUT77), .ZN(n333) );
  XOR2_X1 U377 ( .A(KEYINPUT76), .B(G85GAT), .Z(n331) );
  XNOR2_X1 U378 ( .A(G99GAT), .B(G92GAT), .ZN(n330) );
  XNOR2_X1 U379 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U380 ( .A(n333), .B(n332), .ZN(n373) );
  XOR2_X1 U381 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n335) );
  XNOR2_X1 U382 ( .A(G120GAT), .B(KEYINPUT33), .ZN(n334) );
  XNOR2_X1 U383 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U384 ( .A(n373), .B(n336), .Z(n346) );
  XOR2_X1 U385 ( .A(G176GAT), .B(G64GAT), .Z(n398) );
  XOR2_X1 U386 ( .A(n337), .B(n398), .Z(n339) );
  NAND2_X1 U387 ( .A1(G230GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U388 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U389 ( .A(n340), .B(KEYINPUT78), .Z(n344) );
  XOR2_X1 U390 ( .A(G78GAT), .B(G148GAT), .Z(n342) );
  XNOR2_X1 U391 ( .A(G106GAT), .B(G204GAT), .ZN(n341) );
  XNOR2_X1 U392 ( .A(n342), .B(n341), .ZN(n439) );
  XNOR2_X1 U393 ( .A(n439), .B(KEYINPUT75), .ZN(n343) );
  XNOR2_X1 U394 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U395 ( .A(n346), .B(n345), .ZN(n570) );
  XOR2_X1 U396 ( .A(n570), .B(KEYINPUT41), .Z(n347) );
  XNOR2_X1 U397 ( .A(n347), .B(KEYINPUT65), .ZN(n544) );
  XOR2_X1 U398 ( .A(KEYINPUT29), .B(KEYINPUT69), .Z(n349) );
  XNOR2_X1 U399 ( .A(G141GAT), .B(G8GAT), .ZN(n348) );
  XNOR2_X1 U400 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U401 ( .A(G22GAT), .B(G197GAT), .Z(n351) );
  XNOR2_X1 U402 ( .A(G169GAT), .B(G113GAT), .ZN(n350) );
  XNOR2_X1 U403 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U404 ( .A(n353), .B(n352), .ZN(n367) );
  XOR2_X1 U405 ( .A(G50GAT), .B(n354), .Z(n356) );
  NAND2_X1 U406 ( .A1(G229GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U407 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U408 ( .A(n357), .B(G36GAT), .Z(n365) );
  XOR2_X1 U409 ( .A(KEYINPUT71), .B(KEYINPUT7), .Z(n359) );
  XNOR2_X1 U410 ( .A(G43GAT), .B(G29GAT), .ZN(n358) );
  XNOR2_X1 U411 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U412 ( .A(KEYINPUT8), .B(n360), .Z(n380) );
  XOR2_X1 U413 ( .A(KEYINPUT70), .B(KEYINPUT74), .Z(n362) );
  XNOR2_X1 U414 ( .A(KEYINPUT30), .B(KEYINPUT68), .ZN(n361) );
  XNOR2_X1 U415 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U416 ( .A(n380), .B(n363), .ZN(n364) );
  XNOR2_X1 U417 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U418 ( .A(n367), .B(n366), .ZN(n554) );
  INV_X1 U419 ( .A(n554), .ZN(n567) );
  NOR2_X1 U420 ( .A1(n544), .A2(n567), .ZN(n368) );
  XNOR2_X1 U421 ( .A(n368), .B(KEYINPUT46), .ZN(n369) );
  NOR2_X1 U422 ( .A1(n556), .A2(n369), .ZN(n383) );
  XOR2_X1 U423 ( .A(KEYINPUT79), .B(KEYINPUT11), .Z(n371) );
  XOR2_X1 U424 ( .A(G50GAT), .B(G162GAT), .Z(n448) );
  XOR2_X1 U425 ( .A(G36GAT), .B(G190GAT), .Z(n408) );
  XNOR2_X1 U426 ( .A(n448), .B(n408), .ZN(n370) );
  XNOR2_X1 U427 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U428 ( .A(KEYINPUT10), .B(n372), .Z(n375) );
  XNOR2_X1 U429 ( .A(G218GAT), .B(n373), .ZN(n374) );
  XNOR2_X1 U430 ( .A(n375), .B(n374), .ZN(n379) );
  XOR2_X1 U431 ( .A(KEYINPUT9), .B(G106GAT), .Z(n377) );
  NAND2_X1 U432 ( .A1(G232GAT), .A2(G233GAT), .ZN(n376) );
  XOR2_X1 U433 ( .A(n377), .B(n376), .Z(n378) );
  XNOR2_X1 U434 ( .A(n379), .B(n378), .ZN(n382) );
  XNOR2_X1 U435 ( .A(n380), .B(G134GAT), .ZN(n381) );
  XNOR2_X1 U436 ( .A(n382), .B(n381), .ZN(n552) );
  NAND2_X1 U437 ( .A1(n383), .A2(n552), .ZN(n384) );
  XNOR2_X1 U438 ( .A(n385), .B(n384), .ZN(n394) );
  XOR2_X1 U439 ( .A(KEYINPUT36), .B(KEYINPUT108), .Z(n386) );
  XNOR2_X1 U440 ( .A(n552), .B(n386), .ZN(n576) );
  NAND2_X1 U441 ( .A1(n576), .A2(n556), .ZN(n387) );
  XNOR2_X1 U442 ( .A(n387), .B(KEYINPUT45), .ZN(n388) );
  XNOR2_X1 U443 ( .A(KEYINPUT67), .B(n388), .ZN(n389) );
  INV_X1 U444 ( .A(n389), .ZN(n390) );
  NOR2_X1 U445 ( .A1(n570), .A2(n390), .ZN(n391) );
  XOR2_X1 U446 ( .A(n391), .B(KEYINPUT116), .Z(n392) );
  NOR2_X1 U447 ( .A1(n554), .A2(n392), .ZN(n393) );
  XNOR2_X1 U448 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n395) );
  XNOR2_X1 U449 ( .A(n396), .B(n395), .ZN(n540) );
  XOR2_X1 U450 ( .A(n398), .B(n397), .Z(n400) );
  NAND2_X1 U451 ( .A1(G226GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U452 ( .A(n400), .B(n399), .ZN(n404) );
  XOR2_X1 U453 ( .A(KEYINPUT102), .B(KEYINPUT101), .Z(n402) );
  XNOR2_X1 U454 ( .A(G204GAT), .B(G92GAT), .ZN(n401) );
  XNOR2_X1 U455 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U456 ( .A(n404), .B(n403), .Z(n410) );
  XOR2_X1 U457 ( .A(KEYINPUT21), .B(G218GAT), .Z(n406) );
  XNOR2_X1 U458 ( .A(KEYINPUT94), .B(G211GAT), .ZN(n405) );
  XNOR2_X1 U459 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U460 ( .A(G197GAT), .B(n407), .Z(n452) );
  XNOR2_X1 U461 ( .A(n452), .B(n408), .ZN(n409) );
  XNOR2_X1 U462 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U463 ( .A(n412), .B(n411), .ZN(n517) );
  NOR2_X1 U464 ( .A1(n540), .A2(n517), .ZN(n414) );
  XNOR2_X1 U465 ( .A(KEYINPUT123), .B(KEYINPUT54), .ZN(n413) );
  XNOR2_X1 U466 ( .A(n414), .B(n413), .ZN(n435) );
  XOR2_X1 U467 ( .A(KEYINPUT6), .B(G57GAT), .Z(n416) );
  XNOR2_X1 U468 ( .A(G1GAT), .B(G148GAT), .ZN(n415) );
  XNOR2_X1 U469 ( .A(n416), .B(n415), .ZN(n420) );
  XOR2_X1 U470 ( .A(KEYINPUT4), .B(KEYINPUT97), .Z(n418) );
  XNOR2_X1 U471 ( .A(KEYINPUT1), .B(KEYINPUT5), .ZN(n417) );
  XNOR2_X1 U472 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U473 ( .A(n420), .B(n419), .Z(n425) );
  XOR2_X1 U474 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n422) );
  NAND2_X1 U475 ( .A1(G225GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U476 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U477 ( .A(KEYINPUT100), .B(n423), .ZN(n424) );
  XNOR2_X1 U478 ( .A(n425), .B(n424), .ZN(n431) );
  XOR2_X1 U479 ( .A(G85GAT), .B(G155GAT), .Z(n429) );
  XOR2_X1 U480 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n427) );
  XNOR2_X1 U481 ( .A(G141GAT), .B(KEYINPUT95), .ZN(n426) );
  XNOR2_X1 U482 ( .A(n427), .B(n426), .ZN(n440) );
  XNOR2_X1 U483 ( .A(n440), .B(G162GAT), .ZN(n428) );
  XNOR2_X1 U484 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U485 ( .A(n431), .B(n430), .Z(n434) );
  XNOR2_X1 U486 ( .A(G29GAT), .B(n432), .ZN(n433) );
  XNOR2_X1 U487 ( .A(n434), .B(n433), .ZN(n490) );
  NOR2_X2 U488 ( .A1(n435), .A2(n490), .ZN(n566) );
  XOR2_X1 U489 ( .A(KEYINPUT93), .B(KEYINPUT96), .Z(n437) );
  NAND2_X1 U490 ( .A1(G228GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U492 ( .A(n438), .B(KEYINPUT92), .Z(n442) );
  XNOR2_X1 U493 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U494 ( .A(n442), .B(n441), .ZN(n446) );
  XOR2_X1 U495 ( .A(KEYINPUT22), .B(KEYINPUT91), .Z(n444) );
  XNOR2_X1 U496 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n443) );
  XNOR2_X1 U497 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U498 ( .A(n446), .B(n445), .Z(n450) );
  XNOR2_X1 U499 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U500 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U501 ( .A(n452), .B(n451), .ZN(n466) );
  NAND2_X1 U502 ( .A1(n566), .A2(n466), .ZN(n453) );
  XNOR2_X1 U503 ( .A(n453), .B(KEYINPUT55), .ZN(n454) );
  XNOR2_X1 U504 ( .A(n544), .B(KEYINPUT111), .ZN(n529) );
  NAND2_X1 U505 ( .A1(n288), .A2(n529), .ZN(n458) );
  XOR2_X1 U506 ( .A(G176GAT), .B(KEYINPUT56), .Z(n456) );
  XNOR2_X1 U507 ( .A(KEYINPUT124), .B(KEYINPUT57), .ZN(n455) );
  INV_X1 U508 ( .A(n490), .ZN(n514) );
  NOR2_X1 U509 ( .A1(n567), .A2(n570), .ZN(n487) );
  NAND2_X1 U510 ( .A1(n556), .A2(n552), .ZN(n459) );
  XNOR2_X1 U511 ( .A(n459), .B(KEYINPUT16), .ZN(n460) );
  XNOR2_X1 U512 ( .A(KEYINPUT89), .B(n460), .ZN(n473) );
  XOR2_X1 U513 ( .A(KEYINPUT27), .B(n517), .Z(n464) );
  NAND2_X1 U514 ( .A1(n464), .A2(n490), .ZN(n461) );
  XOR2_X1 U515 ( .A(KEYINPUT103), .B(n461), .Z(n539) );
  XOR2_X1 U516 ( .A(KEYINPUT28), .B(n466), .Z(n499) );
  NOR2_X1 U517 ( .A1(n539), .A2(n499), .ZN(n526) );
  NAND2_X1 U518 ( .A1(n524), .A2(n526), .ZN(n472) );
  NOR2_X1 U519 ( .A1(n496), .A2(n466), .ZN(n463) );
  XNOR2_X1 U520 ( .A(KEYINPUT104), .B(KEYINPUT26), .ZN(n462) );
  XNOR2_X1 U521 ( .A(n463), .B(n462), .ZN(n565) );
  NAND2_X1 U522 ( .A1(n464), .A2(n565), .ZN(n469) );
  INV_X1 U523 ( .A(n517), .ZN(n494) );
  NAND2_X1 U524 ( .A1(n494), .A2(n496), .ZN(n465) );
  NAND2_X1 U525 ( .A1(n466), .A2(n465), .ZN(n467) );
  XOR2_X1 U526 ( .A(KEYINPUT25), .B(n467), .Z(n468) );
  NAND2_X1 U527 ( .A1(n469), .A2(n468), .ZN(n470) );
  NAND2_X1 U528 ( .A1(n470), .A2(n514), .ZN(n471) );
  NAND2_X1 U529 ( .A1(n472), .A2(n471), .ZN(n484) );
  NAND2_X1 U530 ( .A1(n473), .A2(n484), .ZN(n474) );
  XNOR2_X1 U531 ( .A(n474), .B(KEYINPUT105), .ZN(n502) );
  NAND2_X1 U532 ( .A1(n487), .A2(n502), .ZN(n482) );
  NOR2_X1 U533 ( .A1(n514), .A2(n482), .ZN(n476) );
  XNOR2_X1 U534 ( .A(KEYINPUT106), .B(KEYINPUT34), .ZN(n475) );
  XNOR2_X1 U535 ( .A(n476), .B(n475), .ZN(n477) );
  XOR2_X1 U536 ( .A(G1GAT), .B(n477), .Z(G1324GAT) );
  NOR2_X1 U537 ( .A1(n517), .A2(n482), .ZN(n478) );
  XOR2_X1 U538 ( .A(G8GAT), .B(n478), .Z(G1325GAT) );
  NOR2_X1 U539 ( .A1(n524), .A2(n482), .ZN(n480) );
  XNOR2_X1 U540 ( .A(KEYINPUT107), .B(KEYINPUT35), .ZN(n479) );
  XNOR2_X1 U541 ( .A(n480), .B(n479), .ZN(n481) );
  XOR2_X1 U542 ( .A(G15GAT), .B(n481), .Z(G1326GAT) );
  INV_X1 U543 ( .A(n499), .ZN(n521) );
  NOR2_X1 U544 ( .A1(n521), .A2(n482), .ZN(n483) );
  XOR2_X1 U545 ( .A(G22GAT), .B(n483), .Z(G1327GAT) );
  XOR2_X1 U546 ( .A(KEYINPUT39), .B(KEYINPUT110), .Z(n492) );
  NAND2_X1 U547 ( .A1(n576), .A2(n484), .ZN(n485) );
  NOR2_X1 U548 ( .A1(n556), .A2(n485), .ZN(n486) );
  XOR2_X1 U549 ( .A(KEYINPUT37), .B(n486), .Z(n513) );
  NAND2_X1 U550 ( .A1(n487), .A2(n513), .ZN(n488) );
  XNOR2_X1 U551 ( .A(n488), .B(KEYINPUT38), .ZN(n489) );
  XNOR2_X1 U552 ( .A(KEYINPUT109), .B(n489), .ZN(n500) );
  NAND2_X1 U553 ( .A1(n490), .A2(n500), .ZN(n491) );
  XNOR2_X1 U554 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U555 ( .A(G29GAT), .B(n493), .ZN(G1328GAT) );
  NAND2_X1 U556 ( .A1(n500), .A2(n494), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n495), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U558 ( .A1(n500), .A2(n496), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n497), .B(KEYINPUT40), .ZN(n498) );
  XNOR2_X1 U560 ( .A(G43GAT), .B(n498), .ZN(G1330GAT) );
  NAND2_X1 U561 ( .A1(n500), .A2(n499), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n501), .B(G50GAT), .ZN(G1331GAT) );
  AND2_X1 U563 ( .A1(n567), .A2(n529), .ZN(n512) );
  NAND2_X1 U564 ( .A1(n502), .A2(n512), .ZN(n508) );
  NOR2_X1 U565 ( .A1(n514), .A2(n508), .ZN(n504) );
  XNOR2_X1 U566 ( .A(KEYINPUT42), .B(KEYINPUT112), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U568 ( .A(G57GAT), .B(n505), .Z(G1332GAT) );
  NOR2_X1 U569 ( .A1(n517), .A2(n508), .ZN(n506) );
  XOR2_X1 U570 ( .A(G64GAT), .B(n506), .Z(G1333GAT) );
  NOR2_X1 U571 ( .A1(n524), .A2(n508), .ZN(n507) );
  XOR2_X1 U572 ( .A(G71GAT), .B(n507), .Z(G1334GAT) );
  NOR2_X1 U573 ( .A1(n521), .A2(n508), .ZN(n510) );
  XNOR2_X1 U574 ( .A(KEYINPUT113), .B(KEYINPUT43), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U576 ( .A(G78GAT), .B(n511), .Z(G1335GAT) );
  NAND2_X1 U577 ( .A1(n513), .A2(n512), .ZN(n520) );
  NOR2_X1 U578 ( .A1(n514), .A2(n520), .ZN(n515) );
  XOR2_X1 U579 ( .A(G85GAT), .B(n515), .Z(n516) );
  XNOR2_X1 U580 ( .A(KEYINPUT114), .B(n516), .ZN(G1336GAT) );
  NOR2_X1 U581 ( .A1(n517), .A2(n520), .ZN(n518) );
  XOR2_X1 U582 ( .A(G92GAT), .B(n518), .Z(G1337GAT) );
  NOR2_X1 U583 ( .A1(n524), .A2(n520), .ZN(n519) );
  XOR2_X1 U584 ( .A(G99GAT), .B(n519), .Z(G1338GAT) );
  NOR2_X1 U585 ( .A1(n521), .A2(n520), .ZN(n522) );
  XOR2_X1 U586 ( .A(KEYINPUT44), .B(n522), .Z(n523) );
  XNOR2_X1 U587 ( .A(G106GAT), .B(n523), .ZN(G1339GAT) );
  NOR2_X1 U588 ( .A1(n524), .A2(n540), .ZN(n525) );
  NAND2_X1 U589 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U590 ( .A(KEYINPUT117), .B(n527), .ZN(n534) );
  NAND2_X1 U591 ( .A1(n554), .A2(n534), .ZN(n528) );
  XNOR2_X1 U592 ( .A(G113GAT), .B(n528), .ZN(G1340GAT) );
  XOR2_X1 U593 ( .A(G120GAT), .B(KEYINPUT49), .Z(n531) );
  NAND2_X1 U594 ( .A1(n534), .A2(n529), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n531), .B(n530), .ZN(G1341GAT) );
  NAND2_X1 U596 ( .A1(n534), .A2(n556), .ZN(n532) );
  XNOR2_X1 U597 ( .A(n532), .B(KEYINPUT50), .ZN(n533) );
  XNOR2_X1 U598 ( .A(G127GAT), .B(n533), .ZN(G1342GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n536) );
  INV_X1 U600 ( .A(n552), .ZN(n558) );
  NAND2_X1 U601 ( .A1(n534), .A2(n558), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n536), .B(n535), .ZN(n538) );
  XOR2_X1 U603 ( .A(G134GAT), .B(KEYINPUT118), .Z(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(G1343GAT) );
  NOR2_X1 U605 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U606 ( .A1(n565), .A2(n541), .ZN(n551) );
  NOR2_X1 U607 ( .A1(n567), .A2(n551), .ZN(n542) );
  XOR2_X1 U608 ( .A(KEYINPUT120), .B(n542), .Z(n543) );
  XNOR2_X1 U609 ( .A(G141GAT), .B(n543), .ZN(G1344GAT) );
  NOR2_X1 U610 ( .A1(n551), .A2(n544), .ZN(n548) );
  XOR2_X1 U611 ( .A(KEYINPUT52), .B(KEYINPUT121), .Z(n546) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1345GAT) );
  INV_X1 U615 ( .A(n556), .ZN(n574) );
  NOR2_X1 U616 ( .A1(n574), .A2(n551), .ZN(n549) );
  XOR2_X1 U617 ( .A(KEYINPUT122), .B(n549), .Z(n550) );
  XNOR2_X1 U618 ( .A(G155GAT), .B(n550), .ZN(G1346GAT) );
  NOR2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U620 ( .A(G162GAT), .B(n553), .Z(G1347GAT) );
  NAND2_X1 U621 ( .A1(n288), .A2(n554), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n555), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U623 ( .A1(n288), .A2(n556), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n557), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n561) );
  XOR2_X1 U626 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G190GAT), .ZN(G1351GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n564) );
  XNOR2_X1 U630 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n569) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n573) );
  NOR2_X1 U633 ( .A1(n567), .A2(n573), .ZN(n568) );
  XOR2_X1 U634 ( .A(n569), .B(n568), .Z(G1352GAT) );
  INV_X1 U635 ( .A(n573), .ZN(n577) );
  AND2_X1 U636 ( .A1(n570), .A2(n577), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(G1353GAT) );
  NOR2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U640 ( .A(G211GAT), .B(n575), .Z(G1354GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n579) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(n580), .ZN(G1355GAT) );
endmodule

