//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 1 1 1 1 1 0 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 0 0 0 0 0 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 1 1 0 0 0 0 0 1 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1246, new_n1247, new_n1248, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(new_n204), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  INV_X1    g0017(.A(G107), .ZN(new_n218));
  INV_X1    g0018(.A(G264), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n206), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n209), .B(new_n214), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT64), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n225), .A2(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G250), .B(G257), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT65), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT66), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n231), .B(new_n232), .Z(new_n233));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n233), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G50), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT67), .ZN(new_n241));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(KEYINPUT10), .ZN(new_n248));
  AND2_X1   g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  OAI21_X1  g0050(.A(KEYINPUT69), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT69), .ZN(new_n255));
  NAND2_X1  g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n251), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n259), .A2(G222), .A3(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n259), .A2(G223), .A3(G1698), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n261), .B(new_n262), .C1(new_n216), .C2(new_n259), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G41), .ZN(new_n266));
  INV_X1    g0066(.A(G45), .ZN(new_n267));
  AOI21_X1  g0067(.A(G1), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(G1), .A3(G13), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n268), .A2(new_n270), .A3(G274), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT68), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G274), .ZN(new_n274));
  INV_X1    g0074(.A(new_n212), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n274), .B1(new_n275), .B2(new_n269), .ZN(new_n276));
  AOI21_X1  g0076(.A(KEYINPUT68), .B1(new_n276), .B2(new_n268), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n264), .A2(new_n268), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n278), .B1(G226), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(KEYINPUT70), .B1(new_n265), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n265), .A2(KEYINPUT70), .A3(new_n280), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(G200), .A3(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT76), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n248), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n283), .ZN(new_n287));
  OAI21_X1  g0087(.A(G190), .B1(new_n287), .B2(new_n281), .ZN(new_n288));
  NAND3_X1  g0088(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n212), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT8), .B(G58), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT71), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n292), .B1(new_n253), .B2(G20), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n204), .A2(KEYINPUT71), .A3(G33), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n291), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G150), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G20), .A2(G33), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NOR3_X1   g0098(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n299));
  OAI22_X1  g0099(.A1(new_n296), .A2(new_n298), .B1(new_n299), .B2(new_n204), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n290), .B1(new_n295), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n303), .A2(new_n290), .ZN(new_n304));
  INV_X1    g0104(.A(G50), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n305), .B1(new_n203), .B2(G20), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n304), .A2(new_n306), .B1(new_n305), .B2(new_n303), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n301), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n308), .B(KEYINPUT9), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n288), .A2(new_n284), .A3(new_n309), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n286), .B(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G179), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(new_n287), .B2(new_n281), .ZN(new_n313));
  INV_X1    g0113(.A(G169), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n282), .A2(new_n314), .A3(new_n283), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n313), .A2(new_n315), .A3(new_n308), .ZN(new_n316));
  INV_X1    g0116(.A(G13), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n317), .A2(G1), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT74), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n318), .A2(new_n319), .A3(G20), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n302), .A2(KEYINPUT74), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n290), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n322), .B(G77), .C1(G1), .C2(new_n204), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n302), .B(new_n319), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n323), .B1(G77), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n290), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n291), .B1(KEYINPUT73), .B2(new_n298), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n328), .B1(KEYINPUT73), .B2(new_n298), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT15), .B(G87), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n293), .A2(new_n294), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n331), .A2(new_n332), .B1(G20), .B2(G77), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n327), .B1(new_n329), .B2(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n326), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n259), .A2(G232), .A3(new_n260), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n259), .A2(G238), .A3(G1698), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n258), .A2(G107), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT72), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n270), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n336), .A2(new_n337), .A3(KEYINPUT72), .A4(new_n338), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n279), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n273), .A2(new_n277), .B1(new_n344), .B2(new_n217), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n335), .B1(new_n347), .B2(new_n314), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n345), .B1(new_n341), .B2(new_n342), .ZN(new_n349));
  AND3_X1   g0149(.A1(new_n349), .A2(KEYINPUT75), .A3(new_n312), .ZN(new_n350));
  AOI21_X1  g0150(.A(KEYINPUT75), .B1(new_n349), .B2(new_n312), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n348), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n349), .A2(G190), .ZN(new_n353));
  INV_X1    g0153(.A(G200), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n353), .B(new_n335), .C1(new_n354), .C2(new_n349), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n311), .A2(new_n316), .A3(new_n352), .A4(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n278), .B1(G238), .B2(new_n279), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n251), .A2(new_n257), .A3(G226), .A4(new_n260), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n251), .A2(new_n257), .A3(G232), .A4(G1698), .ZN(new_n359));
  NAND2_X1  g0159(.A1(G33), .A2(G97), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  AND3_X1   g0161(.A1(new_n361), .A2(KEYINPUT77), .A3(new_n264), .ZN(new_n362));
  AOI21_X1  g0162(.A(KEYINPUT77), .B1(new_n361), .B2(new_n264), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n357), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT13), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT13), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n357), .B(new_n366), .C1(new_n362), .C2(new_n363), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  XOR2_X1   g0168(.A(KEYINPUT79), .B(KEYINPUT14), .Z(new_n369));
  NAND3_X1  g0169(.A1(new_n368), .A2(G169), .A3(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT80), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n368), .A2(G169), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT14), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n368), .A2(KEYINPUT80), .A3(G169), .A4(new_n369), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n365), .A2(G179), .A3(new_n367), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n372), .A2(new_n374), .A3(new_n375), .A4(new_n376), .ZN(new_n377));
  XNOR2_X1  g0177(.A(KEYINPUT78), .B(KEYINPUT12), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(new_n325), .B2(G68), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT12), .ZN(new_n380));
  INV_X1    g0180(.A(G68), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n318), .A2(new_n380), .A3(G20), .A4(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n332), .A2(G77), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n297), .A2(G50), .B1(G20), .B2(new_n381), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n327), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  OR2_X1    g0186(.A1(new_n386), .A2(KEYINPUT11), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n322), .B(G68), .C1(G1), .C2(new_n204), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n386), .A2(KEYINPUT11), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n383), .A2(new_n387), .A3(new_n388), .A4(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n377), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n390), .ZN(new_n392));
  INV_X1    g0192(.A(G190), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n392), .B1(new_n368), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n354), .B1(new_n365), .B2(new_n367), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n391), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(G58), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n399), .A2(new_n381), .ZN(new_n400));
  NOR2_X1   g0200(.A1(G58), .A2(G68), .ZN(new_n401));
  OAI21_X1  g0201(.A(G20), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n297), .A2(G159), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n249), .A2(new_n250), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n406), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NOR3_X1   g0208(.A1(new_n249), .A2(new_n250), .A3(KEYINPUT69), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n255), .B1(new_n254), .B2(new_n256), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n204), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT7), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n408), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n405), .B1(new_n413), .B2(new_n381), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT16), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(KEYINPUT81), .A3(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT81), .ZN(new_n417));
  AOI21_X1  g0217(.A(G20), .B1(new_n251), .B2(new_n257), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n407), .B1(new_n418), .B2(KEYINPUT7), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n404), .B1(new_n419), .B2(G68), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n417), .B1(new_n420), .B2(KEYINPUT16), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n254), .A2(new_n256), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n412), .B1(new_n422), .B2(G20), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n407), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n404), .B1(new_n424), .B2(G68), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n327), .B1(new_n425), .B2(KEYINPUT16), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n416), .A2(new_n421), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n291), .B1(new_n203), .B2(G20), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n428), .A2(new_n304), .B1(new_n303), .B2(new_n291), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT18), .ZN(new_n431));
  INV_X1    g0231(.A(G223), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n260), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(G226), .B2(new_n260), .ZN(new_n434));
  INV_X1    g0234(.A(G87), .ZN(new_n435));
  OAI22_X1  g0235(.A1(new_n434), .A2(new_n406), .B1(new_n253), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n264), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n264), .A2(new_n268), .A3(new_n235), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n271), .A2(new_n272), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n276), .A2(KEYINPUT68), .A3(new_n268), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT82), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n437), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AOI211_X1 g0243(.A(KEYINPUT82), .B(new_n438), .C1(new_n439), .C2(new_n440), .ZN(new_n444));
  OAI21_X1  g0244(.A(G169), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT82), .B1(new_n278), .B2(new_n438), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n441), .A2(new_n442), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n446), .A2(G179), .A3(new_n447), .A4(new_n437), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n430), .A2(new_n431), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n431), .B1(new_n430), .B2(new_n449), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n354), .B1(new_n443), .B2(new_n444), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n446), .A2(new_n393), .A3(new_n447), .A4(new_n437), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n427), .A2(new_n455), .A3(new_n429), .ZN(new_n456));
  XNOR2_X1  g0256(.A(new_n456), .B(KEYINPUT17), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(G238), .A2(G1698), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n459), .B1(new_n217), .B2(G1698), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n422), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G116), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n270), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n267), .A2(G1), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n276), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G250), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n270), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n314), .B1(new_n463), .B2(new_n469), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n276), .A2(new_n464), .B1(new_n467), .B2(new_n270), .ZN(new_n471));
  INV_X1    g0271(.A(new_n462), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n472), .B1(new_n460), .B2(new_n422), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n471), .B(new_n312), .C1(new_n473), .C2(new_n270), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n422), .A2(new_n204), .A3(G68), .ZN(new_n476));
  INV_X1    g0276(.A(G97), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n477), .B1(new_n293), .B2(new_n294), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT19), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n204), .B1(new_n360), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n435), .A2(new_n477), .A3(new_n218), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n480), .A2(KEYINPUT85), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(KEYINPUT85), .B1(new_n480), .B2(new_n481), .ZN(new_n483));
  OAI221_X1 g0283(.A(new_n476), .B1(new_n478), .B2(KEYINPUT19), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n484), .A2(new_n290), .B1(new_n324), .B2(new_n330), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n304), .B1(G1), .B2(new_n253), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n331), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n475), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n482), .A2(new_n483), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n476), .B1(new_n478), .B2(KEYINPUT19), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n290), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n487), .A2(G87), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n324), .A2(new_n330), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(G200), .B1(new_n463), .B2(new_n469), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n471), .B(G190), .C1(new_n473), .C2(new_n270), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(KEYINPUT86), .B1(new_n489), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n492), .A2(new_n488), .A3(new_n494), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n501), .A2(new_n470), .A3(new_n474), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT86), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n502), .B(new_n503), .C1(new_n495), .C2(new_n498), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT24), .ZN(new_n506));
  NOR3_X1   g0306(.A1(new_n435), .A2(KEYINPUT22), .A3(G20), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n259), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n422), .A2(new_n204), .A3(G87), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT22), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT23), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n512), .B1(new_n204), .B2(G107), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n218), .A2(KEYINPUT23), .A3(G20), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n513), .A2(new_n514), .B1(new_n472), .B2(new_n204), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n506), .B1(new_n511), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n515), .ZN(new_n517));
  AOI211_X1 g0317(.A(KEYINPUT24), .B(new_n517), .C1(new_n508), .C2(new_n510), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n290), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n303), .A2(new_n218), .ZN(new_n520));
  XNOR2_X1  g0320(.A(new_n520), .B(KEYINPUT25), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n521), .B1(new_n487), .B2(G107), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g0323(.A(KEYINPUT5), .B(G41), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n276), .A2(new_n464), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n464), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n270), .ZN(new_n527));
  NOR2_X1   g0327(.A1(G250), .A2(G1698), .ZN(new_n528));
  INV_X1    g0328(.A(G257), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n528), .B1(new_n529), .B2(G1698), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n530), .A2(new_n422), .B1(G33), .B2(G294), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT90), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n264), .B1(new_n531), .B2(new_n532), .ZN(new_n535));
  OAI221_X1 g0335(.A(new_n525), .B1(new_n219), .B2(new_n527), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n314), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n527), .A2(new_n219), .ZN(new_n538));
  INV_X1    g0338(.A(new_n535), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n538), .B1(new_n539), .B2(new_n533), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n540), .A2(new_n312), .A3(new_n525), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n523), .A2(new_n537), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n536), .A2(G200), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n540), .A2(G190), .A3(new_n525), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n519), .A2(new_n543), .A3(new_n544), .A4(new_n522), .ZN(new_n545));
  AND3_X1   g0345(.A1(new_n505), .A2(new_n542), .A3(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(G116), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n547), .B1(new_n203), .B2(G33), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n322), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n324), .A2(new_n547), .ZN(new_n550));
  NAND2_X1  g0350(.A1(G33), .A2(G283), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n551), .B(new_n204), .C1(G33), .C2(new_n477), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n547), .A2(G20), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n552), .A2(new_n290), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT20), .ZN(new_n555));
  AND2_X1   g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n554), .A2(new_n555), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n549), .B(new_n550), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT88), .ZN(new_n559));
  XNOR2_X1  g0359(.A(new_n554), .B(new_n555), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT88), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n560), .A2(new_n561), .A3(new_n550), .A4(new_n549), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G169), .ZN(new_n564));
  INV_X1    g0364(.A(G303), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n251), .B2(new_n257), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n219), .A2(G1698), .ZN(new_n567));
  OAI221_X1 g0367(.A(new_n567), .B1(G257), .B2(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n264), .B1(new_n566), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n264), .B1(new_n464), .B2(new_n524), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n524), .A2(new_n464), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n571), .A2(G270), .B1(new_n572), .B2(new_n276), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT87), .ZN(new_n575));
  XNOR2_X1  g0375(.A(new_n574), .B(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(KEYINPUT21), .B1(new_n564), .B2(new_n576), .ZN(new_n577));
  XNOR2_X1  g0377(.A(new_n574), .B(KEYINPUT87), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT21), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n314), .B1(new_n559), .B2(new_n562), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n574), .A2(new_n312), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n563), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(KEYINPUT89), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT89), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n563), .A2(new_n585), .A3(new_n582), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n577), .A2(new_n581), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n563), .B1(new_n576), .B2(G190), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(new_n354), .B2(new_n576), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n302), .A2(G97), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(new_n486), .B2(new_n477), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT6), .ZN(new_n594));
  NOR3_X1   g0394(.A1(new_n594), .A2(new_n477), .A3(G107), .ZN(new_n595));
  XNOR2_X1  g0395(.A(G97), .B(G107), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n595), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  OAI22_X1  g0397(.A1(new_n597), .A2(new_n204), .B1(new_n216), .B2(new_n298), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n598), .B1(new_n419), .B2(G107), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n593), .B1(new_n599), .B2(new_n327), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n251), .A2(new_n257), .A3(G250), .A4(G1698), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n260), .A2(G244), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT4), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n251), .A2(new_n257), .A3(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n603), .B1(new_n406), .B2(new_n602), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n601), .A2(new_n605), .A3(new_n551), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n264), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n525), .B1(new_n527), .B2(new_n529), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n314), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n609), .B1(new_n607), .B2(new_n264), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n312), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n600), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(KEYINPUT84), .ZN(new_n616));
  INV_X1    g0416(.A(new_n598), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(new_n413), .B2(new_n218), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n592), .B1(new_n618), .B2(new_n290), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n613), .A2(G190), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT83), .ZN(new_n621));
  OAI21_X1  g0421(.A(G200), .B1(new_n613), .B2(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n611), .A2(KEYINPUT83), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n619), .B(new_n620), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT84), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n600), .A2(new_n612), .A3(new_n625), .A4(new_n614), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n616), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n546), .A2(new_n587), .A3(new_n589), .A4(new_n628), .ZN(new_n629));
  NOR4_X1   g0429(.A1(new_n356), .A2(new_n398), .A3(new_n458), .A4(new_n629), .ZN(G372));
  NOR3_X1   g0430(.A1(new_n356), .A2(new_n398), .A3(new_n458), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n489), .A2(new_n499), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n545), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n627), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n584), .A2(new_n586), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n579), .B1(new_n578), .B2(new_n580), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n635), .B(new_n542), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n616), .A2(new_n626), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n640), .A2(new_n505), .A3(KEYINPUT26), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT26), .ZN(new_n642));
  INV_X1    g0442(.A(new_n632), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n642), .B1(new_n643), .B2(new_n615), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n639), .A2(new_n645), .A3(new_n502), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n631), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n316), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n391), .A2(new_n352), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n397), .A2(new_n457), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n452), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n648), .B1(new_n651), .B2(new_n311), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n647), .A2(new_n652), .ZN(G369));
  AND2_X1   g0453(.A1(new_n587), .A2(new_n589), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n318), .A2(new_n204), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n655), .B(KEYINPUT91), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT27), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(new_n659), .A3(G213), .ZN(new_n660));
  INV_X1    g0460(.A(G343), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n563), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n654), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n587), .B2(new_n663), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT92), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n665), .A2(new_n666), .A3(G330), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n666), .B1(new_n665), .B2(G330), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n523), .A2(new_n662), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n542), .A2(new_n545), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g0471(.A(new_n671), .B(KEYINPUT93), .Z(new_n672));
  INV_X1    g0472(.A(new_n542), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n662), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n669), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n672), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n587), .A2(new_n662), .ZN(new_n680));
  INV_X1    g0480(.A(new_n662), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n679), .A2(new_n680), .B1(new_n673), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n678), .A2(new_n682), .ZN(G399));
  INV_X1    g0483(.A(new_n207), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(G41), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(new_n203), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n481), .A2(G116), .ZN(new_n688));
  INV_X1    g0488(.A(new_n685), .ZN(new_n689));
  OAI22_X1  g0489(.A1(new_n687), .A2(new_n688), .B1(new_n210), .B2(new_n689), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT28), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n489), .B1(new_n634), .B2(new_n638), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n662), .B1(new_n692), .B2(new_n645), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n693), .A2(KEYINPUT29), .ZN(new_n694));
  AOI22_X1  g0494(.A1(new_n616), .A2(new_n626), .B1(new_n500), .B2(new_n504), .ZN(new_n695));
  OAI21_X1  g0495(.A(KEYINPUT96), .B1(new_n695), .B2(KEYINPUT26), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n640), .A2(new_n505), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT96), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(new_n698), .A3(new_n642), .ZN(new_n699));
  OR3_X1    g0499(.A1(new_n643), .A2(new_n642), .A3(new_n615), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n696), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n662), .B1(new_n701), .B2(new_n692), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(KEYINPUT29), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n694), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n654), .A2(new_n628), .A3(new_n546), .A4(new_n681), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n463), .A2(new_n469), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n582), .A2(new_n540), .A3(new_n613), .A4(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT94), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(KEYINPUT30), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n706), .A2(G179), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n578), .A2(new_n611), .A3(new_n536), .A4(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT30), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n707), .A2(new_n708), .A3(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n710), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n715), .A2(KEYINPUT31), .A3(new_n662), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(KEYINPUT95), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n705), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n715), .A2(new_n662), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT31), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(KEYINPUT95), .B2(new_n716), .ZN(new_n722));
  OAI21_X1  g0522(.A(G330), .B1(new_n718), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n704), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n691), .B1(new_n725), .B2(G1), .ZN(G364));
  NOR3_X1   g0526(.A1(new_n317), .A2(new_n267), .A3(G20), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT97), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n687), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OAI211_X1 g0530(.A(new_n669), .B(new_n730), .C1(G330), .C2(new_n665), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n259), .A2(G355), .A3(new_n207), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n732), .B1(G116), .B2(new_n207), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n243), .A2(new_n267), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n684), .A2(new_n422), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n736), .B1(new_n267), .B2(new_n211), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n733), .B1(new_n734), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G13), .A2(G33), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G20), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n212), .B1(G20), .B2(new_n314), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n729), .B1(new_n738), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n204), .A2(G179), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G190), .A2(G200), .ZN(new_n747));
  AND2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OR2_X1    g0548(.A1(new_n748), .A2(KEYINPUT98), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(KEYINPUT98), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n746), .A2(new_n393), .A3(G200), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n752), .A2(G329), .B1(G283), .B2(new_n754), .ZN(new_n755));
  XOR2_X1   g0555(.A(new_n755), .B(KEYINPUT101), .Z(new_n756));
  NOR2_X1   g0556(.A1(new_n204), .A2(new_n312), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G200), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n393), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(G190), .ZN(new_n760));
  XNOR2_X1  g0560(.A(KEYINPUT33), .B(G317), .ZN(new_n761));
  AOI22_X1  g0561(.A1(G326), .A2(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n757), .A2(G190), .A3(new_n354), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n757), .A2(new_n747), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n764), .A2(G322), .B1(new_n766), .B2(G311), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n393), .A2(G179), .A3(G200), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n204), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n746), .A2(G190), .A3(G200), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n770), .A2(G294), .B1(new_n772), .B2(G303), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n762), .A2(new_n258), .A3(new_n767), .A4(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G159), .ZN(new_n775));
  OR3_X1    g0575(.A1(new_n751), .A2(KEYINPUT32), .A3(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(KEYINPUT32), .B1(new_n751), .B2(new_n775), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n258), .B1(G87), .B2(new_n772), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n776), .B(new_n777), .C1(KEYINPUT99), .C2(new_n778), .ZN(new_n779));
  AOI22_X1  g0579(.A1(G97), .A2(new_n770), .B1(new_n760), .B2(G68), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT100), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n778), .A2(KEYINPUT99), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n753), .A2(new_n218), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n763), .A2(new_n399), .B1(new_n765), .B2(new_n216), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n783), .B(new_n784), .C1(G50), .C2(new_n759), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n781), .A2(new_n782), .A3(new_n785), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n756), .A2(new_n774), .B1(new_n779), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n745), .B1(new_n787), .B2(new_n742), .ZN(new_n788));
  INV_X1    g0588(.A(new_n741), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n788), .B1(new_n665), .B2(new_n789), .ZN(new_n790));
  AND2_X1   g0590(.A1(new_n731), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(G396));
  INV_X1    g0592(.A(new_n742), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(new_n740), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n729), .B1(G77), .B2(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n764), .A2(G143), .B1(new_n766), .B2(G159), .ZN(new_n796));
  INV_X1    g0596(.A(new_n760), .ZN(new_n797));
  INV_X1    g0597(.A(G137), .ZN(new_n798));
  INV_X1    g0598(.A(new_n759), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n796), .B1(new_n797), .B2(new_n296), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT34), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n752), .A2(G132), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n769), .A2(new_n399), .B1(new_n771), .B2(new_n305), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n406), .B(new_n805), .C1(G68), .C2(new_n754), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n802), .A2(new_n803), .A3(new_n804), .A4(new_n806), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n799), .A2(new_n565), .B1(new_n771), .B2(new_n218), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(G283), .B2(new_n760), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n752), .A2(G311), .ZN(new_n810));
  INV_X1    g0610(.A(G294), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n763), .A2(new_n811), .B1(new_n765), .B2(new_n547), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(new_n259), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n753), .A2(new_n435), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(G97), .B2(new_n770), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n809), .A2(new_n810), .A3(new_n813), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n807), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n795), .B1(new_n817), .B2(new_n742), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n681), .A2(new_n335), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n352), .A2(new_n355), .A3(new_n820), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n348), .B(new_n819), .C1(new_n350), .C2(new_n351), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n818), .B1(new_n823), .B2(new_n740), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT102), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n646), .A2(new_n823), .A3(new_n681), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(KEYINPUT103), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT103), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n693), .A2(new_n828), .A3(new_n823), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n693), .A2(new_n823), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n723), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n730), .ZN(new_n834));
  NOR3_X1   g0634(.A1(new_n831), .A2(new_n723), .A3(new_n832), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n825), .B1(new_n834), .B2(new_n835), .ZN(G384));
  INV_X1    g0636(.A(new_n597), .ZN(new_n837));
  OR2_X1    g0637(.A1(new_n837), .A2(KEYINPUT35), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(KEYINPUT35), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n838), .A2(G116), .A3(new_n213), .A4(new_n839), .ZN(new_n840));
  XOR2_X1   g0640(.A(new_n840), .B(KEYINPUT36), .Z(new_n841));
  OAI211_X1 g0641(.A(new_n211), .B(G77), .C1(new_n399), .C2(new_n381), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n305), .A2(G68), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n203), .B(G13), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT38), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT37), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n426), .B1(KEYINPUT16), .B2(new_n425), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(new_n429), .ZN(new_n849));
  INV_X1    g0649(.A(new_n660), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n849), .B1(new_n449), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n847), .B1(new_n851), .B2(new_n456), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n430), .A2(new_n449), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n456), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n430), .A2(new_n850), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n847), .ZN(new_n856));
  OAI21_X1  g0656(.A(KEYINPUT104), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  AND3_X1   g0657(.A1(new_n427), .A2(new_n429), .A3(new_n455), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n427), .A2(new_n429), .B1(new_n445), .B2(new_n448), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT104), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT37), .B1(new_n430), .B2(new_n850), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n852), .B1(new_n857), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n849), .A2(new_n850), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(new_n452), .B2(new_n457), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n846), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n852), .ZN(new_n868));
  AND4_X1   g0668(.A1(new_n861), .A2(new_n862), .A3(new_n853), .A4(new_n456), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n861), .B1(new_n860), .B2(new_n862), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n865), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n458), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n871), .A2(KEYINPUT38), .A3(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT105), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n867), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  OAI211_X1 g0676(.A(KEYINPUT105), .B(new_n846), .C1(new_n864), .C2(new_n866), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT39), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n377), .A2(new_n390), .A3(new_n681), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT39), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n847), .B1(new_n860), .B2(new_n855), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n883), .B1(new_n857), .B2(new_n863), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n855), .B1(new_n452), .B2(new_n457), .ZN(new_n885));
  OAI211_X1 g0685(.A(KEYINPUT106), .B(new_n846), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n874), .ZN(new_n887));
  INV_X1    g0687(.A(new_n855), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT37), .B1(new_n854), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n869), .B2(new_n870), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n458), .A2(new_n888), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT38), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n892), .A2(KEYINPUT106), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n882), .B1(new_n887), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n879), .A2(new_n881), .A3(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n452), .A2(new_n850), .ZN(new_n896));
  INV_X1    g0696(.A(new_n878), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n662), .A2(new_n390), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n391), .A2(new_n397), .A3(new_n898), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n390), .B(new_n662), .C1(new_n377), .C2(new_n396), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n352), .A2(new_n662), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n902), .B1(new_n830), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n896), .B1(new_n897), .B2(new_n904), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n895), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n631), .A2(new_n694), .A3(new_n703), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n652), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n906), .B(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT40), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n721), .A2(new_n716), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n911), .A2(new_n705), .B1(new_n821), .B2(new_n822), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n901), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n910), .B1(new_n878), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n846), .B1(new_n884), .B2(new_n885), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT106), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(new_n874), .A3(new_n886), .ZN(new_n918));
  AND3_X1   g0718(.A1(new_n912), .A2(new_n901), .A3(KEYINPUT40), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n914), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n911), .A2(new_n705), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n631), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(G330), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(new_n921), .B2(new_n923), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n909), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(G1), .B1(new_n317), .B2(G20), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n909), .B2(new_n925), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n845), .B1(new_n926), .B2(new_n928), .ZN(G367));
  OAI221_X1 g0729(.A(new_n743), .B1(new_n207), .B2(new_n330), .C1(new_n233), .C2(new_n736), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT111), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n730), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n751), .A2(new_n798), .ZN(new_n933));
  OAI221_X1 g0733(.A(new_n259), .B1(new_n305), .B2(new_n765), .C1(new_n296), .C2(new_n763), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n753), .A2(new_n216), .B1(new_n771), .B2(new_n399), .ZN(new_n935));
  NOR3_X1   g0735(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n770), .A2(G68), .ZN(new_n937));
  AOI22_X1  g0737(.A1(G143), .A2(new_n759), .B1(new_n760), .B2(G159), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(G311), .ZN(new_n940));
  OAI221_X1 g0740(.A(new_n406), .B1(new_n565), .B2(new_n763), .C1(new_n799), .C2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(G283), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n769), .A2(new_n218), .B1(new_n765), .B2(new_n942), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n943), .A2(KEYINPUT112), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n797), .A2(new_n811), .B1(new_n477), .B2(new_n753), .ZN(new_n945));
  NOR3_X1   g0745(.A1(new_n941), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(KEYINPUT112), .B2(new_n943), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n772), .A2(KEYINPUT46), .A3(G116), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT46), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n771), .B2(new_n547), .ZN(new_n950));
  INV_X1    g0750(.A(G317), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n948), .B(new_n950), .C1(new_n751), .C2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n939), .B1(new_n947), .B2(new_n952), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n953), .B(KEYINPUT47), .Z(new_n954));
  OAI221_X1 g0754(.A(new_n932), .B1(new_n931), .B2(new_n930), .C1(new_n954), .C2(new_n793), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n662), .A2(new_n495), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n632), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n502), .B2(new_n956), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n958), .A2(new_n789), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n955), .A2(new_n959), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n675), .A2(new_n680), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n679), .A2(new_n680), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n669), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n961), .B(new_n962), .C1(new_n667), .C2(new_n668), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n725), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(KEYINPUT110), .ZN(new_n969));
  OR3_X1    g0769(.A1(new_n966), .A2(KEYINPUT110), .A3(new_n724), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n628), .B1(new_n619), .B2(new_n681), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n615), .A2(new_n681), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n682), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT45), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n974), .B(new_n975), .ZN(new_n976));
  XOR2_X1   g0776(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  OR3_X1    g0778(.A1(new_n682), .A2(new_n973), .A3(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n978), .B1(new_n682), .B2(new_n973), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n976), .A2(new_n678), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n974), .A2(new_n975), .ZN(new_n982));
  AOI21_X1  g0782(.A(KEYINPUT45), .B1(new_n682), .B2(new_n973), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n979), .B(new_n980), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n677), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n969), .A2(new_n970), .A3(new_n981), .A4(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n725), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n685), .B(KEYINPUT41), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n728), .A2(new_n203), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n677), .A2(new_n973), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(KEYINPUT108), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT108), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n677), .A2(new_n994), .A3(new_n973), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n962), .B1(new_n971), .B2(new_n972), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT107), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1002), .A2(KEYINPUT42), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n640), .B1(new_n973), .B2(new_n673), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1004), .A2(new_n662), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(new_n1002), .B2(KEYINPUT42), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n1003), .A2(new_n1006), .B1(KEYINPUT43), .B2(new_n958), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n996), .A2(new_n997), .ZN(new_n1008));
  AND3_X1   g0808(.A1(new_n999), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1007), .B1(new_n999), .B2(new_n1008), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n960), .B1(new_n991), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(G387));
  NAND2_X1  g0813(.A1(new_n966), .A2(new_n724), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n968), .A2(new_n685), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n990), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n676), .A2(new_n741), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n406), .B1(new_n753), .B2(new_n547), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n764), .A2(G317), .B1(new_n766), .B2(G303), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n759), .A2(G322), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1019), .B(new_n1020), .C1(new_n940), .C2(new_n797), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT48), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n770), .A2(G283), .B1(new_n772), .B2(G294), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT49), .Z(new_n1027));
  AOI211_X1 g0827(.A(new_n1018), .B(new_n1027), .C1(G326), .C2(new_n752), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n751), .A2(new_n296), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n770), .A2(new_n331), .B1(new_n772), .B2(G77), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n291), .B2(new_n797), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n422), .B1(new_n765), .B2(new_n381), .C1(new_n305), .C2(new_n763), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n799), .A2(new_n775), .B1(new_n753), .B2(new_n477), .ZN(new_n1033));
  NOR4_X1   g0833(.A1(new_n1029), .A2(new_n1031), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n742), .B1(new_n1028), .B2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n259), .A2(new_n207), .A3(new_n688), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n291), .A2(G50), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT50), .ZN(new_n1038));
  AOI211_X1 g0838(.A(G45), .B(new_n688), .C1(G68), .C2(G77), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n736), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n238), .A2(new_n267), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1036), .B1(G107), .B2(new_n207), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT113), .ZN(new_n1044));
  AND2_X1   g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n743), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1035), .B(new_n729), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT114), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n967), .A2(new_n1016), .B1(new_n1017), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1015), .A2(new_n1049), .ZN(G393));
  NAND3_X1  g0850(.A1(new_n981), .A2(new_n985), .A3(new_n1016), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n743), .B1(new_n477), .B2(new_n207), .C1(new_n736), .C2(new_n246), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n729), .A2(new_n1052), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n799), .A2(new_n296), .B1(new_n775), .B2(new_n763), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT51), .Z(new_n1055));
  NAND2_X1  g0855(.A1(new_n752), .A2(G143), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n771), .A2(new_n381), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n769), .A2(new_n216), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n1057), .B(new_n1058), .C1(G50), .C2(new_n760), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n291), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n406), .B(new_n814), .C1(new_n1060), .C2(new_n766), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1056), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G116), .A2(new_n770), .B1(new_n760), .B2(G303), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n752), .A2(G322), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n783), .B1(G283), .B2(new_n772), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n259), .B1(G294), .B2(new_n766), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G317), .A2(new_n759), .B1(new_n764), .B2(G311), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT52), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n1055), .A2(new_n1062), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1053), .B1(new_n1070), .B2(new_n742), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n973), .B2(new_n789), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1051), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n981), .A2(new_n985), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n689), .B1(new_n1075), .B2(new_n968), .ZN(new_n1076));
  AND3_X1   g0876(.A1(new_n986), .A2(new_n1076), .A3(KEYINPUT115), .ZN(new_n1077));
  AOI21_X1  g0877(.A(KEYINPUT115), .B1(new_n986), .B2(new_n1076), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1074), .B1(new_n1077), .B2(new_n1078), .ZN(G390));
  INV_X1    g0879(.A(new_n903), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n827), .B2(new_n829), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n880), .B1(new_n1081), .B2(new_n902), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n857), .A2(new_n863), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n866), .B1(new_n1083), .B2(new_n868), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n892), .A2(KEYINPUT106), .B1(new_n1084), .B2(KEYINPUT38), .ZN(new_n1085));
  AOI21_X1  g0885(.A(KEYINPUT39), .B1(new_n1085), .B2(new_n917), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n882), .B1(new_n876), .B2(new_n877), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1082), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  OAI211_X1 g0888(.A(G330), .B(new_n823), .C1(new_n718), .C2(new_n722), .ZN(new_n1089));
  OR2_X1    g0889(.A1(new_n1089), .A2(new_n902), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1080), .B1(new_n702), .B2(new_n823), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n918), .B(new_n880), .C1(new_n902), .C2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1088), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n887), .A2(new_n893), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n880), .B1(new_n1091), .B2(new_n902), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n879), .A2(new_n894), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1096), .B1(new_n1097), .B2(new_n1082), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n912), .A2(new_n901), .A3(G330), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1093), .B(new_n1016), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1097), .A2(new_n739), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n729), .B1(new_n1060), .B2(new_n794), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n753), .A2(new_n305), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n797), .A2(new_n798), .B1(new_n775), .B2(new_n769), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n1103), .B(new_n1104), .C1(G128), .C2(new_n759), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n771), .A2(new_n296), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT53), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n752), .A2(G125), .ZN(new_n1108));
  INV_X1    g0908(.A(G132), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(KEYINPUT54), .B(G143), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n763), .A2(new_n1109), .B1(new_n765), .B2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1111), .A2(new_n258), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1105), .A2(new_n1107), .A3(new_n1108), .A4(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1058), .B1(G107), .B2(new_n760), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n942), .B2(new_n799), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n763), .A2(new_n547), .B1(new_n765), .B2(new_n477), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1116), .A2(new_n259), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n772), .A2(G87), .B1(new_n754), .B2(G68), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1117), .B(new_n1118), .C1(new_n751), .C2(new_n811), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1113), .B1(new_n1115), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1102), .B1(new_n1120), .B2(new_n742), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1101), .A2(new_n1121), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n1100), .A2(KEYINPUT117), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(KEYINPUT117), .B1(new_n1100), .B2(new_n1122), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1093), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1089), .A2(new_n902), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n1099), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n831), .B2(new_n1080), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n912), .A2(G330), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n902), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1090), .A2(new_n1091), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1129), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n631), .A2(G330), .A3(new_n922), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n907), .A2(new_n1134), .A3(new_n652), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n689), .B1(new_n1126), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1135), .B1(new_n1129), .B2(new_n1132), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1093), .B(new_n1139), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1140));
  AOI21_X1  g0940(.A(KEYINPUT116), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n1088), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1099), .B1(new_n1088), .B2(new_n1092), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1137), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  AND4_X1   g0944(.A1(KEYINPUT116), .A2(new_n1144), .A3(new_n685), .A4(new_n1140), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1125), .B1(new_n1141), .B2(new_n1145), .ZN(G378));
  NAND2_X1  g0946(.A1(new_n1140), .A2(new_n1136), .ZN(new_n1147));
  INV_X1    g0947(.A(G330), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(new_n918), .B2(new_n919), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n914), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n850), .A2(new_n308), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n311), .A2(new_n316), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1151), .B1(new_n311), .B2(new_n316), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  OR3_X1    g0956(.A1(new_n1153), .A2(new_n1154), .A3(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1156), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1150), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1149), .A2(new_n914), .A3(new_n1159), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n906), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n895), .A2(new_n905), .ZN(new_n1164));
  AND3_X1   g0964(.A1(new_n1149), .A2(new_n914), .A3(new_n1159), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1159), .B1(new_n1149), .B2(new_n914), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1164), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1163), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1147), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT57), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1170), .B1(new_n1163), .B2(new_n1167), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n689), .B1(new_n1172), .B2(new_n1147), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1174));
  NOR3_X1   g0974(.A1(new_n1165), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n1161), .A2(new_n1162), .B1(new_n895), .B2(new_n905), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1016), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1160), .A2(new_n739), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n729), .B1(G50), .B2(new_n794), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n477), .A2(new_n797), .B1(new_n799), .B2(new_n547), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(G58), .B2(new_n754), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n764), .A2(G107), .B1(new_n766), .B2(new_n331), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n937), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(G283), .B2(new_n752), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n266), .B(new_n406), .C1(new_n771), .C2(new_n216), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT118), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1181), .A2(new_n1184), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT58), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n406), .A2(new_n266), .ZN(new_n1189));
  AOI21_X1  g0989(.A(G50), .B1(new_n253), .B2(new_n266), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n1187), .A2(new_n1188), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n759), .A2(G125), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n797), .B2(new_n1109), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n764), .A2(G128), .B1(new_n766), .B2(G137), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n771), .B2(new_n1110), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n1193), .B(new_n1195), .C1(G150), .C2(new_n770), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT59), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1198), .A2(KEYINPUT119), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n752), .A2(G124), .ZN(new_n1200));
  AOI211_X1 g1000(.A(G33), .B(G41), .C1(new_n754), .C2(G159), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT119), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1200), .B(new_n1201), .C1(new_n1197), .C2(new_n1202), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1191), .B1(new_n1188), .B2(new_n1187), .C1(new_n1199), .C2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1179), .B1(new_n1204), .B2(new_n742), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1178), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1177), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1174), .A2(new_n1208), .ZN(G375));
  NAND2_X1  g1009(.A1(new_n1133), .A2(new_n1016), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n729), .B1(G68), .B2(new_n794), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n799), .A2(new_n1109), .B1(new_n771), .B2(new_n775), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(G50), .B2(new_n770), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n752), .A2(G128), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n797), .A2(new_n1110), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n764), .A2(G137), .B1(new_n766), .B2(G150), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n422), .B1(new_n753), .B2(new_n399), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT120), .Z(new_n1219));
  NAND2_X1  g1019(.A1(new_n752), .A2(G303), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n764), .A2(G283), .B1(new_n766), .B2(G107), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n770), .A2(new_n331), .B1(new_n754), .B2(G77), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1220), .A2(new_n258), .A3(new_n1221), .A4(new_n1222), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n760), .A2(G116), .B1(new_n772), .B2(G97), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n811), .B2(new_n799), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n1217), .A2(new_n1219), .B1(new_n1223), .B2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1211), .B1(new_n1226), .B2(new_n742), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n901), .B2(new_n740), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1210), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1129), .A2(new_n1135), .A3(new_n1132), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1137), .A2(new_n988), .A3(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1230), .A2(new_n1232), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(KEYINPUT121), .ZN(G381));
  NAND3_X1  g1034(.A1(new_n1015), .A2(new_n791), .A3(new_n1049), .ZN(new_n1235));
  OR3_X1    g1035(.A1(G390), .A2(G384), .A3(new_n1235), .ZN(new_n1236));
  NOR3_X1   g1036(.A1(new_n1236), .A2(G387), .A3(G381), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1207), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1100), .A2(new_n1122), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT117), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1100), .A2(KEYINPUT117), .A3(new_n1122), .ZN(new_n1243));
  AND3_X1   g1043(.A1(new_n1239), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1237), .A2(new_n1238), .A3(new_n1244), .ZN(G407));
  NAND2_X1  g1045(.A1(new_n661), .A2(G213), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1238), .A2(new_n1244), .A3(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(G407), .A2(G213), .A3(new_n1248), .ZN(G409));
  AOI21_X1  g1049(.A(new_n791), .B1(new_n1015), .B2(new_n1049), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT125), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1251), .A2(new_n1252), .A3(new_n1235), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1235), .ZN(new_n1254));
  OAI21_X1  g1054(.A(KEYINPUT125), .B1(new_n1254), .B2(new_n1250), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(G390), .A2(new_n1253), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n986), .A2(new_n1076), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT115), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n986), .A2(new_n1076), .A3(KEYINPUT115), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1073), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1255), .A2(new_n1253), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  AND3_X1   g1063(.A1(new_n1256), .A2(new_n1012), .A3(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1012), .B1(new_n1263), .B2(new_n1256), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1238), .A2(G378), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT122), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1177), .A2(new_n1269), .A3(new_n1206), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n990), .B1(new_n1163), .B2(new_n1167), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1206), .ZN(new_n1272));
  OAI21_X1  g1072(.A(KEYINPUT122), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1147), .A2(new_n1168), .A3(new_n988), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1270), .A2(new_n1273), .A3(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1244), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1268), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT62), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1129), .A2(new_n1135), .A3(new_n1132), .A4(KEYINPUT60), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n685), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1137), .A2(KEYINPUT60), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1280), .B1(new_n1281), .B2(new_n1231), .ZN(new_n1282));
  OR2_X1    g1082(.A1(G384), .A2(KEYINPUT123), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  OR3_X1    g1084(.A1(new_n1282), .A2(new_n1284), .A3(new_n1229), .ZN(new_n1285));
  AND2_X1   g1085(.A1(G384), .A2(KEYINPUT123), .ZN(new_n1286));
  OAI22_X1  g1086(.A1(new_n1282), .A2(new_n1229), .B1(new_n1284), .B2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1277), .A2(new_n1278), .A3(new_n1246), .A4(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1247), .A2(G2897), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1285), .A2(new_n1287), .A3(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1291), .B1(new_n1285), .B2(new_n1287), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  AOI22_X1  g1094(.A1(new_n1238), .A2(G378), .B1(new_n1275), .B2(new_n1244), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1294), .B1(new_n1295), .B2(new_n1247), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT61), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1290), .A2(new_n1296), .A3(new_n1297), .ZN(new_n1298));
  XOR2_X1   g1098(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1299));
  NOR2_X1   g1099(.A1(new_n1295), .A2(new_n1247), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1299), .B1(new_n1300), .B2(new_n1289), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1267), .B1(new_n1298), .B2(new_n1301), .ZN(new_n1302));
  XOR2_X1   g1102(.A(KEYINPUT124), .B(KEYINPUT63), .Z(new_n1303));
  NAND2_X1  g1103(.A1(new_n1277), .A2(new_n1246), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1303), .B1(new_n1304), .B2(new_n1288), .ZN(new_n1305));
  AOI21_X1  g1105(.A(KEYINPUT61), .B1(new_n1304), .B2(new_n1294), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1300), .A2(KEYINPUT63), .A3(new_n1289), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1305), .A2(new_n1306), .A3(new_n1266), .A4(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1302), .A2(new_n1308), .ZN(G405));
  AND2_X1   g1109(.A1(new_n1238), .A2(G378), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1125), .A2(new_n1239), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1238), .A2(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(KEYINPUT127), .B1(new_n1310), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT127), .ZN(new_n1314));
  OAI211_X1 g1114(.A(new_n1268), .B(new_n1314), .C1(new_n1238), .C2(new_n1311), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1313), .A2(new_n1289), .A3(new_n1315), .ZN(new_n1316));
  OAI211_X1 g1116(.A(KEYINPUT127), .B(new_n1288), .C1(new_n1310), .C2(new_n1312), .ZN(new_n1317));
  AND3_X1   g1117(.A1(new_n1316), .A2(new_n1266), .A3(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1266), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1318), .A2(new_n1319), .ZN(G402));
endmodule


