//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n851, new_n852, new_n853, new_n854, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975, new_n976;
  INV_X1    g000(.A(KEYINPUT104), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G43gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G71gat), .B(G99gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT27), .B(G183gat), .ZN(new_n206));
  INV_X1    g005(.A(G190gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT28), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  AND2_X1   g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT26), .ZN(new_n214));
  AND3_X1   g013(.A1(new_n213), .A2(KEYINPUT68), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216));
  AOI22_X1  g015(.A1(new_n213), .A2(KEYINPUT68), .B1(new_n216), .B2(new_n214), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n210), .B(new_n212), .C1(new_n215), .C2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n211), .A2(KEYINPUT24), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(G183gat), .B2(G190gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n211), .A2(KEYINPUT24), .ZN(new_n221));
  OR2_X1    g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT25), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT66), .B(KEYINPUT23), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(new_n216), .ZN(new_n225));
  INV_X1    g024(.A(new_n213), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(KEYINPUT65), .B(G169gat), .ZN(new_n228));
  INV_X1    g027(.A(G176gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n228), .A2(KEYINPUT23), .A3(new_n229), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n222), .A2(new_n223), .A3(new_n227), .A4(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n218), .A2(new_n231), .ZN(new_n232));
  NOR3_X1   g031(.A1(new_n211), .A2(KEYINPUT67), .A3(KEYINPUT24), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n220), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT67), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n234), .B1(new_n235), .B2(new_n221), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n213), .A2(KEYINPUT23), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n227), .A2(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n223), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n232), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(G127gat), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n241), .A2(KEYINPUT69), .ZN(new_n242));
  INV_X1    g041(.A(G120gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(G113gat), .ZN(new_n244));
  INV_X1    g043(.A(G113gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(G120gat), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT1), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  MUX2_X1   g046(.A(new_n242), .B(new_n241), .S(new_n247), .Z(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(G134gat), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n240), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n239), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n252), .A2(new_n218), .A3(new_n231), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(new_n249), .ZN(new_n254));
  NAND2_X1  g053(.A1(G227gat), .A2(G233gat), .ZN(new_n255));
  XOR2_X1   g054(.A(new_n255), .B(KEYINPUT64), .Z(new_n256));
  NAND3_X1  g055(.A1(new_n251), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT33), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n205), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(KEYINPUT32), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n257), .B(KEYINPUT32), .C1(new_n258), .C2(new_n205), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n251), .A2(new_n254), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(new_n255), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT34), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n256), .A2(KEYINPUT34), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n263), .B(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(KEYINPUT88), .ZN(new_n271));
  NAND2_X1  g070(.A1(G228gat), .A2(G233gat), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT83), .ZN(new_n273));
  XNOR2_X1  g072(.A(G197gat), .B(G204gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n274), .B(KEYINPUT70), .ZN(new_n275));
  NAND2_X1  g074(.A1(G211gat), .A2(G218gat), .ZN(new_n276));
  INV_X1    g075(.A(G211gat), .ZN(new_n277));
  INV_X1    g076(.A(G218gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT22), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n276), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  OR2_X1    g081(.A1(new_n282), .A2(KEYINPUT71), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n275), .A2(KEYINPUT22), .ZN(new_n284));
  AND2_X1   g083(.A1(new_n279), .A2(new_n276), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n282), .A2(KEYINPUT71), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n283), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT29), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT3), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G148gat), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT76), .B1(new_n291), .B2(G141gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT76), .ZN(new_n293));
  INV_X1    g092(.A(G141gat), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n293), .A2(new_n294), .A3(G148gat), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n292), .B(new_n295), .C1(new_n294), .C2(G148gat), .ZN(new_n296));
  OR2_X1    g095(.A1(new_n296), .A2(KEYINPUT77), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(KEYINPUT77), .ZN(new_n298));
  INV_X1    g097(.A(G155gat), .ZN(new_n299));
  INV_X1    g098(.A(G162gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n299), .A2(new_n300), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n302), .B1(new_n303), .B2(KEYINPUT2), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n297), .A2(new_n298), .A3(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT75), .B(KEYINPUT2), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n291), .A2(G141gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n294), .A2(G148gat), .ZN(new_n308));
  OAI22_X1  g107(.A1(new_n306), .A2(new_n301), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n301), .A2(KEYINPUT74), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n303), .A2(KEYINPUT74), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n302), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n309), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  AND2_X1   g112(.A1(new_n305), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n273), .B1(new_n290), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n305), .A2(new_n313), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n287), .A2(new_n286), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT29), .B1(new_n317), .B2(new_n283), .ZN(new_n318));
  OAI211_X1 g117(.A(KEYINPUT83), .B(new_n316), .C1(new_n318), .C2(KEYINPUT3), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT3), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n314), .A2(KEYINPUT78), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT78), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n323), .B1(new_n316), .B2(KEYINPUT3), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n288), .B1(new_n325), .B2(new_n289), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n272), .B1(new_n320), .B2(new_n326), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n272), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT84), .ZN(new_n329));
  INV_X1    g128(.A(new_n288), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n329), .B1(new_n330), .B2(KEYINPUT29), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n288), .A2(KEYINPUT84), .A3(new_n289), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT3), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n328), .B1(new_n333), .B2(new_n314), .ZN(new_n334));
  INV_X1    g133(.A(G22gat), .ZN(new_n335));
  AND3_X1   g134(.A1(new_n327), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n335), .B1(new_n327), .B2(new_n334), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT85), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n327), .A2(new_n334), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(G22gat), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT85), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n327), .A2(new_n334), .A3(new_n335), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(G78gat), .B(G106gat), .ZN(new_n344));
  INV_X1    g143(.A(G50gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n344), .B(new_n345), .ZN(new_n346));
  XOR2_X1   g145(.A(KEYINPUT82), .B(KEYINPUT31), .Z(new_n347));
  XNOR2_X1  g146(.A(new_n346), .B(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n338), .A2(new_n343), .A3(new_n349), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n340), .A2(new_n341), .A3(new_n348), .A4(new_n342), .ZN(new_n351));
  AND2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT30), .ZN(new_n353));
  NAND2_X1  g152(.A1(G226gat), .A2(G233gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(new_n289), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT72), .B1(new_n232), .B2(new_n239), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT72), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n252), .A2(new_n218), .A3(new_n357), .A4(new_n231), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n355), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n253), .A2(new_n354), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n288), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n356), .A2(new_n358), .A3(G226gat), .A4(G233gat), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n253), .A2(new_n289), .A3(new_n354), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n362), .A2(new_n330), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  XOR2_X1   g164(.A(G8gat), .B(G36gat), .Z(new_n366));
  XNOR2_X1  g165(.A(new_n366), .B(KEYINPUT73), .ZN(new_n367));
  XOR2_X1   g166(.A(G64gat), .B(G92gat), .Z(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n353), .B1(new_n365), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n361), .A2(new_n364), .A3(new_n369), .ZN(new_n372));
  MUX2_X1   g171(.A(new_n353), .B(new_n371), .S(new_n372), .Z(new_n373));
  INV_X1    g172(.A(KEYINPUT35), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n249), .B1(KEYINPUT3), .B2(new_n316), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n325), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n249), .A2(KEYINPUT4), .A3(new_n314), .ZN(new_n378));
  NAND2_X1  g177(.A1(G225gat), .A2(G233gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n249), .A2(new_n314), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT4), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n377), .A2(new_n378), .A3(new_n379), .A4(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT5), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  AND2_X1   g187(.A1(new_n382), .A2(new_n378), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n389), .A2(new_n377), .A3(new_n379), .A4(new_n386), .ZN(new_n390));
  XOR2_X1   g189(.A(G1gat), .B(G29gat), .Z(new_n391));
  XNOR2_X1  g190(.A(G57gat), .B(G85gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n391), .B(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n394));
  XOR2_X1   g193(.A(new_n393), .B(new_n394), .Z(new_n395));
  XNOR2_X1  g194(.A(new_n249), .B(new_n314), .ZN(new_n396));
  INV_X1    g195(.A(new_n379), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(KEYINPUT5), .A3(new_n397), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n388), .A2(new_n390), .A3(new_n395), .A4(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT6), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n388), .A2(new_n390), .A3(new_n398), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT81), .ZN(new_n404));
  INV_X1    g203(.A(new_n395), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n404), .B1(new_n403), .B2(new_n405), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n402), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  OR3_X1    g208(.A1(new_n399), .A2(KEYINPUT86), .A3(new_n400), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT86), .B1(new_n399), .B2(new_n400), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n375), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n271), .A2(new_n352), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n270), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n350), .A2(new_n415), .A3(new_n351), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n383), .A2(new_n387), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n398), .B1(new_n383), .B2(new_n387), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n405), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT81), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n401), .B1(new_n420), .B2(new_n406), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n399), .A2(new_n400), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n373), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(KEYINPUT35), .B1(new_n416), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n414), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n365), .A2(KEYINPUT37), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT87), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(new_n427), .A3(new_n370), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT37), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n429), .B1(new_n361), .B2(new_n364), .ZN(new_n430));
  OAI21_X1  g229(.A(KEYINPUT87), .B1(new_n430), .B2(new_n369), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n361), .A2(new_n429), .A3(new_n364), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n428), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT38), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n330), .B1(new_n359), .B2(new_n360), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n362), .A2(new_n288), .A3(new_n363), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(KEYINPUT37), .A3(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n369), .A2(KEYINPUT38), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n432), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n439), .A2(new_n372), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n409), .A2(new_n412), .A3(new_n434), .A4(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n379), .B1(new_n389), .B2(new_n377), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT39), .B1(new_n396), .B2(new_n397), .ZN(new_n443));
  OR2_X1    g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT39), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n444), .A2(new_n405), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT40), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n372), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT30), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n451), .B1(new_n450), .B2(new_n371), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n444), .A2(KEYINPUT40), .A3(new_n405), .A4(new_n446), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n449), .A2(new_n452), .A3(new_n399), .A4(new_n453), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n441), .A2(new_n351), .A3(new_n350), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n350), .A2(new_n351), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n423), .A2(new_n456), .ZN(new_n457));
  XOR2_X1   g256(.A(new_n270), .B(KEYINPUT36), .Z(new_n458));
  NAND3_X1  g257(.A1(new_n455), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n425), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT17), .ZN(new_n461));
  OR3_X1    g260(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n462), .A2(new_n463), .B1(G29gat), .B2(G36gat), .ZN(new_n464));
  INV_X1    g263(.A(G43gat), .ZN(new_n465));
  AND2_X1   g264(.A1(KEYINPUT91), .A2(G50gat), .ZN(new_n466));
  NOR2_X1   g265(.A1(KEYINPUT91), .A2(G50gat), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n465), .A2(G50gat), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT15), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT15), .B1(new_n345), .B2(G43gat), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n472), .A2(new_n469), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n464), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  OR2_X1    g273(.A1(new_n464), .A2(new_n473), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n461), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n335), .A2(G15gat), .ZN(new_n477));
  INV_X1    g276(.A(G15gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(G22gat), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT16), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n477), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n477), .A2(new_n479), .A3(KEYINPUT94), .ZN(new_n482));
  INV_X1    g281(.A(G1gat), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G15gat), .B(G22gat), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n485), .B(KEYINPUT94), .C1(new_n480), .C2(G1gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(G8gat), .ZN(new_n488));
  INV_X1    g287(.A(G8gat), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n484), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n476), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n464), .A2(new_n473), .ZN(new_n493));
  INV_X1    g292(.A(new_n473), .ZN(new_n494));
  XNOR2_X1  g293(.A(KEYINPUT91), .B(G50gat), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n469), .B1(new_n495), .B2(new_n465), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n494), .B1(new_n496), .B2(KEYINPUT15), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n493), .B1(new_n497), .B2(new_n464), .ZN(new_n498));
  XOR2_X1   g297(.A(KEYINPUT92), .B(KEYINPUT17), .Z(new_n499));
  AOI21_X1  g298(.A(KEYINPUT93), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n474), .A2(new_n475), .A3(KEYINPUT93), .A4(new_n499), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n492), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(G229gat), .A2(G233gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n491), .A2(new_n498), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n503), .A2(KEYINPUT18), .A3(new_n504), .A4(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT95), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n484), .A2(new_n486), .A3(new_n489), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n489), .B1(new_n484), .B2(new_n486), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n474), .A2(new_n475), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n474), .A2(new_n475), .A3(new_n499), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT93), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n501), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n513), .B1(new_n517), .B2(new_n492), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n518), .A2(KEYINPUT95), .A3(KEYINPUT18), .A4(new_n504), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n508), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n511), .A2(new_n512), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(new_n505), .ZN(new_n522));
  XOR2_X1   g321(.A(new_n504), .B(KEYINPUT13), .Z(new_n523));
  AND2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n518), .A2(new_n504), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT18), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  XOR2_X1   g326(.A(G169gat), .B(G197gat), .Z(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(KEYINPUT90), .ZN(new_n529));
  XNOR2_X1  g328(.A(G113gat), .B(G141gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  XOR2_X1   g330(.A(KEYINPUT89), .B(KEYINPUT11), .Z(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT12), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n520), .A2(new_n527), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n535), .B1(new_n520), .B2(new_n527), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  XOR2_X1   g338(.A(G183gat), .B(G211gat), .Z(new_n540));
  XOR2_X1   g339(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n541));
  XNOR2_X1  g340(.A(G127gat), .B(G155gat), .ZN(new_n542));
  INV_X1    g341(.A(G231gat), .ZN(new_n543));
  INV_X1    g342(.A(G233gat), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G71gat), .B(G78gat), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  OR2_X1    g347(.A1(G57gat), .A2(G64gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(G57gat), .A2(G64gat), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT96), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n549), .B(new_n550), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n552), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n548), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  OR2_X1    g355(.A1(new_n551), .A2(new_n552), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n549), .A2(new_n550), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n557), .A2(new_n558), .A3(new_n547), .A4(new_n554), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT21), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n546), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  AOI211_X1 g362(.A(KEYINPUT21), .B(new_n545), .C1(new_n556), .C2(new_n559), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n542), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n542), .ZN(new_n567));
  NOR3_X1   g366(.A1(new_n562), .A2(new_n564), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n541), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n560), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n491), .B1(KEYINPUT21), .B2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n563), .A2(new_n565), .A3(new_n542), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n567), .B1(new_n562), .B2(new_n564), .ZN(new_n574));
  INV_X1    g373(.A(new_n541), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n569), .A2(new_n572), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n572), .B1(new_n569), .B2(new_n576), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n540), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n569), .A2(new_n576), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(new_n571), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n569), .A2(new_n572), .A3(new_n576), .ZN(new_n582));
  INV_X1    g381(.A(new_n540), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(G120gat), .B(G148gat), .Z(new_n586));
  XNOR2_X1  g385(.A(G176gat), .B(G204gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G230gat), .A2(G233gat), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT99), .ZN(new_n590));
  NAND2_X1  g389(.A1(G99gat), .A2(G106gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT8), .ZN(new_n592));
  NAND2_X1  g391(.A1(G85gat), .A2(G92gat), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT7), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(G85gat), .ZN(new_n596));
  INV_X1    g395(.A(G92gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n592), .A2(new_n595), .A3(new_n598), .A4(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT98), .ZN(new_n602));
  INV_X1    g401(.A(new_n591), .ZN(new_n603));
  NOR2_X1   g402(.A1(G99gat), .A2(G106gat), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OR2_X1    g404(.A1(G99gat), .A2(G106gat), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n606), .A2(KEYINPUT98), .A3(new_n591), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n590), .B1(new_n601), .B2(new_n608), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n600), .A2(KEYINPUT99), .A3(new_n605), .A4(new_n607), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n601), .A2(new_n608), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(new_n560), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n601), .A2(new_n608), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n615), .B1(KEYINPUT102), .B2(new_n611), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n605), .A2(new_n607), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n617), .A2(KEYINPUT102), .A3(new_n600), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n570), .B1(new_n616), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(KEYINPUT10), .B1(new_n614), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT10), .ZN(new_n622));
  NOR3_X1   g421(.A1(new_n612), .A2(new_n622), .A3(new_n560), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n589), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n589), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n620), .A2(new_n614), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n588), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n624), .A2(new_n626), .A3(new_n588), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT103), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n624), .A2(KEYINPUT103), .A3(new_n626), .A4(new_n588), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n627), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  XOR2_X1   g431(.A(G134gat), .B(G162gat), .Z(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G190gat), .B(G218gat), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n635), .B(KEYINPUT101), .Z(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT100), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n611), .A2(new_n610), .ZN(new_n639));
  AOI21_X1  g438(.A(KEYINPUT99), .B1(new_n617), .B2(new_n600), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n512), .A2(KEYINPUT17), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n609), .A2(KEYINPUT100), .A3(new_n610), .A4(new_n611), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(new_n517), .ZN(new_n645));
  NAND2_X1  g444(.A1(G232gat), .A2(G233gat), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(KEYINPUT41), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n648), .B1(new_n612), .B2(new_n512), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n637), .B1(new_n645), .B2(new_n650), .ZN(new_n651));
  AOI211_X1 g450(.A(new_n636), .B(new_n649), .C1(new_n644), .C2(new_n517), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n634), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n647), .A2(KEYINPUT41), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT97), .ZN(new_n655));
  INV_X1    g454(.A(new_n517), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n650), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n636), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n645), .A2(new_n637), .A3(new_n650), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n659), .A2(new_n660), .A3(new_n633), .ZN(new_n661));
  AND3_X1   g460(.A1(new_n653), .A2(new_n655), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n655), .B1(new_n653), .B2(new_n661), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n585), .B(new_n632), .C1(new_n662), .C2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  AND4_X1   g464(.A1(new_n202), .A2(new_n460), .A3(new_n539), .A4(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n538), .B1(new_n425), .B2(new_n459), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n202), .B1(new_n667), .B2(new_n665), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n409), .B1(new_n400), .B2(new_n399), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(new_n483), .ZN(G1324gat));
  XOR2_X1   g471(.A(KEYINPUT16), .B(G8gat), .Z(new_n673));
  OAI211_X1 g472(.A(new_n452), .B(new_n673), .C1(new_n666), .C2(new_n668), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n674), .A2(KEYINPUT42), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT42), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n452), .B1(new_n666), .B2(new_n668), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n676), .B1(new_n677), .B2(G8gat), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n675), .B1(new_n674), .B2(new_n678), .ZN(G1325gat));
  OAI21_X1  g478(.A(G15gat), .B1(new_n669), .B2(new_n458), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n271), .A2(new_n478), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n680), .B1(new_n669), .B2(new_n681), .ZN(G1326gat));
  NOR2_X1   g481(.A1(new_n669), .A2(new_n352), .ZN(new_n683));
  XOR2_X1   g482(.A(KEYINPUT43), .B(G22gat), .Z(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(G1327gat));
  OR2_X1    g484(.A1(new_n662), .A2(new_n663), .ZN(new_n686));
  INV_X1    g485(.A(new_n632), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n686), .A2(new_n585), .A3(new_n687), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n667), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(G29gat), .ZN(new_n690));
  INV_X1    g489(.A(new_n670), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT45), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n662), .A2(new_n663), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n694), .A2(KEYINPUT44), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n460), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g495(.A(new_n632), .B(KEYINPUT106), .Z(new_n697));
  INV_X1    g496(.A(new_n585), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT105), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n699), .B1(new_n536), .B2(new_n537), .ZN(new_n700));
  INV_X1    g499(.A(new_n504), .ZN(new_n701));
  AOI211_X1 g500(.A(new_n701), .B(new_n513), .C1(new_n517), .C2(new_n492), .ZN(new_n702));
  AOI21_X1  g501(.A(KEYINPUT95), .B1(new_n702), .B2(KEYINPUT18), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n506), .A2(new_n507), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n527), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n535), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n520), .A2(new_n535), .A3(new_n527), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n707), .A2(KEYINPUT105), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n700), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n697), .A2(new_n698), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n457), .A2(KEYINPUT107), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n423), .A2(new_n456), .A3(new_n714), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n713), .A2(new_n458), .A3(new_n455), .A4(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n686), .B1(new_n716), .B2(new_n425), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n696), .B(new_n712), .C1(new_n717), .C2(KEYINPUT44), .ZN(new_n718));
  OAI21_X1  g517(.A(G29gat), .B1(new_n718), .B2(new_n670), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n693), .A2(new_n719), .ZN(G1328gat));
  INV_X1    g519(.A(G36gat), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n689), .A2(new_n721), .A3(new_n452), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT46), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT108), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n718), .A2(new_n725), .A3(new_n373), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n725), .B1(new_n718), .B2(new_n373), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(G36gat), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n724), .B1(new_n726), .B2(new_n728), .ZN(G1329gat));
  NAND2_X1  g528(.A1(new_n689), .A2(new_n271), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n465), .ZN(new_n731));
  INV_X1    g530(.A(new_n458), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(G43gat), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n731), .B1(new_n718), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(KEYINPUT47), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT47), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n731), .B(new_n736), .C1(new_n718), .C2(new_n733), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n735), .A2(new_n737), .ZN(G1330gat));
  NAND2_X1  g537(.A1(new_n689), .A2(new_n456), .ZN(new_n739));
  INV_X1    g538(.A(new_n495), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n456), .A2(new_n495), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n741), .B1(new_n718), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(KEYINPUT48), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT48), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n741), .B(new_n745), .C1(new_n718), .C2(new_n742), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n746), .ZN(G1331gat));
  NAND3_X1  g546(.A1(new_n455), .A2(new_n458), .A3(new_n715), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n714), .B1(new_n423), .B2(new_n456), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n425), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NOR4_X1   g549(.A1(new_n697), .A2(new_n711), .A3(new_n698), .A4(new_n694), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(new_n670), .ZN(new_n753));
  XOR2_X1   g552(.A(KEYINPUT109), .B(G57gat), .Z(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(G1332gat));
  AOI211_X1 g554(.A(new_n373), .B(new_n752), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n756));
  NOR2_X1   g555(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1333gat));
  NAND2_X1  g557(.A1(new_n732), .A2(G71gat), .ZN(new_n759));
  OR3_X1    g558(.A1(new_n752), .A2(KEYINPUT110), .A3(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(G71gat), .ZN(new_n761));
  INV_X1    g560(.A(new_n271), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n761), .B1(new_n752), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(KEYINPUT110), .B1(new_n752), .B2(new_n759), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n760), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n765), .B(new_n766), .ZN(G1334gat));
  NOR2_X1   g566(.A1(new_n752), .A2(new_n352), .ZN(new_n768));
  XOR2_X1   g567(.A(new_n768), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g568(.A1(new_n711), .A2(new_n585), .ZN(new_n770));
  AND3_X1   g569(.A1(new_n717), .A2(KEYINPUT51), .A3(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(KEYINPUT51), .B1(new_n717), .B2(new_n770), .ZN(new_n772));
  OR2_X1    g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n773), .A2(new_n596), .A3(new_n691), .A4(new_n687), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n711), .A2(new_n585), .A3(new_n632), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n696), .B(new_n775), .C1(new_n717), .C2(KEYINPUT44), .ZN(new_n776));
  OAI21_X1  g575(.A(G85gat), .B1(new_n776), .B2(new_n670), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n774), .A2(new_n777), .ZN(G1336gat));
  NOR3_X1   g577(.A1(new_n697), .A2(new_n373), .A3(G92gat), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n779), .B1(new_n771), .B2(new_n772), .ZN(new_n780));
  OAI21_X1  g579(.A(G92gat), .B1(new_n776), .B2(new_n373), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT52), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n780), .A2(new_n781), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(G1337gat));
  NOR3_X1   g585(.A1(new_n762), .A2(G99gat), .A3(new_n632), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n773), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(G99gat), .B1(new_n776), .B2(new_n458), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(G1338gat));
  NOR3_X1   g589(.A1(new_n352), .A2(G106gat), .A3(new_n697), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n791), .B1(new_n771), .B2(new_n772), .ZN(new_n792));
  OAI21_X1  g591(.A(G106gat), .B1(new_n776), .B2(new_n352), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(KEYINPUT53), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n792), .A2(new_n793), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n795), .A2(new_n797), .ZN(G1339gat));
  INV_X1    g597(.A(new_n615), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n611), .A2(KEYINPUT102), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n560), .B1(new_n801), .B2(new_n618), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n612), .A2(new_n570), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n622), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n623), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n625), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n588), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n804), .A2(new_n805), .A3(new_n625), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n624), .A2(new_n809), .A3(KEYINPUT54), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n808), .A2(new_n810), .A3(KEYINPUT55), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n808), .A2(new_n810), .A3(KEYINPUT113), .A4(KEYINPUT55), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n808), .A2(new_n810), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817));
  AOI22_X1  g616(.A1(new_n816), .A2(new_n817), .B1(new_n630), .B2(new_n631), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n700), .A2(new_n709), .A3(new_n815), .A4(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n533), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n518), .A2(new_n504), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n522), .A2(new_n523), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n708), .A2(new_n823), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n824), .A2(new_n632), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n694), .B1(new_n819), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n815), .A2(new_n818), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n827), .A2(new_n686), .A3(new_n824), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n698), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT112), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n665), .A2(new_n710), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n830), .B1(new_n665), .B2(new_n710), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n670), .A2(new_n452), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n352), .A2(new_n271), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(G113gat), .B1(new_n839), .B2(new_n538), .ZN(new_n840));
  INV_X1    g639(.A(new_n836), .ZN(new_n841));
  INV_X1    g640(.A(new_n416), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n711), .A2(new_n245), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n844), .B(KEYINPUT114), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n840), .B1(new_n843), .B2(new_n845), .ZN(G1340gat));
  OAI21_X1  g645(.A(G120gat), .B1(new_n839), .B2(new_n697), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n632), .A2(G120gat), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n848), .B(KEYINPUT115), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n847), .B1(new_n843), .B2(new_n849), .ZN(G1341gat));
  NOR2_X1   g649(.A1(new_n843), .A2(new_n698), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n851), .A2(KEYINPUT116), .ZN(new_n852));
  AOI21_X1  g651(.A(G127gat), .B1(new_n851), .B2(KEYINPUT116), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n698), .A2(new_n241), .ZN(new_n854));
  AOI22_X1  g653(.A1(new_n852), .A2(new_n853), .B1(new_n838), .B2(new_n854), .ZN(G1342gat));
  XNOR2_X1  g654(.A(KEYINPUT69), .B(G134gat), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n841), .A2(new_n842), .A3(new_n694), .A4(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n857), .A2(KEYINPUT56), .ZN(new_n858));
  XOR2_X1   g657(.A(new_n858), .B(KEYINPUT117), .Z(new_n859));
  NAND2_X1  g658(.A1(new_n838), .A2(new_n694), .ZN(new_n860));
  AOI22_X1  g659(.A1(KEYINPUT56), .A2(new_n857), .B1(new_n860), .B2(G134gat), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(G1343gat));
  NOR3_X1   g661(.A1(new_n836), .A2(new_n352), .A3(new_n732), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n863), .A2(new_n294), .A3(new_n539), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n864), .A2(KEYINPUT58), .ZN(new_n865));
  INV_X1    g664(.A(new_n833), .ZN(new_n866));
  OR3_X1    g665(.A1(new_n827), .A2(new_n686), .A3(new_n824), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n825), .B1(new_n827), .B2(new_n538), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n868), .A2(new_n869), .A3(new_n686), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n869), .B1(new_n868), .B2(new_n686), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n867), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n866), .B1(new_n872), .B2(new_n698), .ZN(new_n873));
  OAI21_X1  g672(.A(KEYINPUT57), .B1(new_n873), .B2(new_n352), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n835), .A2(new_n458), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n352), .B1(new_n829), .B2(new_n833), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n874), .A2(new_n539), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(G141gat), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(KEYINPUT119), .B1(new_n874), .B2(new_n878), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n874), .A2(KEYINPUT119), .A3(new_n878), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n883), .A2(new_n711), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n864), .B1(new_n885), .B2(G141gat), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT58), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n881), .B1(new_n886), .B2(new_n887), .ZN(G1344gat));
  NOR2_X1   g687(.A1(new_n732), .A2(new_n352), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n841), .A2(new_n291), .A3(new_n687), .A4(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n835), .A2(new_n458), .A3(new_n687), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n876), .A2(KEYINPUT57), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT120), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n876), .A2(KEYINPUT120), .A3(KEYINPUT57), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n868), .A2(new_n686), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n867), .ZN(new_n899));
  AOI22_X1  g698(.A1(new_n899), .A2(new_n698), .B1(new_n538), .B2(new_n665), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n877), .B1(new_n900), .B2(new_n352), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n892), .B1(new_n897), .B2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n291), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n828), .B1(new_n686), .B2(new_n868), .ZN(new_n905));
  OAI22_X1  g704(.A1(new_n905), .A2(new_n585), .B1(new_n539), .B2(new_n664), .ZN(new_n906));
  AOI21_X1  g705(.A(KEYINPUT57), .B1(new_n906), .B2(new_n456), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n907), .B1(new_n895), .B2(new_n896), .ZN(new_n908));
  OAI21_X1  g707(.A(KEYINPUT121), .B1(new_n908), .B2(new_n892), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n891), .B1(new_n904), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n891), .A2(G148gat), .ZN(new_n911));
  INV_X1    g710(.A(new_n884), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n912), .A2(new_n882), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n911), .B1(new_n913), .B2(new_n687), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n890), .B1(new_n910), .B2(new_n914), .ZN(G1345gat));
  INV_X1    g714(.A(new_n913), .ZN(new_n916));
  OAI21_X1  g715(.A(G155gat), .B1(new_n916), .B2(new_n698), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n863), .A2(new_n299), .A3(new_n585), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(G1346gat));
  OAI21_X1  g718(.A(G162gat), .B1(new_n916), .B2(new_n686), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n863), .A2(new_n300), .A3(new_n694), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1347gat));
  NOR2_X1   g721(.A1(new_n691), .A2(new_n373), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n834), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n924), .A2(new_n837), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(new_n539), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n924), .A2(new_n416), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n711), .A2(new_n228), .ZN(new_n928));
  AOI22_X1  g727(.A1(new_n926), .A2(G169gat), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT122), .ZN(G1348gat));
  INV_X1    g729(.A(new_n697), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n925), .A2(G176gat), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(G176gat), .B1(new_n927), .B2(new_n687), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT123), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n935), .B1(new_n934), .B2(new_n933), .ZN(G1349gat));
  NAND2_X1  g735(.A1(new_n925), .A2(new_n585), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(G183gat), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n927), .A2(new_n206), .A3(new_n585), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n938), .A2(KEYINPUT124), .A3(new_n939), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g740(.A(new_n207), .B1(new_n925), .B2(new_n694), .ZN(new_n942));
  XOR2_X1   g741(.A(new_n942), .B(KEYINPUT61), .Z(new_n943));
  NAND3_X1  g742(.A1(new_n927), .A2(new_n207), .A3(new_n694), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1351gat));
  NOR3_X1   g744(.A1(new_n924), .A2(new_n352), .A3(new_n732), .ZN(new_n946));
  XOR2_X1   g745(.A(new_n946), .B(KEYINPUT125), .Z(new_n947));
  AOI21_X1  g746(.A(G197gat), .B1(new_n947), .B2(new_n711), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n923), .A2(new_n458), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n908), .A2(new_n949), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n539), .A2(G197gat), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(G1352gat));
  INV_X1    g751(.A(G204gat), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n946), .A2(new_n953), .A3(new_n687), .ZN(new_n954));
  XOR2_X1   g753(.A(new_n954), .B(KEYINPUT62), .Z(new_n955));
  NOR3_X1   g754(.A1(new_n908), .A2(new_n697), .A3(new_n949), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n955), .B1(new_n956), .B2(new_n953), .ZN(G1353gat));
  AND4_X1   g756(.A1(KEYINPUT120), .A2(new_n834), .A3(KEYINPUT57), .A4(new_n456), .ZN(new_n958));
  AOI21_X1  g757(.A(KEYINPUT120), .B1(new_n876), .B2(KEYINPUT57), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n901), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(new_n949), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n960), .A2(new_n585), .A3(new_n961), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n962), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT126), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND4_X1  g764(.A1(new_n962), .A2(KEYINPUT126), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n962), .A2(G211gat), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT63), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n965), .A2(new_n966), .A3(new_n969), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n947), .A2(new_n277), .A3(new_n585), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(G1354gat));
  AND2_X1   g771(.A1(new_n950), .A2(KEYINPUT127), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n694), .B1(new_n950), .B2(KEYINPUT127), .ZN(new_n974));
  OAI21_X1  g773(.A(G218gat), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n947), .A2(new_n278), .A3(new_n694), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(G1355gat));
endmodule


