//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 1 0 0 0 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 0 1 1 0 0 0 0 0 0 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  XNOR2_X1  g0009(.A(KEYINPUT64), .B(G77), .ZN(new_n210));
  INV_X1    g0010(.A(G244), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G50), .A2(G226), .ZN(new_n216));
  NAND4_X1  g0016(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n206), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  AND2_X1   g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G20), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n203), .A2(G50), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n209), .B1(KEYINPUT1), .B2(new_n218), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n222), .B1(KEYINPUT1), .B2(new_n218), .ZN(G361));
  XNOR2_X1  g0023(.A(G250), .B(G257), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT65), .ZN(new_n225));
  XOR2_X1   g0025(.A(G264), .B(G270), .Z(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XOR2_X1   g0029(.A(KEYINPUT2), .B(G226), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n227), .B(new_n231), .Z(G358));
  XNOR2_X1  g0032(.A(G50), .B(G68), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G58), .B(G77), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n233), .B(new_n234), .Z(new_n235));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G351));
  NAND3_X1  g0039(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n240));
  NAND2_X1  g0040(.A1(G1), .A2(G13), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g0042(.A(G20), .ZN(new_n243));
  INV_X1    g0043(.A(G33), .ZN(new_n244));
  NAND3_X1  g0044(.A1(new_n243), .A2(new_n244), .A3(KEYINPUT67), .ZN(new_n245));
  INV_X1    g0045(.A(KEYINPUT67), .ZN(new_n246));
  OAI21_X1  g0046(.A(new_n246), .B1(G20), .B2(G33), .ZN(new_n247));
  AND2_X1   g0047(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G150), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  OAI21_X1  g0050(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT8), .B(G58), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n244), .A2(G20), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n251), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n242), .B1(new_n250), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT68), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n256), .B(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G13), .A3(G20), .ZN(new_n260));
  INV_X1    g0060(.A(G50), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n242), .B1(new_n259), .B2(G20), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n262), .B1(new_n263), .B2(new_n261), .ZN(new_n264));
  XOR2_X1   g0064(.A(new_n264), .B(KEYINPUT69), .Z(new_n265));
  NAND2_X1  g0065(.A1(new_n258), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT3), .B(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(G222), .A2(G1698), .ZN(new_n269));
  INV_X1    g0069(.A(G1698), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(G223), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n268), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n241), .B1(G33), .B2(G41), .ZN(new_n273));
  INV_X1    g0073(.A(new_n210), .ZN(new_n274));
  OAI211_X1 g0074(.A(new_n272), .B(new_n273), .C1(new_n274), .C2(new_n268), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n259), .B1(G41), .B2(G45), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT66), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n219), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT66), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n280), .B(new_n259), .C1(G41), .C2(G45), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n277), .A2(G274), .A3(new_n279), .A4(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G226), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n279), .A2(new_n276), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n275), .B(new_n282), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G169), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n287), .B1(G179), .B2(new_n285), .ZN(new_n288));
  OR2_X1    g0088(.A1(new_n267), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT10), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n266), .A2(KEYINPUT9), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT9), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n258), .A2(new_n265), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n285), .A2(G200), .ZN(new_n295));
  INV_X1    g0095(.A(G190), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n295), .B1(new_n296), .B2(new_n285), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n290), .B1(new_n294), .B2(new_n298), .ZN(new_n299));
  AOI211_X1 g0099(.A(KEYINPUT10), .B(new_n297), .C1(new_n291), .C2(new_n293), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n289), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n268), .A2(G238), .A3(G1698), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n268), .A2(G232), .A3(new_n270), .ZN(new_n303));
  INV_X1    g0103(.A(G107), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n302), .B(new_n303), .C1(new_n304), .C2(new_n268), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n305), .A2(new_n273), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n282), .B1(new_n211), .B2(new_n284), .ZN(new_n307));
  OR2_X1    g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n286), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n263), .A2(G77), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT71), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n310), .B(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n248), .A2(new_n252), .ZN(new_n313));
  XNOR2_X1  g0113(.A(KEYINPUT15), .B(G87), .ZN(new_n314));
  OAI22_X1  g0114(.A1(new_n254), .A2(new_n314), .B1(new_n210), .B2(new_n243), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n242), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n260), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n210), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n318), .B(KEYINPUT70), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n312), .A2(new_n316), .A3(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n306), .A2(new_n307), .ZN(new_n321));
  INV_X1    g0121(.A(G179), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n309), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT72), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n320), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(new_n296), .B2(new_n308), .ZN(new_n327));
  INV_X1    g0127(.A(G200), .ZN(new_n328));
  OAI22_X1  g0128(.A1(new_n320), .A2(new_n325), .B1(new_n321), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n324), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  AND2_X1   g0130(.A1(KEYINPUT3), .A2(G33), .ZN(new_n331));
  NOR2_X1   g0131(.A1(KEYINPUT3), .A2(G33), .ZN(new_n332));
  OAI211_X1 g0132(.A(G226), .B(new_n270), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(G33), .A2(G97), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n268), .A2(G232), .A3(G1698), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n279), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n279), .A2(G238), .A3(new_n276), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n282), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(KEYINPUT13), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n336), .A2(new_n333), .A3(new_n334), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n273), .ZN(new_n342));
  AND2_X1   g0142(.A1(new_n282), .A2(new_n338), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT13), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n340), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n346), .A2(new_n296), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n253), .A2(G77), .B1(G20), .B2(new_n202), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(new_n248), .B2(new_n261), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n242), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT11), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n349), .A2(KEYINPUT11), .A3(new_n242), .ZN(new_n353));
  OR3_X1    g0153(.A1(new_n260), .A2(KEYINPUT12), .A3(G68), .ZN(new_n354));
  OAI21_X1  g0154(.A(KEYINPUT12), .B1(new_n260), .B2(G68), .ZN(new_n355));
  AOI22_X1  g0155(.A1(G68), .A2(new_n263), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n352), .A2(new_n353), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n328), .B1(new_n340), .B2(new_n345), .ZN(new_n358));
  OR3_X1    g0158(.A1(new_n347), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT73), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n357), .B(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT14), .ZN(new_n362));
  NOR3_X1   g0162(.A1(new_n337), .A2(KEYINPUT13), .A3(new_n339), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n344), .B1(new_n342), .B2(new_n343), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n362), .B(G169), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n340), .A2(G179), .A3(new_n345), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n362), .B1(new_n346), .B2(G169), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n361), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n359), .A2(new_n369), .ZN(new_n370));
  NOR3_X1   g0170(.A1(new_n301), .A2(new_n330), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n252), .A2(new_n317), .ZN(new_n372));
  INV_X1    g0172(.A(new_n252), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n259), .A2(G20), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n242), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n260), .ZN(new_n377));
  OAI211_X1 g0177(.A(KEYINPUT76), .B(new_n372), .C1(new_n375), .C2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n317), .A2(new_n242), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n380), .A2(new_n373), .A3(new_n374), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT76), .B1(new_n381), .B2(new_n372), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT75), .ZN(new_n384));
  OAI21_X1  g0184(.A(KEYINPUT7), .B1(new_n268), .B2(G20), .ZN(new_n385));
  INV_X1    g0185(.A(new_n332), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT7), .ZN(new_n387));
  NAND2_X1  g0187(.A1(KEYINPUT3), .A2(G33), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n386), .A2(new_n387), .A3(new_n243), .A4(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n385), .A2(G68), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G58), .A2(G68), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT74), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(KEYINPUT74), .A2(G58), .A3(G68), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n393), .A2(new_n203), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n245), .A2(new_n247), .ZN(new_n396));
  AOI22_X1  g0196(.A1(G20), .A2(new_n395), .B1(new_n396), .B2(G159), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n384), .B1(new_n390), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT16), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n242), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AOI211_X1 g0200(.A(new_n384), .B(KEYINPUT16), .C1(new_n390), .C2(new_n397), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n383), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n279), .A2(G232), .A3(new_n276), .ZN(new_n403));
  AND2_X1   g0203(.A1(new_n282), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G87), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT77), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n405), .B(new_n406), .ZN(new_n407));
  OAI211_X1 g0207(.A(G223), .B(new_n270), .C1(new_n331), .C2(new_n332), .ZN(new_n408));
  OAI211_X1 g0208(.A(G226), .B(G1698), .C1(new_n331), .C2(new_n332), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n273), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT78), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n404), .A2(new_n411), .A3(new_n412), .A4(new_n322), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n404), .A2(new_n411), .A3(new_n322), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT78), .ZN(new_n415));
  AOI21_X1  g0215(.A(G169), .B1(new_n404), .B2(new_n411), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n413), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n402), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT18), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT18), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n402), .A2(new_n417), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT17), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n404), .A2(G190), .A3(new_n411), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n328), .B1(new_n404), .B2(new_n411), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n422), .B1(new_n402), .B2(new_n426), .ZN(new_n427));
  OR2_X1    g0227(.A1(new_n398), .A2(new_n399), .ZN(new_n428));
  INV_X1    g0228(.A(new_n401), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n428), .A2(new_n429), .A3(new_n242), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n430), .A2(KEYINPUT17), .A3(new_n383), .A4(new_n425), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n419), .A2(new_n421), .A3(new_n427), .A4(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  OR2_X1    g0233(.A1(new_n433), .A2(KEYINPUT79), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(KEYINPUT79), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n371), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  OAI211_X1 g0236(.A(G244), .B(new_n270), .C1(new_n331), .C2(new_n332), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT4), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(G250), .A2(G1698), .ZN(new_n440));
  NAND2_X1  g0240(.A1(KEYINPUT4), .A2(G244), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n440), .B1(new_n441), .B2(G1698), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n268), .A2(new_n442), .B1(G33), .B2(G283), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n279), .B1(new_n439), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(G45), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n445), .A2(G1), .ZN(new_n446));
  AND2_X1   g0246(.A1(KEYINPUT5), .A2(G41), .ZN(new_n447));
  NOR2_X1   g0247(.A1(KEYINPUT5), .A2(G41), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(G257), .A3(new_n279), .ZN(new_n450));
  XNOR2_X1  g0250(.A(KEYINPUT5), .B(G41), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n451), .A2(new_n279), .A3(G274), .A4(new_n446), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(G200), .B1(new_n444), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT81), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n444), .A2(new_n453), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G190), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT80), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT6), .ZN(new_n461));
  AND2_X1   g0261(.A1(G97), .A2(G107), .ZN(new_n462));
  NOR2_X1   g0262(.A1(G97), .A2(G107), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n304), .A2(KEYINPUT6), .A3(G97), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n466), .A2(G20), .B1(G77), .B2(new_n396), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n385), .A2(G107), .A3(new_n389), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n376), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n260), .A2(G97), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n259), .A2(G33), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n260), .A2(new_n471), .A3(new_n241), .A4(new_n240), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n470), .B1(new_n473), .B2(G97), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n460), .B1(new_n469), .B2(new_n475), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n385), .A2(G107), .A3(new_n389), .ZN(new_n477));
  AND3_X1   g0277(.A1(new_n304), .A2(KEYINPUT6), .A3(G97), .ZN(new_n478));
  XNOR2_X1  g0278(.A(G97), .B(G107), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n478), .B1(new_n479), .B2(new_n461), .ZN(new_n480));
  INV_X1    g0280(.A(G77), .ZN(new_n481));
  OAI22_X1  g0281(.A1(new_n480), .A2(new_n243), .B1(new_n248), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n242), .B1(new_n477), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n483), .A2(KEYINPUT80), .A3(new_n474), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n457), .A2(new_n455), .A3(G190), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n459), .A2(new_n476), .A3(new_n484), .A4(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n446), .A2(G274), .ZN(new_n487));
  OAI21_X1  g0287(.A(G250), .B1(new_n445), .B2(G1), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n487), .B1(new_n273), .B2(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(G244), .B(G1698), .C1(new_n331), .C2(new_n332), .ZN(new_n490));
  OAI211_X1 g0290(.A(G238), .B(new_n270), .C1(new_n331), .C2(new_n332), .ZN(new_n491));
  XNOR2_X1  g0291(.A(KEYINPUT82), .B(G116), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n490), .B(new_n491), .C1(new_n244), .C2(new_n492), .ZN(new_n493));
  AOI211_X1 g0293(.A(G179), .B(new_n489), .C1(new_n493), .C2(new_n273), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n273), .ZN(new_n495));
  INV_X1    g0295(.A(new_n489), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n494), .B1(new_n286), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT19), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n243), .B1(new_n334), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(G87), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n463), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT83), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n500), .A2(new_n502), .A3(KEYINPUT83), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n268), .A2(new_n243), .A3(G68), .ZN(new_n507));
  INV_X1    g0307(.A(G97), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n499), .B1(new_n254), .B2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n505), .A2(new_n506), .A3(new_n507), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n242), .ZN(new_n511));
  INV_X1    g0311(.A(new_n314), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n512), .A2(new_n260), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n473), .A2(new_n512), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n511), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n495), .A2(new_n496), .A3(new_n296), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n489), .B1(new_n493), .B2(new_n273), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n517), .B1(G200), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n472), .A2(new_n501), .ZN(new_n520));
  AOI211_X1 g0320(.A(new_n513), .B(new_n520), .C1(new_n510), .C2(new_n242), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n498), .A2(new_n516), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n457), .A2(G179), .ZN(new_n523));
  OAI21_X1  g0323(.A(G169), .B1(new_n444), .B2(new_n453), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n483), .A2(new_n474), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n243), .B(G87), .C1(new_n331), .C2(new_n332), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(KEYINPUT22), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT22), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n268), .A2(new_n530), .A3(new_n243), .A4(G87), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT24), .ZN(new_n533));
  OAI21_X1  g0333(.A(KEYINPUT23), .B1(new_n243), .B2(G107), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT23), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n535), .A2(new_n304), .A3(G20), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(G116), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT82), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT82), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(G116), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n244), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n537), .B1(new_n542), .B2(new_n243), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n532), .A2(new_n533), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n533), .B1(new_n532), .B2(new_n543), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n242), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n317), .A2(KEYINPUT25), .A3(new_n304), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT25), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n260), .B2(G107), .ZN(new_n549));
  AOI22_X1  g0349(.A1(G107), .A2(new_n473), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  OAI211_X1 g0350(.A(G257), .B(G1698), .C1(new_n331), .C2(new_n332), .ZN(new_n551));
  OAI211_X1 g0351(.A(G250), .B(new_n270), .C1(new_n331), .C2(new_n332), .ZN(new_n552));
  NAND2_X1  g0352(.A1(G33), .A2(G294), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n273), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n451), .A2(new_n446), .B1(new_n219), .B2(new_n278), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(G264), .ZN(new_n557));
  AND4_X1   g0357(.A1(new_n296), .A2(new_n555), .A3(new_n452), .A4(new_n557), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n554), .A2(new_n273), .B1(new_n556), .B2(G264), .ZN(new_n559));
  AOI21_X1  g0359(.A(G200), .B1(new_n559), .B2(new_n452), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n546), .B(new_n550), .C1(new_n558), .C2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n486), .A2(new_n522), .A3(new_n527), .A4(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n268), .A2(G264), .A3(G1698), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n268), .A2(G257), .A3(new_n270), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n331), .A2(new_n332), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G303), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n273), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n449), .A2(G270), .A3(new_n279), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n569), .A2(KEYINPUT84), .A3(new_n452), .ZN(new_n570));
  AOI21_X1  g0370(.A(KEYINPUT84), .B1(new_n569), .B2(new_n452), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n568), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n539), .A2(new_n541), .ZN(new_n573));
  OAI22_X1  g0373(.A1(new_n472), .A2(new_n538), .B1(new_n260), .B2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(G20), .B1(G33), .B2(G283), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n244), .A2(G97), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n576), .A2(new_n577), .B1(new_n240), .B2(new_n241), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n539), .A2(new_n541), .A3(G20), .ZN(new_n579));
  AOI21_X1  g0379(.A(KEYINPUT20), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n578), .A2(KEYINPUT20), .A3(new_n579), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n575), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n572), .A2(KEYINPUT21), .A3(G169), .A4(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n569), .A2(new_n452), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT84), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n569), .A2(KEYINPUT84), .A3(new_n452), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n588), .A2(G179), .A3(new_n568), .A4(new_n582), .ZN(new_n589));
  AND2_X1   g0389(.A1(new_n583), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n559), .A2(new_n452), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n286), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n559), .A2(new_n322), .A3(new_n452), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n532), .A2(new_n543), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(KEYINPUT24), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n532), .A2(new_n533), .A3(new_n543), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n376), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n550), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n592), .B(new_n593), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT21), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n586), .A2(new_n587), .B1(new_n273), .B2(new_n567), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n581), .A2(new_n580), .ZN(new_n602));
  OAI21_X1  g0402(.A(G169), .B1(new_n602), .B2(new_n574), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n600), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n582), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n568), .B(G190), .C1(new_n570), .C2(new_n571), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n605), .B(new_n606), .C1(new_n601), .C2(new_n328), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n590), .A2(new_n599), .A3(new_n604), .A4(new_n607), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n436), .A2(new_n562), .A3(new_n608), .ZN(G372));
  INV_X1    g0409(.A(new_n436), .ZN(new_n610));
  INV_X1    g0410(.A(new_n494), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n497), .A2(new_n286), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n516), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n592), .A2(new_n593), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n614), .B1(new_n546), .B2(new_n550), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n604), .A2(new_n583), .A3(new_n589), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n613), .B1(new_n562), .B2(new_n617), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n523), .A2(new_n524), .B1(new_n483), .B2(new_n474), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n519), .A2(new_n521), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(new_n620), .A3(new_n613), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(KEYINPUT26), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n484), .A2(new_n476), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n522), .A2(new_n525), .A3(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n622), .B1(new_n624), .B2(KEYINPUT26), .ZN(new_n625));
  OR2_X1    g0425(.A1(new_n618), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n610), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n289), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n402), .A2(new_n417), .A3(new_n420), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n420), .B1(new_n402), .B2(new_n417), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n324), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n359), .A2(new_n632), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n633), .A2(new_n369), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n427), .A2(new_n431), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n631), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n297), .B1(new_n291), .B2(new_n293), .ZN(new_n637));
  XNOR2_X1  g0437(.A(new_n637), .B(new_n290), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n628), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n627), .A2(new_n639), .ZN(G369));
  NAND4_X1  g0440(.A1(new_n607), .A2(new_n604), .A3(new_n583), .A4(new_n589), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n259), .A2(new_n243), .A3(G13), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT27), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n643), .A2(KEYINPUT85), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT85), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n646), .B1(new_n642), .B2(KEYINPUT27), .ZN(new_n647));
  OAI221_X1 g0447(.A(G213), .B1(KEYINPUT27), .B2(new_n642), .C1(new_n645), .C2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(G343), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n651), .A2(new_n605), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n641), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n616), .A2(new_n652), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(KEYINPUT86), .B1(new_n655), .B2(G330), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT86), .ZN(new_n657));
  INV_X1    g0457(.A(G330), .ZN(new_n658));
  AOI211_X1 g0458(.A(new_n657), .B(new_n658), .C1(new_n653), .C2(new_n654), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n561), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n651), .B1(new_n546), .B2(new_n550), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n599), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n615), .A2(new_n651), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n616), .A2(new_n651), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n669), .A2(new_n663), .B1(new_n615), .B2(new_n651), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n667), .A2(new_n670), .ZN(G399));
  NOR2_X1   g0471(.A1(new_n502), .A2(G116), .ZN(new_n672));
  INV_X1    g0472(.A(G41), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n207), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n672), .A2(G1), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n221), .B2(new_n674), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT28), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT90), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT26), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n621), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n522), .A2(KEYINPUT26), .A3(new_n525), .A4(new_n623), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n678), .B1(new_n621), .B2(new_n679), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OAI211_X1 g0484(.A(KEYINPUT29), .B(new_n651), .C1(new_n684), .C2(new_n618), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n626), .A2(new_n651), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  XNOR2_X1  g0487(.A(KEYINPUT89), .B(KEYINPUT29), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n685), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  AND3_X1   g0489(.A1(new_n555), .A2(new_n452), .A3(new_n557), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n322), .B1(new_n444), .B2(new_n453), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n518), .A2(KEYINPUT87), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n518), .A2(KEYINPUT87), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n692), .A2(new_n693), .A3(new_n572), .A4(new_n694), .ZN(new_n695));
  AND3_X1   g0495(.A1(new_n457), .A2(new_n518), .A3(new_n559), .ZN(new_n696));
  OAI211_X1 g0496(.A(new_n568), .B(G179), .C1(new_n570), .C2(new_n571), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n696), .A2(new_n698), .A3(KEYINPUT30), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT30), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n457), .A2(new_n518), .A3(new_n559), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n700), .B1(new_n701), .B2(new_n697), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n695), .A2(new_n699), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT31), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n703), .A2(new_n704), .A3(new_n650), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n704), .B1(new_n703), .B2(new_n650), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT88), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n562), .A2(new_n608), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n708), .B1(new_n709), .B2(new_n651), .ZN(new_n710));
  NOR4_X1   g0510(.A1(new_n562), .A2(new_n608), .A3(KEYINPUT88), .A4(new_n650), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n707), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G330), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n689), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n677), .B1(new_n715), .B2(G1), .ZN(G364));
  INV_X1    g0516(.A(new_n655), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n658), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n718), .A2(KEYINPUT91), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n718), .A2(KEYINPUT91), .ZN(new_n720));
  INV_X1    g0520(.A(G13), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(G20), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n259), .B1(new_n722), .B2(G45), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n674), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n719), .A2(new_n720), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n219), .B1(new_n243), .B2(G169), .ZN(new_n728));
  OR2_X1    g0528(.A1(new_n728), .A2(KEYINPUT92), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(KEYINPUT92), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(G13), .A2(G33), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(G20), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n268), .A2(new_n207), .ZN(new_n737));
  INV_X1    g0537(.A(G355), .ZN(new_n738));
  OAI22_X1  g0538(.A1(new_n737), .A2(new_n738), .B1(G116), .B2(new_n207), .ZN(new_n739));
  OR2_X1    g0539(.A1(new_n235), .A2(new_n445), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n565), .A2(new_n207), .ZN(new_n741));
  INV_X1    g0541(.A(new_n221), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n741), .B1(new_n445), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n739), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n243), .A2(new_n296), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n322), .A2(new_n328), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(G326), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n243), .A2(G190), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n322), .A2(G200), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(G311), .ZN(new_n752));
  OAI22_X1  g0552(.A1(new_n747), .A2(new_n748), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G179), .A2(G200), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G190), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n753), .B1(G294), .B2(new_n756), .ZN(new_n757));
  XOR2_X1   g0557(.A(new_n757), .B(KEYINPUT94), .Z(new_n758));
  NOR2_X1   g0558(.A1(new_n328), .A2(G179), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n745), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n745), .A2(new_n750), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI22_X1  g0563(.A1(G303), .A2(new_n761), .B1(new_n763), .B2(G322), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n746), .A2(new_n749), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  XNOR2_X1  g0566(.A(KEYINPUT33), .B(G317), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n749), .A2(new_n754), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n766), .A2(new_n767), .B1(new_n769), .B2(G329), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n764), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n749), .A2(new_n759), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n268), .B(new_n771), .C1(G283), .C2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n756), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n775), .A2(new_n508), .B1(new_n765), .B2(new_n202), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT93), .ZN(new_n777));
  INV_X1    g0577(.A(new_n751), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n565), .B1(new_n778), .B2(new_n274), .ZN(new_n779));
  INV_X1    g0579(.A(G159), .ZN(new_n780));
  OR3_X1    g0580(.A1(new_n768), .A2(KEYINPUT32), .A3(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(KEYINPUT32), .B1(new_n768), .B2(new_n780), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n779), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n760), .A2(new_n501), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n772), .A2(new_n304), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n747), .A2(new_n261), .B1(new_n762), .B2(new_n201), .ZN(new_n786));
  NOR4_X1   g0586(.A1(new_n783), .A2(new_n784), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n758), .A2(new_n774), .B1(new_n777), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n731), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n726), .B1(new_n736), .B2(new_n744), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT95), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n717), .A2(new_n734), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n727), .A2(new_n660), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(G396));
  NAND2_X1  g0594(.A1(new_n789), .A2(new_n733), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n772), .A2(new_n501), .B1(new_n768), .B2(new_n752), .ZN(new_n796));
  XOR2_X1   g0596(.A(new_n796), .B(KEYINPUT96), .Z(new_n797));
  INV_X1    g0597(.A(G303), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n747), .A2(new_n798), .B1(new_n751), .B2(new_n492), .ZN(new_n799));
  INV_X1    g0599(.A(G283), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n304), .A2(new_n760), .B1(new_n765), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G294), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n565), .B1(new_n762), .B2(new_n802), .C1(new_n775), .C2(new_n508), .ZN(new_n803));
  NOR4_X1   g0603(.A1(new_n797), .A2(new_n799), .A3(new_n801), .A4(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(G137), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n747), .A2(new_n805), .B1(new_n765), .B2(new_n249), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n806), .B(KEYINPUT97), .Z(new_n807));
  INV_X1    g0607(.A(G143), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n807), .B1(new_n808), .B2(new_n762), .C1(new_n780), .C2(new_n751), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT34), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n268), .B1(new_n760), .B2(new_n261), .ZN(new_n811));
  INV_X1    g0611(.A(G132), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n772), .A2(new_n202), .B1(new_n768), .B2(new_n812), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n811), .B(new_n813), .C1(G58), .C2(new_n756), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n804), .B1(new_n810), .B2(new_n814), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n726), .B1(G77), .B2(new_n795), .C1(new_n815), .C2(new_n789), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT98), .Z(new_n817));
  NOR2_X1   g0617(.A1(new_n324), .A2(new_n650), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n320), .A2(new_n650), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n327), .B2(new_n329), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n818), .B1(new_n820), .B2(new_n324), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n817), .B1(new_n733), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n820), .A2(new_n324), .ZN(new_n823));
  INV_X1    g0623(.A(new_n818), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n686), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT99), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n821), .B(new_n651), .C1(new_n618), .C2(new_n625), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n686), .A2(KEYINPUT99), .A3(new_n825), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n829), .A2(new_n713), .A3(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n726), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n713), .B1(new_n829), .B2(new_n830), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n822), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT100), .ZN(G384));
  AOI211_X1 g0636(.A(new_n538), .B(new_n220), .C1(new_n466), .C2(KEYINPUT35), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(KEYINPUT35), .B2(new_n466), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT36), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n274), .A2(G50), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n840), .A2(new_n395), .B1(G50), .B2(new_n202), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n841), .A2(G1), .A3(new_n721), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT101), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n828), .A2(new_n824), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n361), .A2(new_n650), .ZN(new_n846));
  AND3_X1   g0646(.A1(new_n359), .A2(new_n369), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n846), .B1(new_n359), .B2(new_n369), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n845), .A2(new_n850), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n381), .A2(new_n372), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n400), .B2(new_n401), .ZN(new_n853));
  INV_X1    g0653(.A(new_n648), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n432), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n853), .A2(new_n417), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n425), .B(new_n383), .C1(new_n401), .C2(new_n400), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n858), .A2(new_n855), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(KEYINPUT37), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n402), .A2(new_n854), .ZN(new_n862));
  XNOR2_X1  g0662(.A(KEYINPUT102), .B(KEYINPUT37), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n418), .A2(new_n862), .A3(new_n859), .A4(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  AND3_X1   g0665(.A1(new_n857), .A2(new_n865), .A3(KEYINPUT38), .ZN(new_n866));
  AOI21_X1  g0666(.A(KEYINPUT38), .B1(new_n857), .B2(new_n865), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n851), .A2(new_n868), .B1(new_n631), .B2(new_n854), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(KEYINPUT103), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT39), .ZN(new_n871));
  NOR3_X1   g0671(.A1(new_n866), .A2(new_n867), .A3(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT38), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n418), .A2(new_n862), .A3(new_n859), .ZN(new_n874));
  INV_X1    g0674(.A(new_n863), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n876), .A2(new_n864), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n427), .A2(new_n431), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n862), .B1(new_n878), .B2(new_n631), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n873), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n857), .A2(new_n865), .A3(KEYINPUT38), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT39), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n872), .A2(new_n882), .ZN(new_n883));
  OR2_X1    g0683(.A1(new_n369), .A2(new_n650), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n631), .A2(new_n854), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n857), .A2(new_n865), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n873), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n881), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n849), .B1(new_n828), .B2(new_n824), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n887), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT103), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n870), .A2(new_n886), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n639), .B1(new_n689), .B2(new_n436), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n895), .B(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n821), .B1(new_n847), .B2(new_n848), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n484), .A2(new_n476), .A3(new_n485), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n454), .A2(new_n455), .B1(new_n457), .B2(G190), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n527), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n546), .A2(new_n550), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n558), .A2(new_n560), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n613), .B(new_n620), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n641), .A2(new_n615), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n905), .A2(new_n906), .A3(new_n651), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(KEYINPUT88), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n905), .A2(new_n906), .A3(new_n708), .A4(new_n651), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n898), .B1(new_n910), .B2(new_n707), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n890), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT40), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n913), .B1(new_n880), .B2(new_n881), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n912), .A2(new_n913), .B1(new_n914), .B2(new_n911), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n705), .A2(new_n706), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n917), .B1(new_n908), .B2(new_n909), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n916), .B1(new_n436), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n915), .A2(new_n610), .A3(new_n712), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n919), .A2(G330), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n897), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n259), .B2(new_n722), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n897), .A2(new_n921), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n844), .B1(new_n923), .B2(new_n924), .ZN(G367));
  NOR2_X1   g0725(.A1(new_n227), .A2(new_n741), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n735), .B1(new_n207), .B2(new_n314), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n726), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n747), .ZN(new_n929));
  XOR2_X1   g0729(.A(KEYINPUT109), .B(G311), .Z(new_n930));
  AOI22_X1  g0730(.A1(new_n929), .A2(new_n930), .B1(new_n773), .B2(G97), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n931), .B(new_n565), .C1(new_n800), .C2(new_n751), .ZN(new_n932));
  NAND2_X1  g0732(.A1(KEYINPUT46), .A2(G116), .ZN(new_n933));
  XNOR2_X1  g0733(.A(KEYINPUT110), .B(G317), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n760), .A2(new_n933), .B1(new_n768), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n760), .A2(new_n492), .ZN(new_n936));
  OAI22_X1  g0736(.A1(new_n936), .A2(KEYINPUT46), .B1(new_n775), .B2(new_n304), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n802), .A2(new_n765), .B1(new_n762), .B2(new_n798), .ZN(new_n938));
  NOR4_X1   g0738(.A1(new_n932), .A2(new_n935), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n760), .A2(new_n201), .B1(new_n772), .B2(new_n210), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n765), .A2(new_n780), .B1(new_n751), .B2(new_n261), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n929), .A2(G143), .B1(new_n769), .B2(G137), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n756), .A2(G68), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n565), .B1(new_n763), .B2(G150), .ZN(new_n945));
  AND3_X1   g0745(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n939), .B1(new_n942), .B2(new_n946), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n947), .A2(KEYINPUT47), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n789), .B1(new_n947), .B2(KEYINPUT47), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n928), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n651), .A2(new_n521), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(KEYINPUT104), .B1(new_n952), .B2(new_n613), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n522), .B2(new_n952), .ZN(new_n954));
  NOR3_X1   g0754(.A1(new_n952), .A2(KEYINPUT104), .A3(new_n613), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n734), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n950), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n623), .A2(new_n525), .A3(new_n650), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT105), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n623), .A2(new_n650), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n486), .A2(new_n964), .A3(new_n527), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n961), .A2(new_n962), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n963), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  NOR3_X1   g0768(.A1(new_n968), .A2(new_n665), .A3(new_n668), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT42), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n969), .B(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n967), .A2(new_n615), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n650), .B1(new_n972), .B2(new_n527), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n960), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT106), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n667), .B2(new_n968), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n666), .A2(KEYINPUT106), .A3(new_n967), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n974), .A2(new_n976), .ZN(new_n983));
  OR3_X1    g0783(.A1(new_n978), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n982), .B1(new_n978), .B2(new_n983), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n670), .A2(new_n967), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT45), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT44), .ZN(new_n989));
  OR3_X1    g0789(.A1(new_n670), .A2(new_n967), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n989), .B1(new_n670), .B2(new_n967), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n990), .A2(KEYINPUT108), .A3(new_n991), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n991), .A2(KEYINPUT108), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n988), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n994), .A2(new_n666), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n666), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n660), .A2(new_n665), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n668), .B1(new_n667), .B2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n998), .ZN(new_n1000));
  NOR3_X1   g0800(.A1(new_n1000), .A2(new_n666), .A3(new_n669), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n715), .B1(new_n997), .B2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(KEYINPUT107), .B(KEYINPUT41), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n674), .B(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n724), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n959), .B1(new_n986), .B2(new_n1007), .ZN(G387));
  NAND2_X1  g0808(.A1(new_n1002), .A2(new_n714), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n715), .B1(new_n1001), .B2(new_n999), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1009), .A2(new_n725), .A3(new_n1010), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n737), .A2(new_n672), .B1(G107), .B2(new_n207), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n741), .B1(new_n231), .B2(G45), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n445), .B1(new_n202), .B2(new_n481), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT111), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1014), .B1(new_n672), .B2(new_n1015), .ZN(new_n1016));
  AND3_X1   g0816(.A1(new_n373), .A2(KEYINPUT50), .A3(new_n261), .ZN(new_n1017));
  AOI21_X1  g0817(.A(KEYINPUT50), .B1(new_n373), .B2(new_n261), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1016), .B1(new_n1015), .B2(new_n672), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1012), .B1(new_n1013), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n726), .B1(new_n1020), .B2(new_n736), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n760), .A2(new_n210), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n268), .B1(new_n772), .B2(new_n508), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1022), .B(new_n1023), .C1(G159), .C2(new_n929), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G68), .A2(new_n778), .B1(new_n769), .B2(G150), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(G50), .A2(new_n763), .B1(new_n766), .B2(new_n373), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n512), .A2(new_n756), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G322), .A2(new_n929), .B1(new_n766), .B2(new_n930), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n798), .B2(new_n751), .C1(new_n762), .C2(new_n934), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT113), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1031), .A2(KEYINPUT48), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n775), .A2(new_n800), .B1(new_n760), .B2(new_n802), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT112), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n1031), .B2(KEYINPUT48), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1032), .A2(KEYINPUT49), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n268), .B1(new_n769), .B2(G326), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1036), .B(new_n1037), .C1(new_n492), .C2(new_n772), .ZN(new_n1038));
  AOI21_X1  g0838(.A(KEYINPUT49), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1028), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1021), .B1(new_n1040), .B2(new_n731), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n665), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1041), .B1(new_n1042), .B2(new_n958), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT114), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n999), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1001), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1044), .B1(new_n1047), .B2(new_n724), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1011), .A2(new_n1048), .ZN(G393));
  NAND3_X1  g0849(.A1(new_n995), .A2(new_n724), .A3(new_n996), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n747), .A2(new_n249), .B1(new_n762), .B2(new_n780), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT51), .Z(new_n1052));
  OAI22_X1  g0852(.A1(new_n765), .A2(new_n261), .B1(new_n768), .B2(new_n808), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n760), .A2(new_n202), .B1(new_n751), .B2(new_n252), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n756), .A2(G77), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1055), .B(new_n268), .C1(new_n501), .C2(new_n772), .ZN(new_n1056));
  OR4_X1    g0856(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .A4(new_n1056), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G317), .A2(new_n929), .B1(new_n763), .B2(G311), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT52), .Z(new_n1059));
  AOI22_X1  g0859(.A1(G303), .A2(new_n766), .B1(new_n778), .B2(G294), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G283), .A2(new_n761), .B1(new_n769), .B2(G322), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n268), .B(new_n785), .C1(new_n573), .C2(new_n756), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n789), .B1(new_n1057), .B2(new_n1063), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n735), .B1(new_n508), .B2(new_n207), .C1(new_n238), .C2(new_n741), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n832), .B1(new_n1065), .B2(KEYINPUT115), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(KEYINPUT115), .B2(new_n1065), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n967), .B2(new_n958), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1047), .A2(new_n715), .A3(new_n996), .A4(new_n995), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n725), .ZN(new_n1071));
  AND2_X1   g0871(.A1(new_n997), .A2(new_n1010), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1050), .B(new_n1069), .C1(new_n1071), .C2(new_n1072), .ZN(G390));
  OAI22_X1  g0873(.A1(new_n872), .A2(new_n882), .B1(new_n891), .B2(new_n885), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n884), .B(KEYINPUT116), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(new_n881), .B2(new_n880), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n651), .B(new_n823), .C1(new_n684), .C2(new_n618), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n824), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n850), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1076), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n898), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n712), .A2(G330), .A3(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1074), .A2(new_n1080), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n851), .A2(new_n884), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n432), .A2(new_n402), .A3(new_n854), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n876), .A2(new_n864), .ZN(new_n1086));
  AOI21_X1  g0886(.A(KEYINPUT38), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n871), .B1(new_n866), .B2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n889), .A2(KEYINPUT39), .A3(new_n881), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n1084), .A2(new_n1090), .B1(new_n1079), .B2(new_n1076), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT117), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1082), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n911), .A2(KEYINPUT117), .A3(G330), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1083), .B1(new_n1091), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n712), .A2(G330), .A3(new_n821), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT118), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1097), .A2(new_n1098), .A3(new_n849), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1098), .B1(new_n1097), .B2(new_n849), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1082), .A2(new_n824), .A3(new_n1077), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1097), .A2(new_n849), .ZN(new_n1103));
  AOI21_X1  g0903(.A(KEYINPUT117), .B1(new_n911), .B2(G330), .ZN(new_n1104));
  NOR4_X1   g0904(.A1(new_n918), .A2(new_n898), .A3(new_n1092), .A4(new_n658), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1103), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1099), .A2(new_n1102), .B1(new_n1106), .B2(new_n845), .ZN(new_n1107));
  OR2_X1    g0907(.A1(new_n436), .A2(new_n713), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1108), .B(new_n639), .C1(new_n436), .C2(new_n689), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1096), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  NOR3_X1   g0910(.A1(new_n918), .A2(new_n658), .A3(new_n825), .ZN(new_n1111));
  OAI21_X1  g0911(.A(KEYINPUT118), .B1(new_n1111), .B2(new_n850), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1078), .B1(new_n911), .B2(G330), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1112), .A2(new_n1099), .A3(new_n1113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1093), .A2(new_n1094), .B1(new_n849), .B2(new_n1097), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n845), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1114), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1074), .A2(new_n1080), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1118), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1108), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n896), .A2(new_n1120), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1117), .A2(new_n1083), .A3(new_n1119), .A4(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1110), .A2(new_n725), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1096), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1090), .A2(new_n732), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n726), .B1(new_n795), .B2(new_n373), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n765), .A2(new_n805), .ZN(new_n1127));
  INV_X1    g0927(.A(G128), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n268), .B1(new_n747), .B2(new_n1128), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n1127), .B(new_n1129), .C1(G125), .C2(new_n769), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n756), .A2(G159), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n760), .A2(new_n249), .ZN(new_n1132));
  XOR2_X1   g0932(.A(KEYINPUT119), .B(KEYINPUT53), .Z(new_n1133));
  XNOR2_X1  g0933(.A(new_n1132), .B(new_n1133), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n762), .A2(new_n812), .B1(new_n772), .B2(new_n261), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(KEYINPUT54), .B(G143), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1135), .B1(new_n778), .B2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1130), .A2(new_n1131), .A3(new_n1134), .A4(new_n1138), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n202), .A2(new_n772), .B1(new_n751), .B2(new_n508), .ZN(new_n1140));
  NOR3_X1   g0940(.A1(new_n1140), .A2(new_n268), .A3(new_n784), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(G283), .A2(new_n929), .B1(new_n763), .B2(G116), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n766), .A2(G107), .B1(new_n769), .B2(G294), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1141), .A2(new_n1055), .A3(new_n1142), .A4(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1139), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1126), .B1(new_n1145), .B2(new_n731), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1124), .A2(new_n724), .B1(new_n1125), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1123), .A2(new_n1147), .ZN(G378));
  AOI22_X1  g0948(.A1(G125), .A2(new_n929), .B1(new_n761), .B2(new_n1137), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n1128), .B2(new_n762), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n765), .A2(new_n812), .B1(new_n751), .B2(new_n805), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT120), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1151), .B(new_n1153), .C1(new_n249), .C2(new_n775), .ZN(new_n1154));
  OR2_X1    g0954(.A1(new_n1154), .A2(KEYINPUT59), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(KEYINPUT59), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n244), .B(new_n673), .C1(new_n772), .C2(new_n780), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT121), .B(G124), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1157), .B1(new_n769), .B2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1155), .A2(new_n1156), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(G50), .B1(new_n388), .B2(new_n673), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n772), .A2(new_n201), .B1(new_n768), .B2(new_n800), .ZN(new_n1162));
  NOR4_X1   g0962(.A1(new_n1162), .A2(new_n1022), .A3(G41), .A4(new_n268), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(G116), .A2(new_n929), .B1(new_n778), .B2(new_n512), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(G107), .A2(new_n763), .B1(new_n766), .B2(G97), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1163), .A2(new_n944), .A3(new_n1164), .A4(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT58), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1161), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1160), .B(new_n1168), .C1(new_n1167), .C2(new_n1166), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n731), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT122), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1171), .B(new_n726), .C1(G50), .C2(new_n795), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n266), .A2(new_n854), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n638), .B2(new_n289), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n289), .B(new_n1175), .C1(new_n299), .C2(new_n300), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1174), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n301), .A2(new_n266), .A3(new_n854), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1180), .A2(new_n1177), .A3(new_n1173), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1172), .B1(new_n1183), .B2(new_n732), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1182), .B1(new_n915), .B2(G330), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n712), .A2(new_n1081), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n913), .B1(new_n1186), .B2(new_n868), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n914), .A2(new_n911), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1187), .A2(new_n1182), .A3(new_n1188), .A4(G330), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n895), .B1(new_n1185), .B2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1187), .A2(G330), .A3(new_n1188), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(new_n1183), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n883), .A2(new_n885), .B1(new_n892), .B2(new_n893), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1193), .A2(new_n1194), .A3(new_n870), .A4(new_n1189), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1191), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1184), .B1(new_n1196), .B2(new_n724), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1121), .B1(new_n1107), .B2(new_n1096), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1196), .A2(new_n1198), .A3(KEYINPUT57), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(new_n725), .ZN(new_n1200));
  AOI21_X1  g1000(.A(KEYINPUT57), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1197), .B1(new_n1200), .B2(new_n1201), .ZN(G375));
  NAND2_X1  g1002(.A1(new_n849), .A2(new_n732), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n726), .B1(new_n795), .B2(G68), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(G150), .A2(new_n778), .B1(new_n769), .B2(G128), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1205), .B1(new_n805), .B2(new_n762), .C1(new_n780), .C2(new_n760), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(G132), .A2(new_n929), .B1(new_n766), .B2(new_n1137), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n565), .B1(new_n773), .B2(G58), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1207), .B(new_n1208), .C1(new_n261), .C2(new_n775), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n565), .B1(new_n772), .B2(new_n481), .ZN(new_n1210));
  XOR2_X1   g1010(.A(new_n1210), .B(KEYINPUT124), .Z(new_n1211));
  AOI22_X1  g1011(.A1(G294), .A2(new_n929), .B1(new_n763), .B2(G283), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(G97), .A2(new_n761), .B1(new_n766), .B2(new_n573), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G107), .A2(new_n778), .B1(new_n769), .B2(G303), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .A4(new_n1027), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n1206), .A2(new_n1209), .B1(new_n1211), .B2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1204), .B1(new_n1216), .B2(new_n731), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n1117), .A2(new_n724), .B1(new_n1203), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1117), .A2(new_n1121), .ZN(new_n1219));
  XOR2_X1   g1019(.A(new_n1005), .B(KEYINPUT123), .Z(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1117), .A2(new_n1121), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1218), .B1(new_n1221), .B2(new_n1222), .ZN(G381));
  NAND2_X1  g1023(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT57), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1226), .A2(new_n725), .A3(new_n1199), .ZN(new_n1227));
  INV_X1    g1027(.A(G378), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1227), .A2(new_n1228), .A3(new_n1197), .ZN(new_n1229));
  INV_X1    g1029(.A(G390), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(G393), .A2(G396), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT100), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n835), .B(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1230), .A2(new_n1231), .A3(new_n1233), .ZN(new_n1234));
  OR4_X1    g1034(.A1(G387), .A2(new_n1229), .A3(new_n1234), .A4(G381), .ZN(G407));
  OAI211_X1 g1035(.A(G407), .B(G213), .C1(G343), .C2(new_n1229), .ZN(G409));
  NAND2_X1  g1036(.A1(G375), .A2(G378), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1106), .A2(new_n845), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1238), .A2(new_n1109), .A3(KEYINPUT60), .A4(new_n1114), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(new_n725), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1219), .A2(KEYINPUT60), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1222), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1240), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1218), .ZN(new_n1244));
  OAI21_X1  g1044(.A(G384), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1239), .A2(new_n725), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT60), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(new_n1117), .B2(new_n1121), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1246), .B1(new_n1248), .B2(new_n1222), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1249), .A2(new_n1233), .A3(new_n1218), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1245), .A2(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1196), .A2(new_n1198), .A3(new_n1220), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1197), .A2(new_n1252), .A3(new_n1123), .A4(new_n1147), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n649), .A2(G213), .ZN(new_n1254));
  AND2_X1   g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1237), .A2(new_n1251), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(KEYINPUT62), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT62), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1237), .A2(new_n1255), .A3(new_n1258), .A4(new_n1251), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1243), .A2(G384), .A3(new_n1244), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1233), .B1(new_n1249), .B2(new_n1218), .ZN(new_n1261));
  INV_X1    g1061(.A(G2897), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n1260), .A2(new_n1261), .B1(new_n1262), .B2(new_n1254), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1254), .A2(new_n1262), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1245), .A2(new_n1250), .A3(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1228), .B1(new_n1227), .B2(new_n1197), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1263), .B(new_n1265), .C1(new_n1266), .C2(new_n1267), .ZN(new_n1268));
  XOR2_X1   g1068(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n1269));
  NAND4_X1  g1069(.A1(new_n1257), .A2(new_n1259), .A3(new_n1268), .A4(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(G387), .A2(new_n1230), .ZN(new_n1271));
  OAI211_X1 g1071(.A(G390), .B(new_n959), .C1(new_n1007), .C2(new_n986), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n793), .B1(new_n1011), .B2(new_n1048), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1231), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1273), .A2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1271), .A2(new_n1272), .A3(new_n1275), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1270), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1256), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT125), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1245), .A2(new_n1250), .A3(new_n1264), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1264), .B1(new_n1245), .B2(new_n1250), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1282), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1263), .A2(KEYINPUT125), .A3(new_n1265), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1237), .A2(new_n1255), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1285), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1281), .B1(new_n1288), .B2(KEYINPUT63), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1271), .A2(new_n1275), .A3(new_n1272), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1275), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(new_n1290), .A2(new_n1291), .A3(KEYINPUT61), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT63), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1292), .B1(new_n1293), .B2(new_n1256), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1280), .B1(new_n1289), .B2(new_n1294), .ZN(G405));
  INV_X1    g1095(.A(new_n1251), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1296), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1277), .A2(new_n1278), .A3(new_n1251), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1229), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1299), .B1(new_n1300), .B2(new_n1266), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1297), .A2(new_n1298), .A3(new_n1229), .A4(new_n1237), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(G402));
endmodule


