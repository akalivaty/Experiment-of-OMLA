

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U548 ( .A1(n519), .A2(KEYINPUT67), .ZN(n520) );
  XNOR2_X2 U549 ( .A(n523), .B(KEYINPUT64), .ZN(n530) );
  XNOR2_X2 U550 ( .A(n515), .B(n514), .ZN(n534) );
  NOR2_X1 U551 ( .A1(n867), .A2(n728), .ZN(n681) );
  NOR2_X1 U552 ( .A1(n1010), .A2(n695), .ZN(n685) );
  NOR2_X1 U553 ( .A1(n690), .A2(n689), .ZN(n701) );
  INV_X1 U554 ( .A(n728), .ZN(n707) );
  INV_X1 U555 ( .A(KEYINPUT66), .ZN(n513) );
  XNOR2_X1 U556 ( .A(n513), .B(KEYINPUT17), .ZN(n514) );
  NOR2_X1 U557 ( .A1(G651), .A2(G543), .ZN(n636) );
  AND2_X1 U558 ( .A1(G2104), .A2(G2105), .ZN(n981) );
  NOR2_X1 U559 ( .A1(G651), .A2(n630), .ZN(n645) );
  AND2_X1 U560 ( .A1(n528), .A2(n527), .ZN(n678) );
  BUF_X1 U561 ( .A(n678), .Z(G160) );
  NOR2_X1 U562 ( .A1(G2104), .A2(G2105), .ZN(n515) );
  NAND2_X1 U563 ( .A1(G137), .A2(n534), .ZN(n518) );
  NAND2_X1 U564 ( .A1(n981), .A2(G113), .ZN(n516) );
  XOR2_X1 U565 ( .A(KEYINPUT65), .B(n516), .Z(n517) );
  NAND2_X1 U566 ( .A1(n518), .A2(n517), .ZN(n519) );
  NAND2_X1 U567 ( .A1(n519), .A2(KEYINPUT67), .ZN(n521) );
  NAND2_X1 U568 ( .A1(n521), .A2(n520), .ZN(n528) );
  INV_X1 U569 ( .A(G2104), .ZN(n522) );
  AND2_X1 U570 ( .A1(n522), .A2(G2105), .ZN(n980) );
  AND2_X1 U571 ( .A1(G125), .A2(n980), .ZN(n526) );
  NOR2_X1 U572 ( .A1(n522), .A2(G2105), .ZN(n523) );
  NAND2_X1 U573 ( .A1(G101), .A2(n530), .ZN(n524) );
  XNOR2_X1 U574 ( .A(KEYINPUT23), .B(n524), .ZN(n525) );
  NOR2_X1 U575 ( .A1(n526), .A2(n525), .ZN(n527) );
  NAND2_X1 U576 ( .A1(G123), .A2(n980), .ZN(n529) );
  XNOR2_X1 U577 ( .A(n529), .B(KEYINPUT18), .ZN(n539) );
  NAND2_X1 U578 ( .A1(n981), .A2(G111), .ZN(n532) );
  NAND2_X1 U579 ( .A1(G99), .A2(n530), .ZN(n531) );
  NAND2_X1 U580 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U581 ( .A(KEYINPUT78), .B(n533), .ZN(n537) );
  NAND2_X1 U582 ( .A1(G135), .A2(n534), .ZN(n535) );
  XNOR2_X1 U583 ( .A(KEYINPUT77), .B(n535), .ZN(n536) );
  NOR2_X1 U584 ( .A1(n537), .A2(n536), .ZN(n538) );
  NAND2_X1 U585 ( .A1(n539), .A2(n538), .ZN(n1006) );
  XNOR2_X1 U586 ( .A(G2096), .B(n1006), .ZN(n540) );
  OR2_X1 U587 ( .A1(G2100), .A2(n540), .ZN(G156) );
  INV_X1 U588 ( .A(G132), .ZN(G219) );
  INV_X1 U589 ( .A(G82), .ZN(G220) );
  XOR2_X1 U590 ( .A(G543), .B(KEYINPUT0), .Z(n630) );
  NAND2_X1 U591 ( .A1(G52), .A2(n645), .ZN(n543) );
  INV_X1 U592 ( .A(G651), .ZN(n544) );
  NOR2_X1 U593 ( .A1(G543), .A2(n544), .ZN(n541) );
  XOR2_X1 U594 ( .A(KEYINPUT1), .B(n541), .Z(n637) );
  NAND2_X1 U595 ( .A1(G64), .A2(n637), .ZN(n542) );
  NAND2_X1 U596 ( .A1(n543), .A2(n542), .ZN(n549) );
  NAND2_X1 U597 ( .A1(G90), .A2(n636), .ZN(n546) );
  NOR2_X1 U598 ( .A1(n630), .A2(n544), .ZN(n641) );
  NAND2_X1 U599 ( .A1(G77), .A2(n641), .ZN(n545) );
  NAND2_X1 U600 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U601 ( .A(KEYINPUT9), .B(n547), .Z(n548) );
  NOR2_X1 U602 ( .A1(n549), .A2(n548), .ZN(G171) );
  NAND2_X1 U603 ( .A1(n636), .A2(G89), .ZN(n550) );
  XNOR2_X1 U604 ( .A(n550), .B(KEYINPUT4), .ZN(n552) );
  NAND2_X1 U605 ( .A1(G76), .A2(n641), .ZN(n551) );
  NAND2_X1 U606 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U607 ( .A(KEYINPUT5), .B(n553), .ZN(n559) );
  NAND2_X1 U608 ( .A1(n637), .A2(G63), .ZN(n554) );
  XOR2_X1 U609 ( .A(KEYINPUT75), .B(n554), .Z(n556) );
  NAND2_X1 U610 ( .A1(n645), .A2(G51), .ZN(n555) );
  NAND2_X1 U611 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U612 ( .A(KEYINPUT6), .B(n557), .Z(n558) );
  NAND2_X1 U613 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U614 ( .A(KEYINPUT7), .B(n560), .ZN(G168) );
  XOR2_X1 U615 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U616 ( .A1(G94), .A2(G452), .ZN(n561) );
  XOR2_X1 U617 ( .A(KEYINPUT70), .B(n561), .Z(G173) );
  NAND2_X1 U618 ( .A1(G7), .A2(G661), .ZN(n562) );
  XNOR2_X1 U619 ( .A(n562), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U620 ( .A(G223), .ZN(n822) );
  NAND2_X1 U621 ( .A1(n822), .A2(G567), .ZN(n563) );
  XOR2_X1 U622 ( .A(KEYINPUT11), .B(n563), .Z(G234) );
  NAND2_X1 U623 ( .A1(G56), .A2(n637), .ZN(n564) );
  XNOR2_X1 U624 ( .A(n564), .B(KEYINPUT14), .ZN(n567) );
  NAND2_X1 U625 ( .A1(G43), .A2(n645), .ZN(n565) );
  XNOR2_X1 U626 ( .A(n565), .B(KEYINPUT72), .ZN(n566) );
  NAND2_X1 U627 ( .A1(n567), .A2(n566), .ZN(n573) );
  NAND2_X1 U628 ( .A1(n636), .A2(G81), .ZN(n568) );
  XNOR2_X1 U629 ( .A(n568), .B(KEYINPUT12), .ZN(n570) );
  NAND2_X1 U630 ( .A1(G68), .A2(n641), .ZN(n569) );
  NAND2_X1 U631 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U632 ( .A(KEYINPUT13), .B(n571), .Z(n572) );
  NOR2_X1 U633 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U634 ( .A(KEYINPUT73), .B(n574), .ZN(n1013) );
  INV_X1 U635 ( .A(n1013), .ZN(n597) );
  NAND2_X1 U636 ( .A1(G860), .A2(n597), .ZN(n575) );
  XNOR2_X1 U637 ( .A(n575), .B(KEYINPUT74), .ZN(G153) );
  INV_X1 U638 ( .A(G171), .ZN(G301) );
  NAND2_X1 U639 ( .A1(G868), .A2(G301), .ZN(n584) );
  NAND2_X1 U640 ( .A1(G92), .A2(n636), .ZN(n577) );
  NAND2_X1 U641 ( .A1(G79), .A2(n641), .ZN(n576) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n581) );
  NAND2_X1 U643 ( .A1(G54), .A2(n645), .ZN(n579) );
  NAND2_X1 U644 ( .A1(G66), .A2(n637), .ZN(n578) );
  NAND2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(KEYINPUT15), .ZN(n1010) );
  INV_X1 U648 ( .A(G868), .ZN(n596) );
  NAND2_X1 U649 ( .A1(n1010), .A2(n596), .ZN(n583) );
  NAND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(G284) );
  NAND2_X1 U651 ( .A1(G53), .A2(n645), .ZN(n586) );
  NAND2_X1 U652 ( .A1(G65), .A2(n637), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n586), .A2(n585), .ZN(n590) );
  NAND2_X1 U654 ( .A1(G91), .A2(n636), .ZN(n588) );
  NAND2_X1 U655 ( .A1(G78), .A2(n641), .ZN(n587) );
  NAND2_X1 U656 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U657 ( .A1(n590), .A2(n589), .ZN(n897) );
  INV_X1 U658 ( .A(n897), .ZN(G299) );
  NOR2_X1 U659 ( .A1(G286), .A2(n596), .ZN(n592) );
  NOR2_X1 U660 ( .A1(G868), .A2(G299), .ZN(n591) );
  NOR2_X1 U661 ( .A1(n592), .A2(n591), .ZN(G297) );
  INV_X1 U662 ( .A(G860), .ZN(n603) );
  NAND2_X1 U663 ( .A1(n603), .A2(G559), .ZN(n593) );
  INV_X1 U664 ( .A(n1010), .ZN(n601) );
  NAND2_X1 U665 ( .A1(n593), .A2(n601), .ZN(n594) );
  XNOR2_X1 U666 ( .A(n594), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U667 ( .A1(G559), .A2(n1010), .ZN(n595) );
  NOR2_X1 U668 ( .A1(n596), .A2(n595), .ZN(n599) );
  NOR2_X1 U669 ( .A1(n597), .A2(G868), .ZN(n598) );
  NOR2_X1 U670 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U671 ( .A(KEYINPUT76), .B(n600), .Z(G282) );
  NAND2_X1 U672 ( .A1(G559), .A2(n601), .ZN(n602) );
  XOR2_X1 U673 ( .A(n1013), .B(n602), .Z(n654) );
  NAND2_X1 U674 ( .A1(n603), .A2(n654), .ZN(n613) );
  NAND2_X1 U675 ( .A1(n645), .A2(G55), .ZN(n604) );
  XNOR2_X1 U676 ( .A(n604), .B(KEYINPUT80), .ZN(n606) );
  NAND2_X1 U677 ( .A1(G67), .A2(n637), .ZN(n605) );
  NAND2_X1 U678 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U679 ( .A(n607), .B(KEYINPUT81), .ZN(n609) );
  NAND2_X1 U680 ( .A1(G80), .A2(n641), .ZN(n608) );
  NAND2_X1 U681 ( .A1(n609), .A2(n608), .ZN(n612) );
  NAND2_X1 U682 ( .A1(G93), .A2(n636), .ZN(n610) );
  XNOR2_X1 U683 ( .A(KEYINPUT79), .B(n610), .ZN(n611) );
  NOR2_X1 U684 ( .A1(n612), .A2(n611), .ZN(n656) );
  XOR2_X1 U685 ( .A(n613), .B(n656), .Z(G145) );
  NAND2_X1 U686 ( .A1(G88), .A2(n636), .ZN(n614) );
  XNOR2_X1 U687 ( .A(n614), .B(KEYINPUT84), .ZN(n621) );
  NAND2_X1 U688 ( .A1(G50), .A2(n645), .ZN(n616) );
  NAND2_X1 U689 ( .A1(G75), .A2(n641), .ZN(n615) );
  NAND2_X1 U690 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U691 ( .A1(G62), .A2(n637), .ZN(n617) );
  XNOR2_X1 U692 ( .A(KEYINPUT83), .B(n617), .ZN(n618) );
  NOR2_X1 U693 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U694 ( .A1(n621), .A2(n620), .ZN(G303) );
  INV_X1 U695 ( .A(G303), .ZN(G166) );
  NAND2_X1 U696 ( .A1(n636), .A2(G85), .ZN(n622) );
  XNOR2_X1 U697 ( .A(KEYINPUT68), .B(n622), .ZN(n629) );
  NAND2_X1 U698 ( .A1(G47), .A2(n645), .ZN(n624) );
  NAND2_X1 U699 ( .A1(G72), .A2(n641), .ZN(n623) );
  NAND2_X1 U700 ( .A1(n624), .A2(n623), .ZN(n627) );
  NAND2_X1 U701 ( .A1(G60), .A2(n637), .ZN(n625) );
  XNOR2_X1 U702 ( .A(KEYINPUT69), .B(n625), .ZN(n626) );
  NOR2_X1 U703 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U704 ( .A1(n629), .A2(n628), .ZN(G290) );
  NAND2_X1 U705 ( .A1(G49), .A2(n645), .ZN(n632) );
  NAND2_X1 U706 ( .A1(G87), .A2(n630), .ZN(n631) );
  NAND2_X1 U707 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U708 ( .A1(n637), .A2(n633), .ZN(n635) );
  NAND2_X1 U709 ( .A1(G651), .A2(G74), .ZN(n634) );
  NAND2_X1 U710 ( .A1(n635), .A2(n634), .ZN(G288) );
  NAND2_X1 U711 ( .A1(G86), .A2(n636), .ZN(n639) );
  NAND2_X1 U712 ( .A1(G61), .A2(n637), .ZN(n638) );
  NAND2_X1 U713 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U714 ( .A(KEYINPUT82), .B(n640), .ZN(n644) );
  NAND2_X1 U715 ( .A1(n641), .A2(G73), .ZN(n642) );
  XOR2_X1 U716 ( .A(KEYINPUT2), .B(n642), .Z(n643) );
  NOR2_X1 U717 ( .A1(n644), .A2(n643), .ZN(n647) );
  NAND2_X1 U718 ( .A1(n645), .A2(G48), .ZN(n646) );
  NAND2_X1 U719 ( .A1(n647), .A2(n646), .ZN(G305) );
  XNOR2_X1 U720 ( .A(n897), .B(G166), .ZN(n653) );
  XNOR2_X1 U721 ( .A(KEYINPUT19), .B(G290), .ZN(n648) );
  XNOR2_X1 U722 ( .A(n648), .B(G288), .ZN(n649) );
  XNOR2_X1 U723 ( .A(KEYINPUT85), .B(n649), .ZN(n651) );
  XNOR2_X1 U724 ( .A(G305), .B(n656), .ZN(n650) );
  XNOR2_X1 U725 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U726 ( .A(n653), .B(n652), .ZN(n1012) );
  XNOR2_X1 U727 ( .A(n654), .B(n1012), .ZN(n655) );
  NAND2_X1 U728 ( .A1(n655), .A2(G868), .ZN(n658) );
  OR2_X1 U729 ( .A1(G868), .A2(n656), .ZN(n657) );
  NAND2_X1 U730 ( .A1(n658), .A2(n657), .ZN(G295) );
  NAND2_X1 U731 ( .A1(G2084), .A2(G2078), .ZN(n659) );
  XOR2_X1 U732 ( .A(KEYINPUT20), .B(n659), .Z(n660) );
  NAND2_X1 U733 ( .A1(G2090), .A2(n660), .ZN(n662) );
  XNOR2_X1 U734 ( .A(KEYINPUT86), .B(KEYINPUT21), .ZN(n661) );
  XNOR2_X1 U735 ( .A(n662), .B(n661), .ZN(n663) );
  NAND2_X1 U736 ( .A1(G2072), .A2(n663), .ZN(G158) );
  XNOR2_X1 U737 ( .A(KEYINPUT71), .B(G57), .ZN(G237) );
  XNOR2_X1 U738 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U739 ( .A1(G108), .A2(G120), .ZN(n664) );
  NOR2_X1 U740 ( .A1(G237), .A2(n664), .ZN(n665) );
  NAND2_X1 U741 ( .A1(G69), .A2(n665), .ZN(n947) );
  NAND2_X1 U742 ( .A1(n947), .A2(G567), .ZN(n670) );
  NOR2_X1 U743 ( .A1(G220), .A2(G219), .ZN(n666) );
  XOR2_X1 U744 ( .A(KEYINPUT22), .B(n666), .Z(n667) );
  NOR2_X1 U745 ( .A1(G218), .A2(n667), .ZN(n668) );
  NAND2_X1 U746 ( .A1(G96), .A2(n668), .ZN(n948) );
  NAND2_X1 U747 ( .A1(n948), .A2(G2106), .ZN(n669) );
  NAND2_X1 U748 ( .A1(n670), .A2(n669), .ZN(n1023) );
  NAND2_X1 U749 ( .A1(G483), .A2(G661), .ZN(n671) );
  NOR2_X1 U750 ( .A1(n1023), .A2(n671), .ZN(n825) );
  NAND2_X1 U751 ( .A1(n825), .A2(G36), .ZN(G176) );
  NAND2_X1 U752 ( .A1(G102), .A2(n530), .ZN(n673) );
  NAND2_X1 U753 ( .A1(G138), .A2(n534), .ZN(n672) );
  NAND2_X1 U754 ( .A1(n673), .A2(n672), .ZN(n677) );
  NAND2_X1 U755 ( .A1(G126), .A2(n980), .ZN(n675) );
  NAND2_X1 U756 ( .A1(G114), .A2(n981), .ZN(n674) );
  NAND2_X1 U757 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U758 ( .A1(n677), .A2(n676), .ZN(G164) );
  NAND2_X1 U759 ( .A1(G1976), .A2(G288), .ZN(n899) );
  XOR2_X1 U760 ( .A(G1996), .B(KEYINPUT96), .Z(n867) );
  NAND2_X1 U761 ( .A1(n678), .A2(G40), .ZN(n755) );
  INV_X1 U762 ( .A(KEYINPUT92), .ZN(n679) );
  XNOR2_X1 U763 ( .A(n755), .B(n679), .ZN(n680) );
  NOR2_X1 U764 ( .A1(G164), .A2(G1384), .ZN(n756) );
  NAND2_X2 U765 ( .A1(n680), .A2(n756), .ZN(n728) );
  XNOR2_X1 U766 ( .A(n681), .B(KEYINPUT26), .ZN(n682) );
  NOR2_X1 U767 ( .A1(n1013), .A2(n682), .ZN(n684) );
  NAND2_X1 U768 ( .A1(G1341), .A2(n728), .ZN(n683) );
  NAND2_X1 U769 ( .A1(n684), .A2(n683), .ZN(n695) );
  XNOR2_X1 U770 ( .A(n685), .B(KEYINPUT97), .ZN(n693) );
  NOR2_X1 U771 ( .A1(n707), .A2(G1348), .ZN(n687) );
  NOR2_X1 U772 ( .A1(G2067), .A2(n728), .ZN(n686) );
  NOR2_X1 U773 ( .A1(n687), .A2(n686), .ZN(n691) );
  NAND2_X1 U774 ( .A1(n707), .A2(G2072), .ZN(n688) );
  XNOR2_X1 U775 ( .A(n688), .B(KEYINPUT27), .ZN(n690) );
  INV_X1 U776 ( .A(G1956), .ZN(n916) );
  NOR2_X1 U777 ( .A1(n916), .A2(n707), .ZN(n689) );
  NAND2_X1 U778 ( .A1(n897), .A2(n701), .ZN(n694) );
  AND2_X1 U779 ( .A1(n691), .A2(n694), .ZN(n692) );
  NAND2_X1 U780 ( .A1(n693), .A2(n692), .ZN(n699) );
  INV_X1 U781 ( .A(n694), .ZN(n697) );
  NAND2_X1 U782 ( .A1(n1010), .A2(n695), .ZN(n696) );
  OR2_X1 U783 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U784 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U785 ( .A(KEYINPUT98), .B(n700), .ZN(n705) );
  OR2_X1 U786 ( .A1(n701), .A2(n897), .ZN(n702) );
  XNOR2_X1 U787 ( .A(n702), .B(KEYINPUT28), .ZN(n703) );
  XNOR2_X1 U788 ( .A(n703), .B(KEYINPUT95), .ZN(n704) );
  NOR2_X1 U789 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U790 ( .A(n706), .B(KEYINPUT29), .ZN(n712) );
  INV_X1 U791 ( .A(G1961), .ZN(n894) );
  NAND2_X1 U792 ( .A1(n728), .A2(n894), .ZN(n709) );
  XNOR2_X1 U793 ( .A(G2078), .B(KEYINPUT25), .ZN(n877) );
  NAND2_X1 U794 ( .A1(n707), .A2(n877), .ZN(n708) );
  NAND2_X1 U795 ( .A1(n709), .A2(n708), .ZN(n717) );
  AND2_X1 U796 ( .A1(n717), .A2(G171), .ZN(n710) );
  XOR2_X1 U797 ( .A(KEYINPUT94), .B(n710), .Z(n711) );
  NAND2_X1 U798 ( .A1(n712), .A2(n711), .ZN(n736) );
  NAND2_X1 U799 ( .A1(G8), .A2(n728), .ZN(n797) );
  NOR2_X1 U800 ( .A1(G1966), .A2(n797), .ZN(n725) );
  NOR2_X1 U801 ( .A1(n728), .A2(G2084), .ZN(n713) );
  XNOR2_X1 U802 ( .A(n713), .B(KEYINPUT93), .ZN(n722) );
  NAND2_X1 U803 ( .A1(G8), .A2(n722), .ZN(n714) );
  NOR2_X1 U804 ( .A1(n725), .A2(n714), .ZN(n715) );
  XOR2_X1 U805 ( .A(KEYINPUT30), .B(n715), .Z(n716) );
  NOR2_X1 U806 ( .A1(G168), .A2(n716), .ZN(n719) );
  NOR2_X1 U807 ( .A1(G171), .A2(n717), .ZN(n718) );
  NOR2_X1 U808 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U809 ( .A(KEYINPUT31), .B(n720), .Z(n734) );
  NAND2_X1 U810 ( .A1(n736), .A2(n734), .ZN(n721) );
  XNOR2_X1 U811 ( .A(n721), .B(KEYINPUT99), .ZN(n727) );
  INV_X1 U812 ( .A(n722), .ZN(n723) );
  AND2_X1 U813 ( .A1(G8), .A2(n723), .ZN(n724) );
  OR2_X1 U814 ( .A1(n725), .A2(n724), .ZN(n726) );
  OR2_X1 U815 ( .A1(n727), .A2(n726), .ZN(n744) );
  NOR2_X1 U816 ( .A1(G1971), .A2(n797), .ZN(n730) );
  NOR2_X1 U817 ( .A1(G2090), .A2(n728), .ZN(n729) );
  NOR2_X1 U818 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U819 ( .A(KEYINPUT100), .B(n731), .Z(n732) );
  NOR2_X1 U820 ( .A1(G166), .A2(n732), .ZN(n733) );
  XNOR2_X1 U821 ( .A(n733), .B(KEYINPUT101), .ZN(n737) );
  AND2_X1 U822 ( .A1(n734), .A2(n737), .ZN(n735) );
  NAND2_X1 U823 ( .A1(n736), .A2(n735), .ZN(n741) );
  INV_X1 U824 ( .A(n737), .ZN(n738) );
  OR2_X1 U825 ( .A1(n738), .A2(G286), .ZN(n739) );
  AND2_X1 U826 ( .A1(n739), .A2(G8), .ZN(n740) );
  NAND2_X1 U827 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U828 ( .A(KEYINPUT32), .B(n742), .ZN(n743) );
  NAND2_X1 U829 ( .A1(n744), .A2(n743), .ZN(n792) );
  NOR2_X1 U830 ( .A1(G1976), .A2(G288), .ZN(n898) );
  NOR2_X1 U831 ( .A1(G1971), .A2(G303), .ZN(n745) );
  NOR2_X1 U832 ( .A1(n898), .A2(n745), .ZN(n746) );
  NAND2_X1 U833 ( .A1(n792), .A2(n746), .ZN(n747) );
  NAND2_X1 U834 ( .A1(n899), .A2(n747), .ZN(n748) );
  NOR2_X1 U835 ( .A1(KEYINPUT33), .A2(n748), .ZN(n749) );
  INV_X1 U836 ( .A(n797), .ZN(n750) );
  NAND2_X1 U837 ( .A1(n749), .A2(n750), .ZN(n753) );
  NAND2_X1 U838 ( .A1(n898), .A2(n750), .ZN(n751) );
  NAND2_X1 U839 ( .A1(n751), .A2(KEYINPUT33), .ZN(n752) );
  NAND2_X1 U840 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U841 ( .A(KEYINPUT102), .B(n754), .ZN(n788) );
  XOR2_X1 U842 ( .A(G1981), .B(G305), .Z(n891) );
  NOR2_X1 U843 ( .A1(n756), .A2(n755), .ZN(n817) );
  NAND2_X1 U844 ( .A1(G104), .A2(n530), .ZN(n757) );
  XOR2_X1 U845 ( .A(KEYINPUT87), .B(n757), .Z(n759) );
  NAND2_X1 U846 ( .A1(G140), .A2(n534), .ZN(n758) );
  NAND2_X1 U847 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U848 ( .A(KEYINPUT34), .B(n760), .ZN(n765) );
  NAND2_X1 U849 ( .A1(G128), .A2(n980), .ZN(n762) );
  NAND2_X1 U850 ( .A1(G116), .A2(n981), .ZN(n761) );
  NAND2_X1 U851 ( .A1(n762), .A2(n761), .ZN(n763) );
  XOR2_X1 U852 ( .A(KEYINPUT35), .B(n763), .Z(n764) );
  NOR2_X1 U853 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U854 ( .A(KEYINPUT36), .B(n766), .ZN(n1007) );
  XNOR2_X1 U855 ( .A(G2067), .B(KEYINPUT37), .ZN(n815) );
  NOR2_X1 U856 ( .A1(n1007), .A2(n815), .ZN(n844) );
  NAND2_X1 U857 ( .A1(n817), .A2(n844), .ZN(n813) );
  NAND2_X1 U858 ( .A1(n530), .A2(G105), .ZN(n767) );
  XNOR2_X1 U859 ( .A(n767), .B(KEYINPUT38), .ZN(n774) );
  NAND2_X1 U860 ( .A1(n981), .A2(G117), .ZN(n769) );
  NAND2_X1 U861 ( .A1(G141), .A2(n534), .ZN(n768) );
  NAND2_X1 U862 ( .A1(n769), .A2(n768), .ZN(n772) );
  NAND2_X1 U863 ( .A1(G129), .A2(n980), .ZN(n770) );
  XNOR2_X1 U864 ( .A(KEYINPUT89), .B(n770), .ZN(n771) );
  NOR2_X1 U865 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U866 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U867 ( .A(KEYINPUT90), .B(n775), .ZN(n1000) );
  NAND2_X1 U868 ( .A1(G1996), .A2(n1000), .ZN(n783) );
  XNOR2_X1 U869 ( .A(G1991), .B(KEYINPUT88), .ZN(n872) );
  NAND2_X1 U870 ( .A1(G119), .A2(n980), .ZN(n777) );
  NAND2_X1 U871 ( .A1(G107), .A2(n981), .ZN(n776) );
  NAND2_X1 U872 ( .A1(n777), .A2(n776), .ZN(n781) );
  NAND2_X1 U873 ( .A1(G95), .A2(n530), .ZN(n779) );
  NAND2_X1 U874 ( .A1(G131), .A2(n534), .ZN(n778) );
  NAND2_X1 U875 ( .A1(n779), .A2(n778), .ZN(n780) );
  OR2_X1 U876 ( .A1(n781), .A2(n780), .ZN(n997) );
  NAND2_X1 U877 ( .A1(n872), .A2(n997), .ZN(n782) );
  NAND2_X1 U878 ( .A1(n783), .A2(n782), .ZN(n840) );
  NAND2_X1 U879 ( .A1(n840), .A2(n817), .ZN(n784) );
  XNOR2_X1 U880 ( .A(n784), .B(KEYINPUT91), .ZN(n809) );
  INV_X1 U881 ( .A(n809), .ZN(n785) );
  NAND2_X1 U882 ( .A1(n813), .A2(n785), .ZN(n801) );
  INV_X1 U883 ( .A(n801), .ZN(n786) );
  AND2_X1 U884 ( .A1(n891), .A2(n786), .ZN(n787) );
  NAND2_X1 U885 ( .A1(n788), .A2(n787), .ZN(n803) );
  NOR2_X1 U886 ( .A1(G2090), .A2(G303), .ZN(n789) );
  XOR2_X1 U887 ( .A(KEYINPUT103), .B(n789), .Z(n790) );
  NAND2_X1 U888 ( .A1(G8), .A2(n790), .ZN(n791) );
  NAND2_X1 U889 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U890 ( .A(n793), .B(KEYINPUT104), .ZN(n794) );
  NAND2_X1 U891 ( .A1(n794), .A2(n797), .ZN(n799) );
  NOR2_X1 U892 ( .A1(G1981), .A2(G305), .ZN(n795) );
  XOR2_X1 U893 ( .A(n795), .B(KEYINPUT24), .Z(n796) );
  OR2_X1 U894 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U895 ( .A1(n799), .A2(n798), .ZN(n800) );
  OR2_X1 U896 ( .A1(n801), .A2(n800), .ZN(n802) );
  NAND2_X1 U897 ( .A1(n803), .A2(n802), .ZN(n805) );
  XNOR2_X1 U898 ( .A(G1986), .B(G290), .ZN(n902) );
  NAND2_X1 U899 ( .A1(n902), .A2(n817), .ZN(n804) );
  NAND2_X1 U900 ( .A1(n805), .A2(n804), .ZN(n820) );
  NOR2_X1 U901 ( .A1(G1996), .A2(n1000), .ZN(n806) );
  XOR2_X1 U902 ( .A(KEYINPUT105), .B(n806), .Z(n834) );
  NOR2_X1 U903 ( .A1(n997), .A2(n872), .ZN(n837) );
  NOR2_X1 U904 ( .A1(G1986), .A2(G290), .ZN(n807) );
  NOR2_X1 U905 ( .A1(n837), .A2(n807), .ZN(n808) );
  NOR2_X1 U906 ( .A1(n809), .A2(n808), .ZN(n810) );
  XNOR2_X1 U907 ( .A(n810), .B(KEYINPUT106), .ZN(n811) );
  NOR2_X1 U908 ( .A1(n834), .A2(n811), .ZN(n812) );
  XNOR2_X1 U909 ( .A(n812), .B(KEYINPUT39), .ZN(n814) );
  NAND2_X1 U910 ( .A1(n814), .A2(n813), .ZN(n816) );
  NAND2_X1 U911 ( .A1(n1007), .A2(n815), .ZN(n846) );
  NAND2_X1 U912 ( .A1(n816), .A2(n846), .ZN(n818) );
  NAND2_X1 U913 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U914 ( .A1(n820), .A2(n819), .ZN(n821) );
  XNOR2_X1 U915 ( .A(KEYINPUT40), .B(n821), .ZN(G329) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n822), .ZN(G217) );
  AND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n823) );
  NAND2_X1 U918 ( .A1(G661), .A2(n823), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n824) );
  NAND2_X1 U920 ( .A1(n825), .A2(n824), .ZN(G188) );
  NAND2_X1 U922 ( .A1(n980), .A2(G124), .ZN(n826) );
  XNOR2_X1 U923 ( .A(n826), .B(KEYINPUT44), .ZN(n828) );
  NAND2_X1 U924 ( .A1(G112), .A2(n981), .ZN(n827) );
  NAND2_X1 U925 ( .A1(n828), .A2(n827), .ZN(n832) );
  NAND2_X1 U926 ( .A1(G100), .A2(n530), .ZN(n830) );
  NAND2_X1 U927 ( .A1(G136), .A2(n534), .ZN(n829) );
  NAND2_X1 U928 ( .A1(n830), .A2(n829), .ZN(n831) );
  NOR2_X1 U929 ( .A1(n832), .A2(n831), .ZN(G162) );
  XOR2_X1 U930 ( .A(G2090), .B(G162), .Z(n833) );
  NOR2_X1 U931 ( .A1(n834), .A2(n833), .ZN(n835) );
  XOR2_X1 U932 ( .A(KEYINPUT51), .B(n835), .Z(n842) );
  XOR2_X1 U933 ( .A(G160), .B(G2084), .Z(n836) );
  NOR2_X1 U934 ( .A1(n837), .A2(n836), .ZN(n838) );
  NAND2_X1 U935 ( .A1(n838), .A2(n1006), .ZN(n839) );
  NOR2_X1 U936 ( .A1(n840), .A2(n839), .ZN(n841) );
  NAND2_X1 U937 ( .A1(n842), .A2(n841), .ZN(n843) );
  NOR2_X1 U938 ( .A1(n844), .A2(n843), .ZN(n845) );
  XNOR2_X1 U939 ( .A(n845), .B(KEYINPUT120), .ZN(n847) );
  NAND2_X1 U940 ( .A1(n847), .A2(n846), .ZN(n862) );
  NAND2_X1 U941 ( .A1(G103), .A2(n530), .ZN(n848) );
  XNOR2_X1 U942 ( .A(KEYINPUT115), .B(n848), .ZN(n856) );
  NAND2_X1 U943 ( .A1(G127), .A2(n980), .ZN(n850) );
  NAND2_X1 U944 ( .A1(G115), .A2(n981), .ZN(n849) );
  NAND2_X1 U945 ( .A1(n850), .A2(n849), .ZN(n851) );
  XNOR2_X1 U946 ( .A(n851), .B(KEYINPUT116), .ZN(n852) );
  XNOR2_X1 U947 ( .A(n852), .B(KEYINPUT47), .ZN(n854) );
  NAND2_X1 U948 ( .A1(G139), .A2(n534), .ZN(n853) );
  NAND2_X1 U949 ( .A1(n854), .A2(n853), .ZN(n855) );
  NOR2_X1 U950 ( .A1(n856), .A2(n855), .ZN(n993) );
  XNOR2_X1 U951 ( .A(G2072), .B(n993), .ZN(n858) );
  XNOR2_X1 U952 ( .A(G164), .B(G2078), .ZN(n857) );
  NAND2_X1 U953 ( .A1(n858), .A2(n857), .ZN(n859) );
  XOR2_X1 U954 ( .A(KEYINPUT121), .B(n859), .Z(n860) );
  XNOR2_X1 U955 ( .A(KEYINPUT50), .B(n860), .ZN(n861) );
  NOR2_X1 U956 ( .A1(n862), .A2(n861), .ZN(n863) );
  XNOR2_X1 U957 ( .A(KEYINPUT52), .B(n863), .ZN(n865) );
  INV_X1 U958 ( .A(KEYINPUT55), .ZN(n864) );
  NAND2_X1 U959 ( .A1(n865), .A2(n864), .ZN(n866) );
  NAND2_X1 U960 ( .A1(n866), .A2(G29), .ZN(n945) );
  XOR2_X1 U961 ( .A(G29), .B(KEYINPUT124), .Z(n889) );
  XNOR2_X1 U962 ( .A(G32), .B(n867), .ZN(n868) );
  XNOR2_X1 U963 ( .A(n868), .B(KEYINPUT122), .ZN(n876) );
  XNOR2_X1 U964 ( .A(G2067), .B(G26), .ZN(n870) );
  XNOR2_X1 U965 ( .A(G33), .B(G2072), .ZN(n869) );
  NOR2_X1 U966 ( .A1(n870), .A2(n869), .ZN(n871) );
  NAND2_X1 U967 ( .A1(G28), .A2(n871), .ZN(n874) );
  XNOR2_X1 U968 ( .A(G25), .B(n872), .ZN(n873) );
  NOR2_X1 U969 ( .A1(n874), .A2(n873), .ZN(n875) );
  NAND2_X1 U970 ( .A1(n876), .A2(n875), .ZN(n879) );
  XOR2_X1 U971 ( .A(G27), .B(n877), .Z(n878) );
  NOR2_X1 U972 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U973 ( .A(KEYINPUT53), .B(n880), .Z(n884) );
  XNOR2_X1 U974 ( .A(KEYINPUT54), .B(G34), .ZN(n881) );
  XNOR2_X1 U975 ( .A(n881), .B(KEYINPUT123), .ZN(n882) );
  XNOR2_X1 U976 ( .A(G2084), .B(n882), .ZN(n883) );
  NAND2_X1 U977 ( .A1(n884), .A2(n883), .ZN(n886) );
  XNOR2_X1 U978 ( .A(G35), .B(G2090), .ZN(n885) );
  NOR2_X1 U979 ( .A1(n886), .A2(n885), .ZN(n887) );
  XNOR2_X1 U980 ( .A(n887), .B(KEYINPUT55), .ZN(n888) );
  NAND2_X1 U981 ( .A1(n889), .A2(n888), .ZN(n890) );
  NAND2_X1 U982 ( .A1(G11), .A2(n890), .ZN(n943) );
  XNOR2_X1 U983 ( .A(G16), .B(KEYINPUT56), .ZN(n915) );
  XNOR2_X1 U984 ( .A(G1966), .B(G168), .ZN(n892) );
  NAND2_X1 U985 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U986 ( .A(n893), .B(KEYINPUT57), .ZN(n913) );
  XNOR2_X1 U987 ( .A(G171), .B(n894), .ZN(n896) );
  XNOR2_X1 U988 ( .A(G1348), .B(n1010), .ZN(n895) );
  NOR2_X1 U989 ( .A1(n896), .A2(n895), .ZN(n909) );
  XNOR2_X1 U990 ( .A(n897), .B(G1956), .ZN(n904) );
  INV_X1 U991 ( .A(n898), .ZN(n900) );
  NAND2_X1 U992 ( .A1(n900), .A2(n899), .ZN(n901) );
  NOR2_X1 U993 ( .A1(n902), .A2(n901), .ZN(n903) );
  NAND2_X1 U994 ( .A1(n904), .A2(n903), .ZN(n907) );
  XOR2_X1 U995 ( .A(G1971), .B(G303), .Z(n905) );
  XNOR2_X1 U996 ( .A(KEYINPUT125), .B(n905), .ZN(n906) );
  NOR2_X1 U997 ( .A1(n907), .A2(n906), .ZN(n908) );
  NAND2_X1 U998 ( .A1(n909), .A2(n908), .ZN(n911) );
  XNOR2_X1 U999 ( .A(G1341), .B(n1013), .ZN(n910) );
  NOR2_X1 U1000 ( .A1(n911), .A2(n910), .ZN(n912) );
  NAND2_X1 U1001 ( .A1(n913), .A2(n912), .ZN(n914) );
  NAND2_X1 U1002 ( .A1(n915), .A2(n914), .ZN(n941) );
  INV_X1 U1003 ( .A(G16), .ZN(n939) );
  XNOR2_X1 U1004 ( .A(G20), .B(n916), .ZN(n920) );
  XNOR2_X1 U1005 ( .A(G1341), .B(G19), .ZN(n918) );
  XNOR2_X1 U1006 ( .A(G6), .B(G1981), .ZN(n917) );
  NOR2_X1 U1007 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1008 ( .A1(n920), .A2(n919), .ZN(n923) );
  XOR2_X1 U1009 ( .A(KEYINPUT59), .B(G1348), .Z(n921) );
  XNOR2_X1 U1010 ( .A(G4), .B(n921), .ZN(n922) );
  NOR2_X1 U1011 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1012 ( .A(KEYINPUT60), .B(n924), .ZN(n934) );
  XNOR2_X1 U1013 ( .A(G1966), .B(KEYINPUT126), .ZN(n925) );
  XNOR2_X1 U1014 ( .A(n925), .B(G21), .ZN(n932) );
  XNOR2_X1 U1015 ( .A(G1971), .B(G22), .ZN(n927) );
  XNOR2_X1 U1016 ( .A(G23), .B(G1976), .ZN(n926) );
  NOR2_X1 U1017 ( .A1(n927), .A2(n926), .ZN(n929) );
  XOR2_X1 U1018 ( .A(G1986), .B(G24), .Z(n928) );
  NAND2_X1 U1019 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1020 ( .A(KEYINPUT58), .B(n930), .ZN(n931) );
  NOR2_X1 U1021 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1022 ( .A1(n934), .A2(n933), .ZN(n936) );
  XNOR2_X1 U1023 ( .A(G5), .B(G1961), .ZN(n935) );
  NOR2_X1 U1024 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1025 ( .A(KEYINPUT61), .B(n937), .ZN(n938) );
  NAND2_X1 U1026 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1027 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1028 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1029 ( .A1(n945), .A2(n944), .ZN(n946) );
  XOR2_X1 U1030 ( .A(KEYINPUT62), .B(n946), .Z(G311) );
  XNOR2_X1 U1031 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1032 ( .A(G120), .ZN(G236) );
  INV_X1 U1033 ( .A(G108), .ZN(G238) );
  INV_X1 U1034 ( .A(G96), .ZN(G221) );
  INV_X1 U1035 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1036 ( .A1(n948), .A2(n947), .ZN(G325) );
  INV_X1 U1037 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U1038 ( .A(G1341), .B(G2454), .ZN(n949) );
  XNOR2_X1 U1039 ( .A(n949), .B(G2430), .ZN(n950) );
  XNOR2_X1 U1040 ( .A(n950), .B(G1348), .ZN(n956) );
  XOR2_X1 U1041 ( .A(G2443), .B(G2427), .Z(n952) );
  XNOR2_X1 U1042 ( .A(G2438), .B(G2446), .ZN(n951) );
  XNOR2_X1 U1043 ( .A(n952), .B(n951), .ZN(n954) );
  XOR2_X1 U1044 ( .A(G2451), .B(G2435), .Z(n953) );
  XNOR2_X1 U1045 ( .A(n954), .B(n953), .ZN(n955) );
  XNOR2_X1 U1046 ( .A(n956), .B(n955), .ZN(n957) );
  NAND2_X1 U1047 ( .A1(n957), .A2(G14), .ZN(n958) );
  XNOR2_X1 U1048 ( .A(KEYINPUT107), .B(n958), .ZN(G401) );
  XOR2_X1 U1049 ( .A(KEYINPUT111), .B(KEYINPUT41), .Z(n960) );
  XNOR2_X1 U1050 ( .A(G1961), .B(G1976), .ZN(n959) );
  XNOR2_X1 U1051 ( .A(n960), .B(n959), .ZN(n970) );
  XOR2_X1 U1052 ( .A(KEYINPUT109), .B(G2474), .Z(n962) );
  XNOR2_X1 U1053 ( .A(G1996), .B(G1986), .ZN(n961) );
  XNOR2_X1 U1054 ( .A(n962), .B(n961), .ZN(n966) );
  XOR2_X1 U1055 ( .A(G1981), .B(G1971), .Z(n964) );
  XNOR2_X1 U1056 ( .A(G1991), .B(G1956), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(n964), .B(n963), .ZN(n965) );
  XOR2_X1 U1058 ( .A(n966), .B(n965), .Z(n968) );
  XNOR2_X1 U1059 ( .A(G1966), .B(KEYINPUT110), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(n968), .B(n967), .ZN(n969) );
  XOR2_X1 U1061 ( .A(n970), .B(n969), .Z(G229) );
  XOR2_X1 U1062 ( .A(G2100), .B(G2096), .Z(n972) );
  XNOR2_X1 U1063 ( .A(G2090), .B(KEYINPUT43), .ZN(n971) );
  XNOR2_X1 U1064 ( .A(n972), .B(n971), .ZN(n973) );
  XOR2_X1 U1065 ( .A(n973), .B(G2678), .Z(n975) );
  XNOR2_X1 U1066 ( .A(G2072), .B(KEYINPUT108), .ZN(n974) );
  XNOR2_X1 U1067 ( .A(n975), .B(n974), .ZN(n979) );
  XOR2_X1 U1068 ( .A(KEYINPUT42), .B(G2078), .Z(n977) );
  XNOR2_X1 U1069 ( .A(G2067), .B(G2084), .ZN(n976) );
  XNOR2_X1 U1070 ( .A(n977), .B(n976), .ZN(n978) );
  XNOR2_X1 U1071 ( .A(n979), .B(n978), .ZN(G227) );
  NAND2_X1 U1072 ( .A1(G130), .A2(n980), .ZN(n983) );
  NAND2_X1 U1073 ( .A1(G118), .A2(n981), .ZN(n982) );
  NAND2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n989) );
  NAND2_X1 U1075 ( .A1(G106), .A2(n530), .ZN(n985) );
  NAND2_X1 U1076 ( .A1(G142), .A2(n534), .ZN(n984) );
  NAND2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1078 ( .A(KEYINPUT45), .B(n986), .Z(n987) );
  XNOR2_X1 U1079 ( .A(KEYINPUT112), .B(n987), .ZN(n988) );
  NOR2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n1004) );
  XOR2_X1 U1081 ( .A(KEYINPUT117), .B(KEYINPUT46), .Z(n991) );
  XNOR2_X1 U1082 ( .A(KEYINPUT48), .B(KEYINPUT118), .ZN(n990) );
  XNOR2_X1 U1083 ( .A(n991), .B(n990), .ZN(n992) );
  XOR2_X1 U1084 ( .A(n992), .B(KEYINPUT114), .Z(n995) );
  XNOR2_X1 U1085 ( .A(n993), .B(KEYINPUT113), .ZN(n994) );
  XNOR2_X1 U1086 ( .A(n995), .B(n994), .ZN(n999) );
  XOR2_X1 U1087 ( .A(G160), .B(G162), .Z(n996) );
  XNOR2_X1 U1088 ( .A(n997), .B(n996), .ZN(n998) );
  XOR2_X1 U1089 ( .A(n999), .B(n998), .Z(n1002) );
  XNOR2_X1 U1090 ( .A(G164), .B(n1000), .ZN(n1001) );
  XNOR2_X1 U1091 ( .A(n1002), .B(n1001), .ZN(n1003) );
  XOR2_X1 U1092 ( .A(n1004), .B(n1003), .Z(n1005) );
  XNOR2_X1 U1093 ( .A(n1006), .B(n1005), .ZN(n1008) );
  XNOR2_X1 U1094 ( .A(n1008), .B(n1007), .ZN(n1009) );
  NOR2_X1 U1095 ( .A1(G37), .A2(n1009), .ZN(G395) );
  XNOR2_X1 U1096 ( .A(G286), .B(n1010), .ZN(n1011) );
  XNOR2_X1 U1097 ( .A(n1011), .B(G301), .ZN(n1015) );
  XNOR2_X1 U1098 ( .A(n1013), .B(n1012), .ZN(n1014) );
  XNOR2_X1 U1099 ( .A(n1015), .B(n1014), .ZN(n1016) );
  NOR2_X1 U1100 ( .A1(G37), .A2(n1016), .ZN(n1017) );
  XOR2_X1 U1101 ( .A(KEYINPUT119), .B(n1017), .Z(G397) );
  OR2_X1 U1102 ( .A1(n1023), .A2(G401), .ZN(n1020) );
  NOR2_X1 U1103 ( .A1(G229), .A2(G227), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(KEYINPUT49), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1022) );
  NOR2_X1 U1106 ( .A1(G395), .A2(G397), .ZN(n1021) );
  NAND2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(G225) );
  INV_X1 U1108 ( .A(G225), .ZN(G308) );
  INV_X1 U1109 ( .A(n1023), .ZN(G319) );
endmodule

