//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 1 1 0 0 0 0 1 0 0 0 0 0 0 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:59 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n540, new_n541,
    new_n542, new_n543, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n608, new_n609, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT66), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  XNOR2_X1  g040(.A(KEYINPUT3), .B(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G137), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT67), .B(G2105), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n471));
  NOR2_X1   g046(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AND2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  OAI21_X1  g050(.A(G125), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n473), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n470), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT68), .ZN(G160));
  NOR2_X1   g056(.A1(new_n474), .A2(new_n475), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(new_n473), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n482), .A2(G2105), .ZN(new_n484));
  AOI22_X1  g059(.A1(G124), .A2(new_n483), .B1(new_n484), .B2(G136), .ZN(new_n485));
  OAI221_X1 g060(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n473), .C2(G112), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n489), .A2(new_n491), .A3(G2104), .ZN(new_n492));
  AND2_X1   g067(.A1(G126), .A2(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n493), .B1(new_n474), .B2(new_n475), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(G138), .B1(new_n474), .B2(new_n475), .ZN(new_n496));
  OAI21_X1  g071(.A(KEYINPUT4), .B1(new_n496), .B2(new_n468), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n473), .A2(new_n466), .A3(new_n498), .A4(G138), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n495), .B1(new_n497), .B2(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT6), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT69), .B1(new_n501), .B2(G651), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n503), .A2(new_n504), .A3(KEYINPUT6), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n502), .A2(new_n505), .B1(new_n501), .B2(G651), .ZN(new_n506));
  OR2_X1    g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XOR2_X1   g084(.A(KEYINPUT71), .B(G88), .Z(new_n510));
  NAND3_X1  g085(.A1(new_n506), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G62), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n512), .B1(new_n507), .B2(new_n508), .ZN(new_n513));
  AND2_X1   g088(.A1(G75), .A2(G543), .ZN(new_n514));
  OAI21_X1  g089(.A(G651), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n502), .A2(new_n505), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n501), .A2(G651), .ZN(new_n518));
  AND2_X1   g093(.A1(G50), .A2(G543), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT70), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n506), .A2(KEYINPUT70), .A3(new_n519), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n516), .A2(new_n524), .ZN(G166));
  NAND3_X1  g100(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n506), .A2(G543), .ZN(new_n527));
  INV_X1    g102(.A(G51), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(KEYINPUT72), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT72), .ZN(new_n531));
  OAI211_X1 g106(.A(new_n531), .B(new_n526), .C1(new_n527), .C2(new_n528), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n517), .A2(new_n518), .A3(new_n509), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G89), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n530), .A2(new_n532), .A3(new_n534), .A4(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  NAND3_X1  g114(.A1(new_n506), .A2(G52), .A3(G543), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  OAI221_X1 g117(.A(new_n540), .B1(new_n541), .B2(new_n504), .C1(new_n542), .C2(new_n535), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(G171));
  INV_X1    g119(.A(new_n527), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G43), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n536), .A2(G81), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n548), .A2(new_n504), .ZN(new_n549));
  AND3_X1   g124(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  XOR2_X1   g130(.A(KEYINPUT75), .B(G65), .Z(new_n556));
  INV_X1    g131(.A(KEYINPUT74), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n509), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n507), .A2(KEYINPUT74), .A3(new_n508), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n556), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AND2_X1   g135(.A1(G78), .A2(G543), .ZN(new_n561));
  OAI21_X1  g136(.A(G651), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n536), .A2(G91), .ZN(new_n563));
  AND2_X1   g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n517), .A2(G53), .A3(G543), .A4(new_n518), .ZN(new_n565));
  AND2_X1   g140(.A1(KEYINPUT73), .A2(KEYINPUT9), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n565), .B(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n564), .A2(new_n567), .ZN(G299));
  XNOR2_X1  g143(.A(new_n543), .B(KEYINPUT76), .ZN(G301));
  NAND2_X1  g144(.A1(new_n516), .A2(new_n524), .ZN(G303));
  NAND4_X1  g145(.A1(new_n517), .A2(G49), .A3(G543), .A4(new_n518), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n572));
  INV_X1    g147(.A(G87), .ZN(new_n573));
  OAI211_X1 g148(.A(new_n571), .B(new_n572), .C1(new_n535), .C2(new_n573), .ZN(G288));
  NAND3_X1  g149(.A1(new_n506), .A2(G86), .A3(new_n509), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n517), .A2(G48), .A3(G543), .A4(new_n518), .ZN(new_n576));
  INV_X1    g151(.A(G61), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n577), .B1(new_n507), .B2(new_n508), .ZN(new_n578));
  AND2_X1   g153(.A1(G73), .A2(G543), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n575), .A2(new_n576), .A3(new_n580), .ZN(G305));
  AOI22_X1  g156(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n504), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT77), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n583), .B(new_n584), .ZN(new_n585));
  XNOR2_X1  g160(.A(KEYINPUT78), .B(G47), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n545), .A2(new_n586), .B1(new_n536), .B2(G85), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n585), .A2(new_n587), .ZN(G290));
  INV_X1    g163(.A(G66), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n589), .B1(new_n558), .B2(new_n559), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT79), .ZN(new_n591));
  AND2_X1   g166(.A1(G79), .A2(G543), .ZN(new_n592));
  OR3_X1    g167(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n591), .B1(new_n590), .B2(new_n592), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n593), .A2(G651), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n536), .A2(KEYINPUT10), .A3(G92), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n597));
  INV_X1    g172(.A(G92), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n535), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n596), .A2(new_n599), .B1(G54), .B2(new_n545), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n595), .A2(new_n600), .ZN(new_n601));
  MUX2_X1   g176(.A(new_n601), .B(G301), .S(G868), .Z(G321));
  XNOR2_X1  g177(.A(G321), .B(KEYINPUT80), .ZN(G284));
  INV_X1    g178(.A(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(G299), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(new_n604), .B2(G168), .ZN(G297));
  OAI21_X1  g181(.A(new_n605), .B1(new_n604), .B2(G168), .ZN(G280));
  INV_X1    g182(.A(new_n601), .ZN(new_n608));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(G860), .ZN(G148));
  NAND2_X1  g185(.A1(new_n608), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g189(.A1(new_n482), .A2(new_n463), .ZN(new_n615));
  XNOR2_X1  g190(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT13), .ZN(new_n618));
  INV_X1    g193(.A(G2100), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n619), .ZN(new_n621));
  AOI22_X1  g196(.A1(G123), .A2(new_n483), .B1(new_n484), .B2(G135), .ZN(new_n622));
  OAI221_X1 g197(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n473), .C2(G111), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(G2096), .Z(new_n625));
  NAND3_X1  g200(.A1(new_n620), .A2(new_n621), .A3(new_n625), .ZN(G156));
  XOR2_X1   g201(.A(KEYINPUT15), .B(G2435), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2438), .ZN(new_n628));
  XOR2_X1   g203(.A(G2427), .B(G2430), .Z(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(KEYINPUT83), .B(KEYINPUT14), .Z(new_n631));
  NAND2_X1  g206(.A1(new_n628), .A2(new_n629), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G1341), .B(G1348), .Z(new_n634));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n633), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G2451), .B(G2454), .Z(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(G14), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n642), .B1(new_n637), .B2(new_n640), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(G401));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  XNOR2_X1  g221(.A(G2072), .B(G2078), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT85), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT84), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT18), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(KEYINPUT86), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n648), .B1(new_n654), .B2(new_n647), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n655), .B1(new_n654), .B2(new_n647), .ZN(new_n656));
  INV_X1    g231(.A(new_n646), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT87), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n647), .B(KEYINPUT17), .Z(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g236(.A1(new_n660), .A2(new_n646), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n661), .B1(new_n663), .B2(new_n648), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2096), .B(G2100), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n653), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n666), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n668), .B1(new_n652), .B2(new_n664), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n669), .ZN(G227));
  XOR2_X1   g245(.A(G1991), .B(G1996), .Z(new_n671));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1956), .B(G2474), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1961), .B(G1966), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n679));
  OR2_X1    g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n678), .A2(new_n679), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n675), .A2(new_n676), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n674), .A2(new_n683), .ZN(new_n684));
  OR3_X1    g259(.A1(new_n674), .A2(new_n677), .A3(new_n683), .ZN(new_n685));
  NAND4_X1  g260(.A1(new_n680), .A2(new_n681), .A3(new_n684), .A4(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT90), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n690), .B1(new_n688), .B2(new_n689), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n671), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n693), .ZN(new_n695));
  INV_X1    g270(.A(new_n671), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n695), .A2(new_n696), .A3(new_n691), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1981), .B(G1986), .ZN(new_n698));
  AND3_X1   g273(.A1(new_n694), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n698), .B1(new_n694), .B2(new_n697), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(G229));
  INV_X1    g276(.A(G29), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G33), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT25), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G139), .B2(new_n484), .ZN(new_n706));
  NAND2_X1  g281(.A1(G115), .A2(G2104), .ZN(new_n707));
  INV_X1    g282(.A(G127), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(new_n482), .B2(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n473), .B1(new_n709), .B2(KEYINPUT95), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(KEYINPUT95), .B2(new_n709), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n706), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(KEYINPUT96), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT96), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n706), .A2(new_n714), .A3(new_n711), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n703), .B1(new_n717), .B2(new_n702), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(G2072), .Z(new_n719));
  NAND2_X1  g294(.A1(new_n702), .A2(G35), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT102), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n487), .B2(G29), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT29), .B(G2090), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(G27), .A2(G29), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G164), .B2(G29), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n724), .B1(G2078), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n702), .A2(G26), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT28), .Z(new_n729));
  AOI22_X1  g304(.A1(G128), .A2(new_n483), .B1(new_n484), .B2(G140), .ZN(new_n730));
  OAI221_X1 g305(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n473), .C2(G116), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n729), .B1(new_n732), .B2(G29), .ZN(new_n733));
  INV_X1    g308(.A(G2067), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(G2078), .ZN(new_n736));
  INV_X1    g311(.A(new_n726), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G16), .ZN(new_n739));
  AOI21_X1  g314(.A(KEYINPUT23), .B1(new_n739), .B2(G20), .ZN(new_n740));
  AND3_X1   g315(.A1(new_n739), .A2(KEYINPUT23), .A3(G20), .ZN(new_n741));
  AOI211_X1 g316(.A(new_n740), .B(new_n741), .C1(G299), .C2(G16), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT103), .B(G1956), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n727), .A2(new_n738), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n702), .A2(G32), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n484), .A2(G141), .ZN(new_n747));
  INV_X1    g322(.A(G105), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(new_n463), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n483), .A2(G129), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT26), .Z(new_n752));
  NAND2_X1  g327(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n746), .B1(new_n754), .B2(new_n702), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT27), .B(G1996), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT97), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n755), .B(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT31), .B(G11), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT98), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT30), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n761), .A2(G28), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n702), .B1(new_n761), .B2(G28), .ZN(new_n763));
  OAI221_X1 g338(.A(new_n760), .B1(new_n762), .B2(new_n763), .C1(new_n624), .C2(new_n702), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n758), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n550), .A2(G16), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G16), .B2(G19), .ZN(new_n767));
  INV_X1    g342(.A(G1341), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(G160), .A2(G29), .ZN(new_n771));
  INV_X1    g346(.A(G34), .ZN(new_n772));
  AOI21_X1  g347(.A(G29), .B1(new_n772), .B2(KEYINPUT24), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(KEYINPUT24), .B2(new_n772), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(G2084), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n767), .A2(new_n768), .ZN(new_n778));
  NOR4_X1   g353(.A1(new_n745), .A2(new_n770), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n719), .A2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT104), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n775), .A2(new_n776), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n782), .A2(KEYINPUT101), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n782), .A2(KEYINPUT101), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n742), .A2(new_n743), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(G4), .A2(G16), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(new_n608), .B2(G16), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT94), .B(G1348), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n739), .A2(G5), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G171), .B2(new_n739), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT99), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n794), .A2(G1961), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT100), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n739), .A2(G21), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G168), .B2(new_n739), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G1966), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n794), .A2(G1961), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n796), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n780), .A2(new_n781), .A3(new_n791), .A4(new_n803), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n719), .A2(new_n779), .A3(new_n790), .A4(new_n786), .ZN(new_n805));
  OAI21_X1  g380(.A(KEYINPUT104), .B1(new_n805), .B2(new_n802), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n739), .A2(G22), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G166), .B2(new_n739), .ZN(new_n808));
  INV_X1    g383(.A(G1971), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  MUX2_X1   g385(.A(G23), .B(G288), .S(G16), .Z(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT33), .B(G1976), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  MUX2_X1   g388(.A(G6), .B(G305), .S(G16), .Z(new_n814));
  XOR2_X1   g389(.A(KEYINPUT32), .B(G1981), .Z(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n810), .A2(new_n813), .A3(new_n816), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n817), .A2(KEYINPUT34), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(KEYINPUT34), .ZN(new_n819));
  MUX2_X1   g394(.A(G24), .B(G290), .S(G16), .Z(new_n820));
  AND2_X1   g395(.A1(new_n820), .A2(G1986), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n820), .A2(G1986), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n702), .A2(G25), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n483), .A2(G119), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT91), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n473), .A2(G107), .ZN(new_n827));
  OAI21_X1  g402(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n827), .A2(new_n829), .B1(new_n484), .B2(G131), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n823), .B1(new_n831), .B2(G29), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT35), .B(G1991), .Z(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NOR3_X1   g409(.A1(new_n821), .A2(new_n822), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n818), .A2(new_n819), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(KEYINPUT36), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(KEYINPUT93), .ZN(new_n838));
  XOR2_X1   g413(.A(KEYINPUT92), .B(KEYINPUT36), .Z(new_n839));
  OAI21_X1  g414(.A(new_n838), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n836), .A2(new_n839), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(KEYINPUT93), .ZN(new_n842));
  AOI22_X1  g417(.A1(new_n804), .A2(new_n806), .B1(new_n840), .B2(new_n842), .ZN(G311));
  NAND2_X1  g418(.A1(new_n840), .A2(new_n842), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n804), .A2(new_n806), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(G150));
  NAND3_X1  g421(.A1(new_n506), .A2(G55), .A3(G543), .ZN(new_n847));
  AOI22_X1  g422(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n848));
  INV_X1    g423(.A(G93), .ZN(new_n849));
  OAI221_X1 g424(.A(new_n847), .B1(new_n848), .B2(new_n504), .C1(new_n849), .C2(new_n535), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(G860), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT37), .Z(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(KEYINPUT105), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n536), .A2(G93), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n848), .A2(new_n504), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT105), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n854), .A2(new_n855), .A3(new_n856), .A4(new_n847), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n550), .A2(new_n853), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n859), .A2(KEYINPUT105), .A3(new_n850), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT38), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n608), .A2(G559), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT39), .ZN(new_n865));
  AOI21_X1  g440(.A(G860), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n866), .B1(new_n865), .B2(new_n864), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT106), .ZN(new_n868));
  AND2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n867), .A2(new_n868), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n852), .B1(new_n869), .B2(new_n870), .ZN(G145));
  INV_X1    g446(.A(new_n495), .ZN(new_n872));
  INV_X1    g447(.A(G138), .ZN(new_n873));
  OR2_X1    g448(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n874));
  NAND2_X1  g449(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n498), .B1(new_n876), .B2(new_n473), .ZN(new_n877));
  NOR3_X1   g452(.A1(new_n496), .A2(new_n468), .A3(KEYINPUT4), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n872), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n732), .B(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(new_n754), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n732), .B(G164), .ZN(new_n882));
  INV_X1    g457(.A(new_n754), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n716), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(KEYINPUT107), .B1(new_n884), .B2(new_n881), .ZN(new_n886));
  INV_X1    g461(.A(new_n712), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n881), .A2(new_n884), .A3(KEYINPUT107), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n885), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AOI22_X1  g465(.A1(G130), .A2(new_n483), .B1(new_n484), .B2(G142), .ZN(new_n891));
  OAI221_X1 g466(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n473), .C2(G118), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(new_n617), .ZN(new_n894));
  INV_X1    g469(.A(new_n831), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n894), .B(new_n895), .ZN(new_n896));
  OR3_X1    g471(.A1(new_n890), .A2(KEYINPUT108), .A3(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(G160), .B(new_n624), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(G162), .ZN(new_n899));
  OR2_X1    g474(.A1(new_n896), .A2(KEYINPUT108), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n899), .B1(new_n890), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n897), .A2(new_n901), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n890), .A2(new_n896), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n890), .A2(new_n896), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n899), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(G37), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n902), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g483(.A1(new_n850), .A2(new_n604), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n611), .B(new_n861), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT41), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n595), .A2(new_n567), .A3(new_n564), .A4(new_n600), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  AOI22_X1  g488(.A1(new_n595), .A2(new_n600), .B1(new_n564), .B2(new_n567), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n911), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n601), .A2(G299), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n916), .A2(KEYINPUT41), .A3(new_n912), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n910), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT109), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n913), .A2(new_n914), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n910), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n919), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n920), .B1(new_n919), .B2(new_n922), .ZN(new_n924));
  XNOR2_X1  g499(.A(G290), .B(G166), .ZN(new_n925));
  XOR2_X1   g500(.A(G305), .B(G288), .Z(new_n926));
  XNOR2_X1  g501(.A(new_n925), .B(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT42), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n927), .B(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n923), .B1(new_n924), .B2(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n927), .B(KEYINPUT42), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n931), .A2(new_n920), .A3(new_n922), .A4(new_n919), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n909), .B1(new_n933), .B2(new_n604), .ZN(G295));
  OAI21_X1  g509(.A(new_n909), .B1(new_n933), .B2(new_n604), .ZN(G331));
  NAND2_X1  g510(.A1(G286), .A2(new_n543), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(G301), .B2(G286), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n858), .A2(new_n860), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT76), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n543), .B(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(G168), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n861), .B1(new_n942), .B2(new_n936), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n921), .B1(new_n939), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n937), .A2(new_n938), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n942), .A2(new_n861), .A3(new_n936), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n915), .A2(new_n945), .A3(new_n917), .A4(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n927), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT43), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n927), .A2(new_n944), .A3(new_n947), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n950), .A2(new_n951), .A3(new_n906), .A4(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT110), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n950), .A2(new_n906), .A3(new_n952), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n956));
  AOI21_X1  g531(.A(G37), .B1(new_n948), .B2(new_n949), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT110), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n957), .A2(new_n958), .A3(new_n951), .A4(new_n952), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n954), .A2(new_n956), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n956), .A2(KEYINPUT44), .A3(new_n953), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(G397));
  XNOR2_X1  g539(.A(KEYINPUT111), .B(KEYINPUT45), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n965), .B1(G164), .B2(G1384), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G40), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n469), .A2(new_n968), .A3(new_n478), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  XOR2_X1   g546(.A(new_n831), .B(new_n833), .Z(new_n972));
  XNOR2_X1  g547(.A(new_n754), .B(G1996), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n732), .B(new_n734), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(G290), .B(G1986), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n971), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(G164), .A2(G1384), .ZN(new_n980));
  INV_X1    g555(.A(new_n965), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n982), .B(new_n969), .C1(KEYINPUT45), .C2(new_n980), .ZN(new_n983));
  INV_X1    g558(.A(G1966), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT50), .ZN(new_n986));
  INV_X1    g561(.A(G1384), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n879), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n988), .A2(new_n969), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n776), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n985), .A2(G168), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(G8), .ZN(new_n993));
  AOI21_X1  g568(.A(G168), .B1(new_n985), .B2(new_n991), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT51), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n992), .A2(new_n996), .A3(G8), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT62), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n470), .A2(G40), .A3(new_n479), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n879), .A2(new_n987), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1000), .B1(new_n1001), .B2(new_n965), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n879), .A2(KEYINPUT45), .A3(new_n987), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1002), .A2(new_n736), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n988), .A2(new_n989), .A3(new_n969), .ZN(new_n1006));
  XOR2_X1   g581(.A(KEYINPUT122), .B(G1961), .Z(new_n1007));
  AOI22_X1  g582(.A1(new_n1004), .A2(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  OR2_X1    g583(.A1(new_n980), .A2(KEYINPUT45), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1005), .A2(G2078), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1009), .A2(new_n982), .A3(new_n969), .A4(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(G301), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(G305), .A2(G1981), .ZN(new_n1013));
  INV_X1    g588(.A(G1981), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n575), .A2(new_n1014), .A3(new_n580), .A4(new_n576), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT49), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1013), .A2(KEYINPUT49), .A3(new_n1015), .ZN(new_n1019));
  INV_X1    g594(.A(G8), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1020), .B1(new_n980), .B2(new_n969), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1018), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n980), .A2(new_n969), .ZN(new_n1023));
  INV_X1    g598(.A(G1976), .ZN(new_n1024));
  OR2_X1    g599(.A1(G288), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1023), .A2(new_n1025), .A3(G8), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT52), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT52), .B1(G288), .B2(new_n1024), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1021), .A2(new_n1025), .A3(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1022), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1003), .A2(new_n966), .A3(new_n969), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n809), .ZN(new_n1032));
  XOR2_X1   g607(.A(KEYINPUT112), .B(G2090), .Z(new_n1033));
  NAND4_X1  g608(.A1(new_n988), .A2(new_n989), .A3(new_n969), .A4(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1020), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1020), .B1(new_n516), .B2(new_n524), .ZN(new_n1036));
  NAND2_X1  g611(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1037), .ZN(new_n1039));
  NOR2_X1   g614(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  AOI211_X1 g617(.A(new_n1020), .B(new_n1042), .C1(new_n516), .C2(new_n524), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT114), .B1(new_n1038), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1036), .A2(new_n1041), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1045), .B(new_n1046), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1044), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1030), .B1(new_n1035), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1045), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1050));
  AOI22_X1  g625(.A1(new_n990), .A2(new_n1033), .B1(new_n1031), .B2(new_n809), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1050), .B1(new_n1051), .B2(new_n1020), .ZN(new_n1052));
  AND2_X1   g627(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT62), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n995), .A2(new_n1054), .A3(new_n997), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n999), .A2(new_n1012), .A3(new_n1053), .A4(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT115), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1048), .A2(new_n1035), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1022), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1059));
  NAND2_X1  g634(.A1(G168), .A2(G8), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1060), .B1(new_n985), .B2(new_n991), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1058), .A2(new_n1052), .A3(new_n1059), .A4(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT63), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1049), .A2(KEYINPUT63), .A3(new_n1052), .A4(new_n1061), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1021), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1015), .ZN(new_n1068));
  NOR2_X1   g643(.A1(G288), .A2(G1976), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1068), .B1(new_n1022), .B2(new_n1069), .ZN(new_n1070));
  OAI22_X1  g645(.A1(new_n1058), .A2(new_n1030), .B1(new_n1067), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1057), .B1(new_n1066), .B2(new_n1072), .ZN(new_n1073));
  AOI211_X1 g648(.A(KEYINPUT115), .B(new_n1071), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1056), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1005), .B1(new_n1031), .B2(G2078), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1011), .A2(new_n1076), .A3(G301), .A4(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT124), .ZN(new_n1079));
  XNOR2_X1  g654(.A(new_n1078), .B(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT123), .B1(new_n967), .B2(new_n1000), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1082), .A2(new_n1003), .A3(new_n1010), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n967), .A2(KEYINPUT123), .A3(new_n1000), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1076), .B(new_n1077), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1081), .B1(new_n1085), .B2(G171), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1080), .A2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1085), .A2(new_n941), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1081), .B1(new_n1088), .B2(new_n1012), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1087), .A2(new_n998), .A3(new_n1089), .A4(new_n1053), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n1091));
  XOR2_X1   g666(.A(KEYINPUT58), .B(G1341), .Z(new_n1092));
  NAND2_X1  g667(.A1(new_n1023), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(G1996), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1003), .A2(new_n966), .A3(new_n1094), .A4(new_n969), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n859), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT59), .B1(new_n1096), .B2(KEYINPUT119), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1096), .A2(KEYINPUT118), .ZN(new_n1099));
  NAND3_X1  g674(.A1(KEYINPUT118), .A2(KEYINPUT119), .A3(KEYINPUT59), .ZN(new_n1100));
  AOI211_X1 g675(.A(new_n859), .B(new_n1100), .C1(new_n1093), .C2(new_n1095), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(KEYINPUT56), .B(G2072), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1003), .A2(new_n966), .A3(new_n969), .A4(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT116), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1104), .B(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(G1956), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1006), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n567), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n562), .A2(new_n563), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT57), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT57), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n564), .A2(new_n1112), .A3(new_n567), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1108), .A2(new_n1111), .A3(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT61), .B1(new_n1106), .B2(new_n1114), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1113), .A2(new_n1111), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1002), .A2(new_n1105), .A3(new_n1003), .A4(new_n1103), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1104), .A2(KEYINPUT116), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1116), .B1(new_n1119), .B2(new_n1108), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1098), .B(new_n1102), .C1(new_n1115), .C2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1116), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1108), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1124), .B1(new_n1106), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1119), .A2(new_n1108), .A3(new_n1116), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1123), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1091), .B1(new_n1121), .B2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1106), .A2(new_n1114), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1122), .B1(new_n1130), .B2(new_n1120), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1126), .A2(KEYINPUT61), .A3(new_n1127), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n1097), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1131), .A2(new_n1132), .A3(KEYINPUT121), .A4(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1023), .A2(G2067), .ZN(new_n1135));
  INV_X1    g710(.A(G1348), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1135), .B1(new_n1136), .B2(new_n1006), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n1137), .A2(KEYINPUT60), .A3(new_n601), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n601), .B1(new_n1137), .B2(KEYINPUT60), .ZN(new_n1139));
  OAI22_X1  g714(.A1(new_n1138), .A2(new_n1139), .B1(KEYINPUT60), .B2(new_n1137), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1129), .A2(new_n1134), .A3(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1137), .A2(new_n601), .ZN(new_n1142));
  XOR2_X1   g717(.A(new_n1142), .B(KEYINPUT117), .Z(new_n1143));
  OAI21_X1  g718(.A(new_n1127), .B1(new_n1143), .B2(new_n1120), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1090), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n979), .B1(new_n1075), .B2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n970), .B1(new_n974), .B2(new_n754), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1147), .B(KEYINPUT126), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n970), .A2(G1996), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n1149), .B(KEYINPUT46), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  XOR2_X1   g726(.A(new_n1151), .B(KEYINPUT47), .Z(new_n1152));
  NAND2_X1  g727(.A1(new_n895), .A2(new_n833), .ZN(new_n1153));
  OAI22_X1  g728(.A1(new_n975), .A2(new_n1153), .B1(G2067), .B2(new_n732), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(new_n971), .ZN(new_n1155));
  XOR2_X1   g730(.A(new_n1155), .B(KEYINPUT125), .Z(new_n1156));
  OR3_X1    g731(.A1(new_n970), .A2(G290), .A3(G1986), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1157), .ZN(new_n1158));
  AOI22_X1  g733(.A1(new_n977), .A2(new_n971), .B1(KEYINPUT48), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1159), .B1(KEYINPUT48), .B2(new_n1158), .ZN(new_n1160));
  AND3_X1   g735(.A1(new_n1152), .A2(new_n1156), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1146), .A2(new_n1161), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g737(.A1(new_n644), .A2(G319), .ZN(new_n1164));
  INV_X1    g738(.A(new_n1164), .ZN(new_n1165));
  INV_X1    g739(.A(KEYINPUT127), .ZN(new_n1166));
  NAND4_X1  g740(.A1(new_n1165), .A2(new_n1166), .A3(new_n667), .A4(new_n669), .ZN(new_n1167));
  OAI21_X1  g741(.A(KEYINPUT127), .B1(G227), .B2(new_n1164), .ZN(new_n1168));
  OAI211_X1 g742(.A(new_n1167), .B(new_n1168), .C1(new_n699), .C2(new_n700), .ZN(new_n1169));
  INV_X1    g743(.A(new_n1169), .ZN(new_n1170));
  AND3_X1   g744(.A1(new_n960), .A2(new_n1170), .A3(new_n907), .ZN(G308));
  NAND3_X1  g745(.A1(new_n960), .A2(new_n1170), .A3(new_n907), .ZN(G225));
endmodule


