//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 0 1 0 1 1 0 1 0 0 0 1 1 0 1 0 1 1 0 1 0 0 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 0 0 0 1 0 0 1 0 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942;
  INV_X1    g000(.A(KEYINPUT81), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT10), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G143), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G146), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT1), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G128), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  OR2_X1    g009(.A1(KEYINPUT64), .A2(G143), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(KEYINPUT64), .A2(G143), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n196), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n195), .B1(new_n199), .B2(KEYINPUT1), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n194), .B1(new_n192), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G104), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G107), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n202), .A2(G107), .ZN(new_n205));
  OAI21_X1  g019(.A(G101), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT3), .B1(new_n202), .B2(G107), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n208));
  INV_X1    g022(.A(G107), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n209), .A3(G104), .ZN(new_n210));
  INV_X1    g024(.A(G101), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n207), .A2(new_n210), .A3(new_n211), .A4(new_n203), .ZN(new_n212));
  AND2_X1   g026(.A1(new_n206), .A2(new_n212), .ZN(new_n213));
  AND3_X1   g027(.A1(new_n201), .A2(KEYINPUT80), .A3(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(KEYINPUT80), .B1(new_n201), .B2(new_n213), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n188), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G134), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(G137), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT65), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n220), .A2(KEYINPUT11), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n220), .A2(KEYINPUT11), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n219), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G131), .ZN(new_n224));
  INV_X1    g038(.A(G137), .ZN(new_n225));
  OAI211_X1 g039(.A(G134), .B(new_n225), .C1(new_n220), .C2(KEYINPUT11), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n217), .A2(G137), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n223), .A2(new_n224), .A3(new_n226), .A4(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT65), .B(KEYINPUT11), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n226), .B(new_n227), .C1(new_n229), .C2(new_n218), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G131), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT0), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n234), .A2(new_n195), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n192), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(KEYINPUT0), .A2(G128), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n189), .A2(G146), .ZN(new_n239));
  AOI211_X1 g053(.A(new_n235), .B(new_n238), .C1(new_n199), .C2(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT67), .B1(new_n237), .B2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n235), .B1(new_n199), .B2(new_n239), .ZN(new_n242));
  INV_X1    g056(.A(new_n238), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n242), .A2(new_n243), .B1(new_n192), .B2(new_n235), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT67), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n241), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n207), .A2(new_n210), .A3(new_n203), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(new_n249), .A3(G101), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(G101), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(KEYINPUT4), .A3(new_n212), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n247), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n199), .A2(new_n239), .ZN(new_n254));
  OAI21_X1  g068(.A(G128), .B1(new_n190), .B2(new_n193), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n194), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(KEYINPUT10), .A3(new_n213), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n216), .A2(new_n233), .A3(new_n253), .A4(new_n258), .ZN(new_n259));
  OAI22_X1  g073(.A1(new_n214), .A2(new_n215), .B1(new_n257), .B2(new_n213), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n260), .A2(KEYINPUT12), .A3(new_n232), .ZN(new_n261));
  AOI21_X1  g075(.A(KEYINPUT12), .B1(new_n260), .B2(new_n232), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n259), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(G110), .B(G140), .ZN(new_n264));
  INV_X1    g078(.A(G953), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n265), .A2(G227), .ZN(new_n266));
  XOR2_X1   g080(.A(new_n264), .B(new_n266), .Z(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n263), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n259), .A2(new_n267), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n216), .A2(new_n253), .A3(new_n258), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(new_n232), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(G902), .B1(new_n269), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G469), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n187), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  XOR2_X1   g091(.A(KEYINPUT73), .B(G902), .Z(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  AND3_X1   g093(.A1(new_n259), .A2(KEYINPUT82), .A3(new_n267), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n261), .A2(new_n262), .ZN(new_n281));
  AOI21_X1  g095(.A(KEYINPUT82), .B1(new_n259), .B2(new_n267), .ZN(new_n282));
  NOR3_X1   g096(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n267), .B1(new_n273), .B2(new_n259), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n276), .B(new_n279), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  AOI22_X1  g099(.A1(new_n263), .A2(new_n268), .B1(new_n271), .B2(new_n273), .ZN(new_n286));
  OAI211_X1 g100(.A(KEYINPUT81), .B(G469), .C1(new_n286), .C2(G902), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n277), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(G214), .B1(G237), .B2(G902), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  XOR2_X1   g104(.A(G116), .B(G119), .Z(new_n291));
  XNOR2_X1  g105(.A(KEYINPUT2), .B(G113), .ZN(new_n292));
  OR2_X1    g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n292), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(new_n252), .A3(new_n250), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT5), .ZN(new_n297));
  INV_X1    g111(.A(G119), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n298), .A3(G116), .ZN(new_n299));
  OAI211_X1 g113(.A(G113), .B(new_n299), .C1(new_n291), .C2(new_n297), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n213), .A2(new_n293), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n296), .A2(new_n301), .ZN(new_n302));
  XOR2_X1   g116(.A(G110), .B(G122), .Z(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT6), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n303), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n296), .A2(new_n307), .A3(new_n301), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT83), .ZN(new_n309));
  OR2_X1    g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n309), .ZN(new_n311));
  AOI22_X1  g125(.A1(new_n310), .A2(new_n311), .B1(new_n303), .B2(new_n302), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n306), .B1(new_n312), .B2(new_n305), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT85), .B(G224), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n265), .ZN(new_n315));
  XOR2_X1   g129(.A(new_n315), .B(KEYINPUT86), .Z(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(KEYINPUT84), .ZN(new_n317));
  INV_X1    g131(.A(G125), .ZN(new_n318));
  MUX2_X1   g132(.A(new_n244), .B(new_n257), .S(new_n318), .Z(new_n319));
  XNOR2_X1  g133(.A(new_n317), .B(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n313), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT7), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  AND2_X1   g137(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n319), .A2(new_n323), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n303), .B(KEYINPUT8), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n300), .A2(new_n293), .ZN(new_n327));
  OR2_X1    g141(.A1(new_n327), .A2(new_n213), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n326), .B1(new_n328), .B2(new_n301), .ZN(new_n329));
  NOR3_X1   g143(.A1(new_n324), .A2(new_n325), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n310), .A2(new_n311), .ZN(new_n331));
  AOI21_X1  g145(.A(G902), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n321), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(G210), .B1(G237), .B2(G902), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n321), .A2(new_n334), .A3(new_n332), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n290), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G221), .ZN(new_n339));
  XOR2_X1   g153(.A(KEYINPUT9), .B(G234), .Z(new_n340));
  INV_X1    g154(.A(G902), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  XOR2_X1   g156(.A(new_n342), .B(KEYINPUT79), .Z(new_n343));
  NAND3_X1  g157(.A1(new_n288), .A2(new_n338), .A3(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G237), .ZN(new_n346));
  AND4_X1   g160(.A1(KEYINPUT87), .A2(new_n346), .A3(new_n265), .A4(G214), .ZN(new_n347));
  NOR2_X1   g161(.A1(G237), .A2(G953), .ZN(new_n348));
  AOI21_X1  g162(.A(KEYINPUT87), .B1(new_n348), .B2(G214), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n191), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT88), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n348), .A2(G143), .A3(G214), .ZN(new_n353));
  OAI211_X1 g167(.A(KEYINPUT88), .B(new_n191), .C1(new_n347), .C2(new_n349), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(G131), .ZN(new_n356));
  XNOR2_X1  g170(.A(G125), .B(G140), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT19), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n357), .B1(KEYINPUT90), .B2(new_n358), .ZN(new_n359));
  XOR2_X1   g173(.A(KEYINPUT90), .B(KEYINPUT19), .Z(new_n360));
  AOI21_X1  g174(.A(new_n359), .B1(new_n357), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n197), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT76), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n357), .A2(new_n363), .A3(KEYINPUT16), .ZN(new_n364));
  INV_X1    g178(.A(G140), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G125), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n318), .A2(G140), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n366), .A2(new_n367), .A3(KEYINPUT16), .ZN(new_n368));
  OAI21_X1  g182(.A(KEYINPUT76), .B1(new_n366), .B2(KEYINPUT16), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n364), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G146), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n362), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n356), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n355), .A2(KEYINPUT18), .A3(G131), .ZN(new_n374));
  AND2_X1   g188(.A1(KEYINPUT18), .A2(G131), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n352), .A2(new_n376), .A3(new_n353), .A4(new_n354), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n357), .B(new_n197), .ZN(new_n378));
  AND4_X1   g192(.A1(KEYINPUT89), .A2(new_n374), .A3(new_n377), .A4(new_n378), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n377), .A2(new_n378), .ZN(new_n380));
  AOI21_X1  g194(.A(KEYINPUT89), .B1(new_n380), .B2(new_n374), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n373), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT91), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(G113), .B(G122), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n385), .B(new_n202), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  OAI211_X1 g201(.A(KEYINPUT91), .B(new_n373), .C1(new_n379), .C2(new_n381), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n384), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(KEYINPUT92), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT93), .ZN(new_n391));
  OR3_X1    g205(.A1(new_n356), .A2(new_n391), .A3(KEYINPUT17), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n355), .A2(KEYINPUT17), .A3(G131), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT77), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n364), .B(new_n197), .C1(new_n368), .C2(new_n369), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n371), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n370), .A2(KEYINPUT77), .A3(G146), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n391), .B1(new_n356), .B2(KEYINPUT17), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n392), .A2(new_n393), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  OR2_X1    g214(.A1(new_n379), .A2(new_n381), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n400), .A2(new_n386), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT92), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n384), .A2(new_n403), .A3(new_n387), .A4(new_n388), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n390), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(G475), .A2(G902), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT94), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n405), .A2(KEYINPUT94), .A3(new_n406), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(KEYINPUT20), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n191), .A2(G128), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT96), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n195), .A2(G143), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n191), .A2(KEYINPUT96), .A3(G128), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n417), .B(G134), .ZN(new_n418));
  XNOR2_X1  g232(.A(KEYINPUT95), .B(G122), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G116), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n209), .B1(new_n420), .B2(KEYINPUT14), .ZN(new_n421));
  INV_X1    g235(.A(G122), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n420), .B1(G116), .B2(new_n422), .ZN(new_n423));
  XOR2_X1   g237(.A(new_n421), .B(new_n423), .Z(new_n424));
  NAND2_X1  g238(.A1(new_n418), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n425), .B(KEYINPUT97), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT13), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n217), .B1(new_n415), .B2(new_n427), .ZN(new_n428));
  XOR2_X1   g242(.A(new_n417), .B(new_n428), .Z(new_n429));
  XNOR2_X1  g243(.A(new_n423), .B(G107), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n340), .A2(G217), .A3(new_n265), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n433), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n426), .A2(new_n431), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n278), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(G478), .ZN(new_n438));
  NOR3_X1   g252(.A1(new_n437), .A2(KEYINPUT15), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G952), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n440), .A2(G953), .ZN(new_n441));
  INV_X1    g255(.A(G234), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n441), .B1(new_n442), .B2(new_n346), .ZN(new_n443));
  AOI211_X1 g257(.A(new_n265), .B(new_n279), .C1(G234), .C2(G237), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  XOR2_X1   g259(.A(KEYINPUT21), .B(G898), .Z(new_n446));
  OAI21_X1  g260(.A(new_n443), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n438), .A2(KEYINPUT15), .ZN(new_n449));
  AOI211_X1 g263(.A(new_n278), .B(new_n449), .C1(new_n434), .C2(new_n436), .ZN(new_n450));
  NOR3_X1   g264(.A1(new_n439), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n402), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n386), .B1(new_n400), .B2(new_n401), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n341), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(G475), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT20), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n407), .A2(new_n408), .A3(new_n456), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n411), .A2(new_n451), .A3(new_n455), .A4(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT98), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n458), .A2(new_n459), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n345), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT99), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI211_X1 g279(.A(KEYINPUT99), .B(new_n345), .C1(new_n461), .C2(new_n462), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n247), .A2(new_n232), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n295), .B(KEYINPUT69), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n219), .A2(new_n227), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT66), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(new_n472), .A3(G131), .ZN(new_n473));
  AND2_X1   g287(.A1(new_n228), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n472), .B1(new_n471), .B2(G131), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n475), .B1(new_n194), .B2(new_n256), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n468), .A2(new_n470), .A3(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  OR2_X1    g293(.A1(new_n479), .A2(KEYINPUT28), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT71), .ZN(new_n481));
  AOI22_X1  g295(.A1(new_n474), .A2(new_n476), .B1(new_n232), .B2(new_n244), .ZN(new_n482));
  INV_X1    g296(.A(new_n295), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n478), .A2(new_n484), .ZN(new_n485));
  NOR3_X1   g299(.A1(new_n482), .A2(new_n481), .A3(new_n483), .ZN(new_n486));
  OAI21_X1  g300(.A(KEYINPUT28), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n480), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n489), .B(G101), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n348), .A2(G210), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n490), .B(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n468), .A2(KEYINPUT68), .A3(KEYINPUT30), .A4(new_n477), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n233), .B1(new_n241), .B2(new_n246), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n474), .A2(new_n476), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT30), .ZN(new_n497));
  NOR3_X1   g311(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT68), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n499), .B1(new_n482), .B2(KEYINPUT30), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n494), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n479), .B1(new_n501), .B2(new_n295), .ZN(new_n502));
  INV_X1    g316(.A(new_n492), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(KEYINPUT29), .B1(new_n493), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n469), .B1(new_n495), .B2(new_n496), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT72), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n478), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n468), .A2(new_n470), .A3(KEYINPUT72), .A4(new_n477), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(KEYINPUT28), .A3(new_n509), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n510), .A2(new_n480), .A3(KEYINPUT29), .A4(new_n492), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n279), .ZN(new_n512));
  OAI21_X1  g326(.A(G472), .B1(new_n505), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n501), .A2(new_n295), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT70), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n514), .A2(new_n515), .A3(new_n478), .A4(new_n492), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(KEYINPUT31), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n488), .A2(new_n503), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT31), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n502), .A2(new_n515), .A3(new_n519), .A4(new_n492), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n517), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT32), .ZN(new_n522));
  NOR2_X1   g336(.A1(G472), .A2(G902), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n522), .B1(new_n521), .B2(new_n523), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n513), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n265), .A2(G221), .A3(G234), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(KEYINPUT22), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(new_n225), .ZN(new_n529));
  INV_X1    g343(.A(G110), .ZN(new_n530));
  OAI21_X1  g344(.A(KEYINPUT23), .B1(new_n195), .B2(G119), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n531), .B(KEYINPUT74), .C1(new_n298), .C2(G128), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n298), .A2(G128), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT74), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n533), .B1(new_n534), .B2(KEYINPUT23), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n530), .B1(new_n536), .B2(KEYINPUT75), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n537), .B1(KEYINPUT75), .B2(new_n536), .ZN(new_n538));
  XOR2_X1   g352(.A(KEYINPUT24), .B(G110), .Z(new_n539));
  XNOR2_X1  g353(.A(G119), .B(G128), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n538), .A2(new_n396), .A3(new_n397), .A4(new_n541), .ZN(new_n542));
  OAI22_X1  g356(.A1(new_n536), .A2(G110), .B1(new_n540), .B2(new_n539), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n357), .A2(new_n197), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(new_n371), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT78), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n529), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n546), .A2(new_n547), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n548), .B(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT25), .B1(new_n550), .B2(new_n278), .ZN(new_n551));
  OAI21_X1  g365(.A(G217), .B1(new_n278), .B2(new_n442), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT25), .ZN(new_n554));
  INV_X1    g368(.A(new_n548), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n555), .A2(new_n549), .ZN(new_n556));
  NOR3_X1   g370(.A1(new_n548), .A2(new_n547), .A3(new_n546), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n554), .B(new_n279), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n551), .A2(new_n553), .A3(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n553), .A2(G902), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n560), .B1(new_n556), .B2(new_n557), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n526), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n467), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(G101), .ZN(G3));
  AND2_X1   g381(.A1(new_n521), .A2(new_n523), .ZN(new_n568));
  INV_X1    g382(.A(G472), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n569), .B1(new_n521), .B2(new_n279), .ZN(new_n570));
  OR2_X1    g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NOR4_X1   g385(.A1(new_n571), .A2(new_n344), .A3(new_n448), .A4(new_n562), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n411), .A2(new_n455), .A3(new_n457), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT33), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n434), .A2(new_n574), .A3(new_n436), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n574), .B1(new_n434), .B2(new_n436), .ZN(new_n576));
  OAI211_X1 g390(.A(G478), .B(new_n279), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  XOR2_X1   g391(.A(KEYINPUT100), .B(G478), .Z(new_n578));
  OAI21_X1  g392(.A(new_n577), .B1(new_n437), .B2(new_n578), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n573), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n572), .A2(new_n580), .ZN(new_n581));
  XOR2_X1   g395(.A(KEYINPUT34), .B(G104), .Z(new_n582));
  XNOR2_X1  g396(.A(new_n581), .B(new_n582), .ZN(G6));
  NOR2_X1   g397(.A1(new_n439), .A2(new_n450), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n411), .A2(new_n585), .A3(new_n455), .A4(new_n457), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n572), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT35), .B(G107), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(KEYINPUT101), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n588), .B(new_n590), .ZN(G9));
  NOR2_X1   g405(.A1(new_n529), .A2(KEYINPUT36), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n546), .B(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n560), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n559), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n571), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(KEYINPUT102), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n467), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(KEYINPUT37), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(new_n530), .ZN(G12));
  INV_X1    g415(.A(new_n513), .ZN(new_n602));
  INV_X1    g416(.A(new_n525), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n605), .A2(new_n344), .A3(new_n596), .ZN(new_n606));
  INV_X1    g420(.A(new_n443), .ZN(new_n607));
  INV_X1    g421(.A(G900), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n607), .B1(new_n444), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n586), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G128), .ZN(G30));
  NOR2_X1   g426(.A1(new_n502), .A2(new_n503), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n492), .B1(new_n508), .B2(new_n509), .ZN(new_n614));
  OR3_X1    g428(.A1(new_n613), .A2(G902), .A3(new_n614), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n603), .A2(new_n604), .B1(G472), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n616), .A2(new_n595), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n288), .A2(new_n343), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n609), .B(KEYINPUT39), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n617), .B1(new_n622), .B2(KEYINPUT40), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n623), .A2(new_n290), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n336), .A2(new_n337), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(KEYINPUT38), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n573), .A2(new_n585), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n627), .B1(new_n622), .B2(KEYINPUT40), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n624), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(new_n629), .B(new_n191), .Z(G45));
  INV_X1    g444(.A(new_n609), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n606), .A2(new_n580), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G146), .ZN(G48));
  NOR2_X1   g447(.A1(new_n283), .A2(new_n284), .ZN(new_n634));
  OAI21_X1  g448(.A(G469), .B1(new_n634), .B2(new_n278), .ZN(new_n635));
  INV_X1    g449(.A(new_n342), .ZN(new_n636));
  AND4_X1   g450(.A1(new_n338), .A2(new_n635), .A3(new_n636), .A4(new_n285), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n526), .A2(new_n637), .A3(new_n447), .A4(new_n563), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n573), .A2(new_n579), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT41), .B(G113), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G15));
  AND4_X1   g456(.A1(new_n447), .A2(new_n526), .A3(new_n637), .A4(new_n563), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT103), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n643), .A2(new_n644), .A3(new_n587), .ZN(new_n645));
  OAI21_X1  g459(.A(KEYINPUT103), .B1(new_n638), .B2(new_n586), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G116), .ZN(G18));
  NOR2_X1   g462(.A1(new_n605), .A2(new_n596), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n649), .B(new_n637), .C1(new_n461), .C2(new_n462), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G119), .ZN(G21));
  NAND2_X1  g465(.A1(new_n510), .A2(new_n480), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n503), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n517), .A2(new_n653), .A3(new_n520), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n654), .A2(new_n523), .ZN(new_n655));
  NOR4_X1   g469(.A1(new_n655), .A2(new_n570), .A3(new_n562), .A4(new_n448), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n656), .A2(new_n573), .A3(new_n585), .A4(new_n637), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G122), .ZN(G24));
  NAND4_X1  g472(.A1(new_n573), .A2(new_n579), .A3(new_n631), .A4(new_n637), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n655), .A2(new_n570), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n595), .ZN(new_n661));
  OR2_X1    g475(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT104), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(new_n318), .ZN(G27));
  NAND3_X1  g478(.A1(new_n573), .A2(new_n579), .A3(new_n631), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n336), .A2(new_n289), .A3(new_n337), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n285), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n275), .A2(new_n276), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n636), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n564), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT42), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n667), .A2(KEYINPUT105), .A3(new_n675), .A4(new_n671), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(new_n224), .ZN(G33));
  INV_X1    g492(.A(new_n666), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n671), .A2(new_n610), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G134), .ZN(G36));
  NOR2_X1   g495(.A1(new_n286), .A2(KEYINPUT45), .ZN(new_n682));
  OR3_X1    g496(.A1(new_n682), .A2(KEYINPUT106), .A3(new_n276), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n286), .A2(KEYINPUT45), .ZN(new_n684));
  OAI21_X1  g498(.A(KEYINPUT106), .B1(new_n682), .B2(new_n276), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(G469), .A2(G902), .ZN(new_n687));
  AOI21_X1  g501(.A(KEYINPUT46), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n668), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT46), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n686), .A2(new_n687), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n689), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n620), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n692), .A2(new_n636), .A3(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT107), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n411), .A2(new_n455), .A3(new_n457), .A4(new_n579), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT108), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(KEYINPUT43), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n700), .B1(new_n697), .B2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n702), .A2(new_n571), .A3(new_n595), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n704));
  OR2_X1    g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n666), .B1(new_n703), .B2(new_n704), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n696), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G137), .ZN(G39));
  INV_X1    g522(.A(KEYINPUT47), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n691), .A2(new_n690), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n710), .A2(new_n688), .A3(new_n668), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n709), .B1(new_n711), .B2(new_n342), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n692), .A2(KEYINPUT47), .A3(new_n636), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n605), .A2(new_n562), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n714), .A2(new_n667), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(KEYINPUT109), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT109), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n714), .A2(new_n719), .A3(new_n667), .A4(new_n716), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G140), .ZN(G42));
  INV_X1    g536(.A(new_n660), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n723), .A2(new_n562), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n702), .A2(new_n607), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n635), .A2(new_n285), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n342), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n626), .A2(new_n289), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n725), .A2(KEYINPUT50), .A3(new_n727), .A4(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT50), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n702), .A2(new_n607), .A3(new_n727), .A4(new_n724), .ZN(new_n731));
  INV_X1    g545(.A(new_n728), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT111), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n729), .A2(new_n733), .A3(KEYINPUT111), .ZN(new_n737));
  AOI21_X1  g551(.A(KEYINPUT51), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n712), .B(new_n713), .C1(new_n343), .C2(new_n726), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n739), .A2(new_n679), .A3(new_n725), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n616), .A2(new_n563), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n726), .A2(new_n342), .A3(new_n666), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n607), .ZN(new_n743));
  NOR4_X1   g557(.A1(new_n741), .A2(new_n743), .A3(new_n573), .A4(new_n579), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n697), .A2(new_n699), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n697), .A2(new_n701), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n607), .B(new_n742), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT112), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT112), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n702), .A2(new_n749), .A3(new_n607), .A4(new_n742), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n661), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n744), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n738), .A2(new_n740), .A3(new_n753), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n753), .A2(new_n734), .A3(KEYINPUT113), .ZN(new_n755));
  AOI21_X1  g569(.A(KEYINPUT113), .B1(new_n753), .B2(new_n734), .ZN(new_n756));
  INV_X1    g570(.A(new_n740), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n755), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n754), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n741), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n761), .A2(new_n580), .A3(new_n607), .A4(new_n742), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n564), .B1(new_n748), .B2(new_n750), .ZN(new_n763));
  OR2_X1    g577(.A1(KEYINPUT114), .A2(KEYINPUT48), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n765), .B1(KEYINPUT114), .B2(KEYINPUT48), .ZN(new_n766));
  INV_X1    g580(.A(new_n338), .ZN(new_n767));
  OAI221_X1 g581(.A(new_n441), .B1(new_n767), .B2(new_n731), .C1(new_n763), .C2(new_n764), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n760), .A2(new_n762), .A3(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n657), .B1(new_n639), .B2(new_n638), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n647), .A2(new_n774), .A3(new_n650), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n606), .B(new_n631), .C1(new_n580), .C2(new_n587), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n662), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n627), .A2(new_n767), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n670), .A2(new_n609), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n779), .A2(new_n617), .A3(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n776), .B1(new_n778), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n779), .A2(new_n617), .A3(new_n780), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n783), .A2(new_n777), .A3(new_n662), .A4(KEYINPUT52), .ZN(new_n784));
  AOI211_X1 g598(.A(new_n775), .B(new_n677), .C1(new_n782), .C2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n671), .A2(new_n610), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n618), .A2(new_n526), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n584), .A2(new_n631), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n787), .A2(new_n573), .A3(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n665), .A2(new_n723), .ZN(new_n790));
  INV_X1    g604(.A(new_n670), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n786), .B1(new_n792), .B2(new_n596), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n679), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n639), .A2(new_n586), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n572), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n465), .B(new_n466), .C1(new_n565), .C2(new_n598), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n794), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(KEYINPUT53), .B1(new_n785), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n782), .A2(new_n784), .ZN(new_n800));
  INV_X1    g614(.A(new_n775), .ZN(new_n801));
  INV_X1    g615(.A(new_n677), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n794), .A2(new_n796), .A3(new_n797), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(KEYINPUT54), .B1(new_n799), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT110), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n775), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n647), .A2(new_n774), .A3(new_n650), .A4(KEYINPUT110), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n805), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n798), .A2(new_n802), .A3(new_n800), .A4(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n805), .B1(new_n803), .B2(new_n804), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n807), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n760), .A2(KEYINPUT115), .A3(new_n762), .A4(new_n769), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n772), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n440), .A2(new_n265), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n697), .A2(new_n290), .A3(new_n626), .ZN(new_n821));
  XOR2_X1   g635(.A(new_n726), .B(KEYINPUT49), .Z(new_n822));
  NAND4_X1  g636(.A1(new_n821), .A2(new_n761), .A3(new_n343), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n820), .A2(new_n823), .ZN(G75));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n313), .B(new_n320), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(KEYINPUT55), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n812), .A2(new_n813), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n828), .A2(KEYINPUT116), .A3(new_n278), .A4(new_n335), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT56), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n279), .B1(new_n812), .B2(new_n813), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT116), .B1(new_n832), .B2(new_n335), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n825), .B(new_n827), .C1(new_n831), .C2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n809), .A2(new_n810), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n836), .A2(KEYINPUT53), .A3(new_n802), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n800), .A2(new_n794), .A3(new_n796), .A4(new_n797), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n278), .B(new_n335), .C1(new_n799), .C2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n842), .A2(new_n830), .A3(new_n829), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n825), .B1(new_n843), .B2(new_n827), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n265), .A2(G952), .ZN(new_n845));
  XOR2_X1   g659(.A(new_n845), .B(KEYINPUT118), .Z(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n840), .ZN(new_n848));
  OR2_X1    g662(.A1(new_n827), .A2(KEYINPUT56), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n835), .A2(new_n844), .A3(new_n850), .ZN(G51));
  INV_X1    g665(.A(KEYINPUT120), .ZN(new_n852));
  INV_X1    g666(.A(new_n845), .ZN(new_n853));
  OAI21_X1  g667(.A(KEYINPUT54), .B1(new_n799), .B2(new_n839), .ZN(new_n854));
  AOI22_X1  g668(.A1(new_n854), .A2(new_n815), .B1(KEYINPUT57), .B2(new_n687), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n687), .A2(KEYINPUT57), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n634), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  XOR2_X1   g671(.A(new_n686), .B(KEYINPUT119), .Z(new_n858));
  AND2_X1   g672(.A1(new_n832), .A2(new_n858), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n852), .B(new_n853), .C1(new_n857), .C2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n687), .A2(KEYINPUT57), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n814), .B1(new_n812), .B2(new_n813), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n856), .B(new_n861), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n634), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n859), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT120), .B1(new_n866), .B2(new_n845), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n860), .A2(new_n867), .ZN(G54));
  NAND3_X1  g682(.A1(new_n832), .A2(KEYINPUT58), .A3(G475), .ZN(new_n869));
  INV_X1    g683(.A(new_n405), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n869), .A2(new_n870), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n871), .A2(new_n872), .A3(new_n845), .ZN(G60));
  NOR2_X1   g687(.A1(new_n575), .A2(new_n576), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n874), .B(KEYINPUT121), .Z(new_n875));
  XOR2_X1   g689(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n876));
  NOR2_X1   g690(.A1(new_n438), .A2(new_n341), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n876), .B(new_n877), .ZN(new_n878));
  AOI211_X1 g692(.A(new_n875), .B(new_n878), .C1(new_n854), .C2(new_n815), .ZN(new_n879));
  OAI211_X1 g693(.A(KEYINPUT123), .B(new_n875), .C1(new_n816), .C2(new_n878), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT123), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n878), .B1(new_n807), .B2(new_n815), .ZN(new_n882));
  INV_X1    g696(.A(new_n875), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI211_X1 g698(.A(new_n846), .B(new_n879), .C1(new_n880), .C2(new_n884), .ZN(G63));
  NAND2_X1  g699(.A1(G217), .A2(G902), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n886), .B(KEYINPUT60), .Z(new_n887));
  NAND2_X1  g701(.A1(new_n828), .A2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n593), .ZN(new_n889));
  OR3_X1    g703(.A1(new_n888), .A2(KEYINPUT124), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n846), .B1(new_n888), .B2(new_n550), .ZN(new_n891));
  OAI21_X1  g705(.A(KEYINPUT124), .B1(new_n888), .B2(new_n889), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT61), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n890), .A2(KEYINPUT61), .A3(new_n891), .A4(new_n892), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(G66));
  AOI21_X1  g711(.A(new_n265), .B1(new_n446), .B2(new_n314), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n797), .A2(new_n801), .A3(new_n796), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n898), .B1(new_n899), .B2(new_n265), .ZN(new_n900));
  INV_X1    g714(.A(new_n313), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n901), .B1(G898), .B2(new_n265), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n900), .B(new_n902), .Z(G69));
  AOI21_X1  g717(.A(new_n265), .B1(G227), .B2(G900), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n501), .B(new_n361), .Z(new_n905));
  NOR3_X1   g719(.A1(new_n627), .A2(new_n767), .A3(new_n564), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n778), .B1(new_n696), .B2(new_n906), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n802), .A2(new_n680), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n721), .A2(new_n907), .A3(new_n707), .A4(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n265), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n608), .A2(G953), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(KEYINPUT126), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT126), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n910), .A2(new_n914), .A3(new_n911), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n905), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n905), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n629), .A2(new_n662), .A3(new_n777), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT62), .Z(new_n919));
  NAND4_X1  g733(.A1(new_n795), .A2(new_n565), .A3(new_n621), .A4(new_n679), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT125), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n919), .A2(new_n707), .A3(new_n721), .A4(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n917), .B1(new_n922), .B2(new_n265), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n904), .B1(new_n916), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n915), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n914), .B1(new_n910), .B2(new_n911), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n917), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n904), .ZN(new_n928));
  INV_X1    g742(.A(new_n923), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n924), .A2(new_n930), .ZN(G72));
  NAND2_X1  g745(.A1(G472), .A2(G902), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT63), .Z(new_n933));
  OAI21_X1  g747(.A(new_n933), .B1(new_n922), .B2(new_n899), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n613), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n933), .B1(new_n909), .B2(new_n899), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n504), .B(KEYINPUT127), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n845), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n613), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n933), .B1(new_n799), .B2(new_n806), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(new_n503), .B2(new_n502), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n939), .B1(new_n940), .B2(new_n942), .ZN(G57));
endmodule


