//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 1 0 0 1 1 1 0 1 1 0 1 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n763, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n864, new_n865, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980;
  INV_X1    g000(.A(KEYINPUT87), .ZN(new_n202));
  XNOR2_X1  g001(.A(G8gat), .B(G36gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  XNOR2_X1  g004(.A(G197gat), .B(G204gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT22), .ZN(new_n207));
  INV_X1    g006(.A(G211gat), .ZN(new_n208));
  INV_X1    g007(.A(G218gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n206), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G211gat), .B(G218gat), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(new_n206), .A3(new_n210), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT72), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT72), .B1(new_n214), .B2(new_n215), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(G226gat), .A2(G233gat), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G169gat), .ZN(new_n223));
  INV_X1    g022(.A(G176gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT26), .ZN(new_n226));
  NAND2_X1  g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NOR2_X1   g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229));
  AOI22_X1  g028(.A1(new_n229), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT66), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n228), .A2(new_n230), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT27), .B(G183gat), .ZN(new_n236));
  INV_X1    g035(.A(G190gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT28), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n236), .A2(KEYINPUT28), .A3(new_n237), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n235), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT25), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT23), .ZN(new_n245));
  OAI22_X1  g044(.A1(KEYINPUT64), .A2(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n227), .B(new_n245), .C1(new_n246), .C2(new_n248), .ZN(new_n249));
  AND3_X1   g048(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n251));
  OAI21_X1  g050(.A(G190gat), .B1(KEYINPUT24), .B2(G183gat), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n244), .B1(new_n249), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n252), .A2(new_n251), .ZN(new_n255));
  NAND3_X1  g054(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AND2_X1   g056(.A1(G169gat), .A2(G176gat), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n258), .B1(KEYINPUT23), .B2(new_n229), .ZN(new_n259));
  OR2_X1    g058(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n260), .A2(new_n225), .A3(new_n247), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n257), .A2(KEYINPUT25), .A3(new_n259), .A4(new_n261), .ZN(new_n262));
  AND3_X1   g061(.A1(new_n254), .A2(KEYINPUT65), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT65), .B1(new_n254), .B2(new_n262), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n222), .B(new_n243), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n222), .A2(KEYINPUT29), .ZN(new_n266));
  AND2_X1   g065(.A1(new_n254), .A2(new_n262), .ZN(new_n267));
  AOI22_X1  g066(.A1(new_n232), .A2(new_n234), .B1(new_n240), .B2(new_n241), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n220), .B1(new_n265), .B2(new_n269), .ZN(new_n270));
  NOR3_X1   g069(.A1(new_n267), .A2(new_n268), .A3(new_n221), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n243), .B1(new_n263), .B2(new_n264), .ZN(new_n272));
  XNOR2_X1  g071(.A(KEYINPUT73), .B(KEYINPUT29), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n274), .A2(new_n222), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n271), .B1(new_n272), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n270), .B1(new_n220), .B2(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(KEYINPUT85), .B(KEYINPUT37), .Z(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n277), .A2(KEYINPUT86), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT86), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n269), .ZN(new_n282));
  OR2_X1    g081(.A1(new_n218), .A2(new_n219), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n254), .A2(new_n262), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n243), .A2(new_n222), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT65), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n254), .A2(KEYINPUT65), .A3(new_n262), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n268), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n275), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n220), .B(new_n286), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n284), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n281), .B1(new_n293), .B2(new_n278), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n205), .B1(new_n280), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(KEYINPUT37), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT38), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n202), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT37), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n295), .B1(new_n300), .B2(new_n277), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n301), .A2(KEYINPUT87), .A3(KEYINPUT38), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n300), .B1(new_n276), .B2(new_n283), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n282), .A2(new_n220), .ZN(new_n304));
  AOI21_X1  g103(.A(KEYINPUT38), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n295), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT80), .B(KEYINPUT6), .ZN(new_n307));
  NOR2_X1   g106(.A1(G155gat), .A2(G162gat), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT75), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT2), .ZN(new_n311));
  AOI22_X1  g110(.A1(new_n310), .A2(new_n311), .B1(G155gat), .B2(G162gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(G141gat), .B(G148gat), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n311), .B1(G155gat), .B2(G162gat), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n309), .B(new_n312), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  AND2_X1   g114(.A1(G141gat), .A2(G148gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(G141gat), .A2(G148gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(G155gat), .ZN(new_n319));
  INV_X1    g118(.A(G162gat), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT2), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(KEYINPUT75), .B1(new_n319), .B2(new_n320), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n318), .B(new_n321), .C1(new_n308), .C2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n315), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(G134gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G127gat), .ZN(new_n326));
  INV_X1    g125(.A(G127gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G134gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G113gat), .B(G120gat), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n329), .B1(new_n330), .B2(KEYINPUT1), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT67), .ZN(new_n332));
  INV_X1    g131(.A(G113gat), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n332), .B1(new_n333), .B2(G120gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(G120gat), .ZN(new_n335));
  INV_X1    g134(.A(G120gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n336), .A2(KEYINPUT67), .A3(G113gat), .ZN(new_n337));
  AND3_X1   g136(.A1(new_n334), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT1), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n326), .A2(new_n328), .A3(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n331), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n340), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n334), .A2(new_n335), .A3(new_n337), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n345), .A2(new_n323), .A3(new_n315), .A4(new_n331), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT77), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n342), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(G225gat), .A2(G233gat), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n324), .A2(new_n341), .A3(KEYINPUT77), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n348), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n352), .A2(KEYINPUT5), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT76), .B1(new_n324), .B2(KEYINPUT3), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT76), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT3), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n315), .A2(new_n323), .A3(new_n355), .A4(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  AOI22_X1  g157(.A1(new_n324), .A2(KEYINPUT3), .B1(new_n345), .B2(new_n331), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n341), .A2(KEYINPUT68), .ZN(new_n361));
  INV_X1    g160(.A(new_n324), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT68), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n345), .A2(new_n363), .A3(new_n331), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n361), .A2(new_n362), .A3(KEYINPUT4), .A4(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT4), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n346), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n360), .A2(new_n349), .A3(new_n365), .A4(new_n367), .ZN(new_n368));
  AOI211_X1 g167(.A(KEYINPUT5), .B(new_n350), .C1(new_n358), .C2(new_n359), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n346), .A2(new_n366), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n361), .A2(new_n362), .A3(new_n364), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n370), .B1(new_n371), .B2(new_n366), .ZN(new_n372));
  AOI22_X1  g171(.A1(new_n353), .A2(new_n368), .B1(new_n369), .B2(new_n372), .ZN(new_n373));
  XOR2_X1   g172(.A(G1gat), .B(G29gat), .Z(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(G57gat), .B(G85gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n376), .B(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT79), .B1(new_n373), .B2(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n373), .A2(new_n378), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n307), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n353), .A2(new_n368), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n369), .A2(new_n372), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n382), .A2(KEYINPUT79), .A3(new_n383), .A4(new_n378), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n307), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n382), .A2(new_n383), .ZN(new_n386));
  INV_X1    g185(.A(new_n378), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n381), .A2(new_n389), .B1(new_n277), .B2(new_n205), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n299), .A2(new_n302), .A3(new_n306), .A4(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n274), .B1(new_n354), .B2(new_n357), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n283), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n216), .ZN(new_n394));
  OR2_X1    g193(.A1(new_n394), .A2(KEYINPUT29), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n362), .B1(new_n395), .B2(new_n356), .ZN(new_n396));
  OAI211_X1 g195(.A(G228gat), .B(G233gat), .C1(new_n393), .C2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(G22gat), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n356), .B1(new_n394), .B2(new_n274), .ZN(new_n399));
  AOI22_X1  g198(.A1(new_n399), .A2(new_n324), .B1(G228gat), .B2(G233gat), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n400), .B1(new_n392), .B2(new_n283), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n397), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n398), .B1(new_n397), .B2(new_n401), .ZN(new_n404));
  XNOR2_X1  g203(.A(G78gat), .B(G106gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT31), .B(G50gat), .ZN(new_n406));
  XOR2_X1   g205(.A(new_n405), .B(new_n406), .Z(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  OAI22_X1  g207(.A1(new_n403), .A2(new_n404), .B1(KEYINPUT82), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n404), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n407), .B(KEYINPUT82), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n410), .A2(new_n402), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n348), .A2(new_n351), .ZN(new_n415));
  OAI21_X1  g214(.A(KEYINPUT39), .B1(new_n415), .B2(new_n350), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n349), .B1(new_n372), .B2(new_n360), .ZN(new_n417));
  OR2_X1    g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT39), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n418), .A2(new_n378), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT84), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT40), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NOR2_X1   g223(.A1(KEYINPUT84), .A2(KEYINPUT40), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  NOR3_X1   g225(.A1(new_n424), .A2(new_n380), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT83), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT74), .B1(new_n277), .B2(new_n205), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT74), .ZN(new_n430));
  INV_X1    g229(.A(new_n205), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n293), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n284), .A2(new_n292), .A3(new_n205), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT30), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT30), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n284), .A2(new_n436), .A3(new_n292), .A4(new_n205), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n428), .B1(new_n433), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n433), .A2(new_n428), .A3(new_n438), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n427), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n391), .A2(new_n414), .A3(new_n443), .ZN(new_n444));
  AOI22_X1  g243(.A1(new_n429), .A2(new_n432), .B1(new_n435), .B2(new_n437), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n381), .A2(new_n445), .A3(new_n389), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT81), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT81), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n381), .A2(new_n445), .A3(new_n389), .A4(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n414), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(G227gat), .A2(G233gat), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n361), .A2(new_n364), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n290), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n272), .A2(new_n452), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n451), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT32), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OR2_X1    g257(.A1(new_n456), .A2(KEYINPUT33), .ZN(new_n459));
  XOR2_X1   g258(.A(G15gat), .B(G43gat), .Z(new_n460));
  XNOR2_X1  g259(.A(new_n460), .B(KEYINPUT69), .ZN(new_n461));
  XOR2_X1   g260(.A(G71gat), .B(G99gat), .Z(new_n462));
  XNOR2_X1  g261(.A(new_n462), .B(KEYINPUT70), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n461), .B(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n458), .A2(new_n459), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n454), .A2(new_n455), .A3(new_n451), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT34), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(KEYINPUT71), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n467), .B1(new_n466), .B2(KEYINPUT71), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n455), .ZN(new_n472));
  INV_X1    g271(.A(new_n451), .ZN(new_n473));
  AOI221_X4 g272(.A(new_n457), .B1(KEYINPUT33), .B2(new_n464), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n465), .A2(new_n471), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n470), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(new_n468), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n464), .B1(new_n456), .B2(KEYINPUT33), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n456), .A2(new_n457), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n478), .B1(new_n481), .B2(new_n474), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n476), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT36), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n476), .A2(new_n482), .A3(KEYINPUT36), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n450), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n382), .A2(new_n378), .A3(new_n383), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT79), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n388), .ZN(new_n492));
  AOI22_X1  g291(.A1(new_n492), .A2(new_n307), .B1(new_n388), .B2(new_n385), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n493), .B1(new_n441), .B2(new_n439), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT88), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n493), .B(KEYINPUT88), .C1(new_n441), .C2(new_n439), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT35), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n483), .A2(new_n498), .A3(new_n414), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n496), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n476), .A2(new_n482), .B1(new_n409), .B2(new_n413), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n447), .A2(new_n449), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT35), .ZN(new_n503));
  AOI22_X1  g302(.A1(new_n444), .A2(new_n488), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  XOR2_X1   g303(.A(KEYINPUT89), .B(KEYINPUT11), .Z(new_n505));
  XNOR2_X1  g304(.A(new_n505), .B(KEYINPUT90), .ZN(new_n506));
  XOR2_X1   g305(.A(G113gat), .B(G141gat), .Z(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  XOR2_X1   g307(.A(G169gat), .B(G197gat), .Z(new_n509));
  XNOR2_X1  g308(.A(new_n508), .B(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(KEYINPUT12), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(G229gat), .A2(G233gat), .ZN(new_n513));
  XOR2_X1   g312(.A(new_n513), .B(KEYINPUT13), .Z(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(KEYINPUT14), .B(G29gat), .ZN(new_n516));
  INV_X1    g315(.A(G36gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(G29gat), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n519), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(G43gat), .B(G50gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT15), .ZN(new_n523));
  OR2_X1    g322(.A1(new_n522), .A2(KEYINPUT15), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n521), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  OR2_X1    g324(.A1(new_n525), .A2(KEYINPUT91), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(KEYINPUT91), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n521), .A2(new_n523), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G15gat), .B(G22gat), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT92), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(G1gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n530), .A2(new_n531), .A3(G1gat), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT16), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n530), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n534), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(G8gat), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n529), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n529), .A2(new_n539), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n515), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT93), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI211_X1 g343(.A(KEYINPUT93), .B(new_n515), .C1(new_n540), .C2(new_n541), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n529), .A2(KEYINPUT17), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT17), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n526), .A2(new_n547), .A3(new_n527), .A4(new_n528), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n539), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n513), .ZN(new_n550));
  INV_X1    g349(.A(new_n541), .ZN(new_n551));
  NOR3_X1   g350(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  OAI22_X1  g351(.A1(new_n544), .A2(new_n545), .B1(new_n552), .B2(KEYINPUT18), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n546), .A2(new_n548), .ZN(new_n554));
  INV_X1    g353(.A(new_n539), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n556), .A2(new_n513), .A3(new_n541), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT18), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n512), .B1(new_n553), .B2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n542), .B(new_n543), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n552), .A2(KEYINPUT18), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n557), .A2(new_n558), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n561), .A2(new_n511), .A3(new_n562), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n504), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT94), .B1(G71gat), .B2(G78gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(G57gat), .B(G64gat), .ZN(new_n569));
  AOI21_X1  g368(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G71gat), .B(G78gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT95), .B(KEYINPUT21), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G127gat), .B(G155gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n573), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n539), .B1(KEYINPUT21), .B2(new_n578), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n577), .A2(new_n579), .ZN(new_n581));
  NAND2_X1  g380(.A1(G231gat), .A2(G233gat), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n582), .B(KEYINPUT97), .Z(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT96), .ZN(new_n584));
  XNOR2_X1  g383(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(G183gat), .B(G211gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  AND3_X1   g387(.A1(new_n580), .A2(new_n581), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n588), .B1(new_n580), .B2(new_n581), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AND2_X1   g390(.A1(G232gat), .A2(G233gat), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n592), .A2(KEYINPUT41), .ZN(new_n593));
  XNOR2_X1  g392(.A(G134gat), .B(G162gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G99gat), .B(G106gat), .ZN(new_n597));
  INV_X1    g396(.A(G99gat), .ZN(new_n598));
  INV_X1    g397(.A(G106gat), .ZN(new_n599));
  OAI21_X1  g398(.A(KEYINPUT8), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(KEYINPUT99), .B(G92gat), .Z(new_n601));
  OAI221_X1 g400(.A(new_n600), .B1(new_n597), .B2(KEYINPUT100), .C1(new_n601), .C2(G85gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(G85gat), .A2(G92gat), .ZN(new_n603));
  OAI21_X1  g402(.A(KEYINPUT7), .B1(new_n603), .B2(KEYINPUT98), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT98), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n605), .B1(G85gat), .B2(G92gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n604), .B(new_n606), .ZN(new_n607));
  OAI211_X1 g406(.A(KEYINPUT100), .B(new_n597), .C1(new_n602), .C2(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n602), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n597), .A2(KEYINPUT100), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n554), .A2(new_n608), .A3(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(G190gat), .B(G218gat), .Z(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n611), .A2(new_n608), .ZN(new_n615));
  AOI22_X1  g414(.A1(new_n529), .A2(new_n615), .B1(KEYINPUT41), .B2(new_n592), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n612), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n614), .B1(new_n612), .B2(new_n616), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n596), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n619), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n621), .A2(new_n595), .A3(new_n617), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n591), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G120gat), .B(G148gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT102), .ZN(new_n625));
  XNOR2_X1  g424(.A(G176gat), .B(G204gat), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n625), .B(new_n626), .Z(new_n627));
  NAND2_X1  g426(.A1(new_n615), .A2(new_n578), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n611), .A2(new_n573), .A3(new_n608), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G230gat), .A2(G233gat), .ZN(new_n631));
  OAI21_X1  g430(.A(KEYINPUT101), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n631), .B1(new_n628), .B2(new_n629), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT101), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n631), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT10), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n628), .A2(new_n638), .A3(new_n629), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n615), .A2(KEYINPUT10), .A3(new_n578), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n627), .B1(new_n636), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n639), .A2(new_n640), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n631), .ZN(new_n644));
  INV_X1    g443(.A(new_n627), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n644), .A2(new_n632), .A3(new_n645), .A4(new_n635), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT103), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n642), .A2(new_n646), .A3(KEYINPUT103), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n623), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT104), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n623), .A2(new_n649), .A3(KEYINPUT104), .A4(new_n650), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n567), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n656), .A2(new_n493), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(new_n533), .ZN(G1324gat));
  INV_X1    g457(.A(G8gat), .ZN(new_n659));
  INV_X1    g458(.A(new_n656), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n442), .A2(new_n440), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n659), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT16), .B(G8gat), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n656), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(KEYINPUT42), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n666), .B1(KEYINPUT42), .B2(new_n665), .ZN(G1325gat));
  INV_X1    g466(.A(new_n487), .ZN(new_n668));
  OAI21_X1  g467(.A(G15gat), .B1(new_n656), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(G15gat), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n483), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n669), .B1(new_n656), .B2(new_n671), .ZN(G1326gat));
  OR3_X1    g471(.A1(new_n656), .A2(KEYINPUT105), .A3(new_n414), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT105), .B1(new_n656), .B2(new_n414), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(KEYINPUT43), .B(G22gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1327gat));
  NAND2_X1  g476(.A1(new_n649), .A2(new_n650), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(new_n591), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n680), .A2(new_n566), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n444), .A2(new_n488), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n500), .A2(KEYINPUT107), .A3(new_n503), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT107), .B1(new_n500), .B2(new_n503), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n683), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n620), .A2(new_n622), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(KEYINPUT44), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT44), .B1(new_n504), .B2(new_n687), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n682), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(G29gat), .B1(new_n692), .B2(new_n493), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n504), .A2(new_n682), .A3(new_n687), .ZN(new_n694));
  INV_X1    g493(.A(new_n493), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n694), .A2(new_n519), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n696), .A2(new_n697), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n693), .A2(new_n698), .A3(new_n699), .ZN(G1328gat));
  NOR2_X1   g499(.A1(new_n661), .A2(G36gat), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n694), .A2(new_n701), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n702), .A2(KEYINPUT108), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n702), .A2(KEYINPUT108), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT46), .ZN(new_n705));
  OR3_X1    g504(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(G36gat), .B1(new_n692), .B2(new_n661), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n705), .B1(new_n703), .B2(new_n704), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(G1329gat));
  INV_X1    g508(.A(KEYINPUT47), .ZN(new_n710));
  INV_X1    g509(.A(G43gat), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n711), .B1(new_n691), .B2(new_n487), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n500), .A2(new_n503), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n683), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n687), .ZN(new_n715));
  AOI21_X1  g514(.A(G43gat), .B1(new_n476), .B2(new_n482), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n714), .A2(new_n715), .A3(new_n681), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT109), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n710), .B1(new_n712), .B2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n688), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT107), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n713), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n500), .A2(KEYINPUT107), .A3(new_n503), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n720), .B1(new_n724), .B2(new_n683), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n726), .B1(new_n714), .B2(new_n715), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n487), .B(new_n681), .C1(new_n725), .C2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT110), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n691), .A2(KEYINPUT110), .A3(new_n487), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n730), .A2(new_n731), .A3(G43gat), .ZN(new_n732));
  OR2_X1    g531(.A1(new_n718), .A2(new_n710), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n719), .B1(new_n732), .B2(new_n733), .ZN(G1330gat));
  INV_X1    g533(.A(G50gat), .ZN(new_n735));
  INV_X1    g534(.A(new_n414), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n735), .B1(new_n691), .B2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT111), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n414), .A2(new_n739), .A3(G50gat), .ZN(new_n740));
  AOI21_X1  g539(.A(KEYINPUT111), .B1(new_n736), .B2(new_n735), .ZN(new_n741));
  NOR4_X1   g540(.A1(new_n680), .A2(new_n687), .A3(new_n740), .A4(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n567), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n738), .A2(KEYINPUT48), .A3(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT48), .ZN(new_n745));
  INV_X1    g544(.A(new_n743), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(new_n737), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n744), .A2(new_n747), .ZN(G1331gat));
  NAND3_X1  g547(.A1(new_n678), .A2(new_n566), .A3(new_n623), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n749), .B1(new_n724), .B2(new_n683), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n695), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g551(.A(new_n661), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  OR2_X1    g553(.A1(new_n754), .A2(KEYINPUT112), .ZN(new_n755));
  NOR2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(KEYINPUT112), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n755), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n756), .B1(new_n755), .B2(new_n757), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n758), .A2(new_n759), .ZN(G1333gat));
  NAND2_X1  g559(.A1(new_n750), .A2(new_n487), .ZN(new_n761));
  AOI21_X1  g560(.A(G71gat), .B1(new_n476), .B2(new_n482), .ZN(new_n762));
  AOI22_X1  g561(.A1(new_n761), .A2(G71gat), .B1(new_n750), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g563(.A1(new_n750), .A2(new_n736), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G78gat), .ZN(G1335gat));
  INV_X1    g565(.A(new_n591), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n565), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n769), .A2(new_n679), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(new_n725), .B2(new_n727), .ZN(new_n771));
  OAI21_X1  g570(.A(G85gat), .B1(new_n771), .B2(new_n493), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n769), .A2(new_n687), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n686), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n686), .A2(KEYINPUT51), .A3(new_n773), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  OR3_X1    g578(.A1(new_n679), .A2(G85gat), .A3(new_n493), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n772), .B1(new_n779), .B2(new_n780), .ZN(G1336gat));
  INV_X1    g580(.A(KEYINPUT113), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n782), .A2(KEYINPUT52), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(KEYINPUT52), .ZN(new_n784));
  INV_X1    g583(.A(new_n601), .ZN(new_n785));
  INV_X1    g584(.A(new_n770), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n786), .B1(new_n689), .B2(new_n690), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n785), .B1(new_n787), .B2(new_n662), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n679), .A2(new_n661), .A3(G92gat), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n790), .B1(new_n776), .B2(new_n777), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n783), .B(new_n784), .C1(new_n788), .C2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n601), .B1(new_n771), .B2(new_n661), .ZN(new_n793));
  INV_X1    g592(.A(new_n777), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT51), .B1(new_n686), .B2(new_n773), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n789), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n793), .A2(new_n796), .A3(new_n782), .A4(KEYINPUT52), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n792), .A2(new_n797), .ZN(G1337gat));
  OAI21_X1  g597(.A(G99gat), .B1(new_n771), .B2(new_n668), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n678), .A2(new_n598), .A3(new_n483), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n799), .B1(new_n779), .B2(new_n800), .ZN(G1338gat));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n679), .A2(G106gat), .A3(new_n414), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n802), .B1(new_n779), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n599), .B1(new_n787), .B2(new_n736), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n787), .A2(new_n736), .ZN(new_n807));
  XOR2_X1   g606(.A(new_n803), .B(KEYINPUT114), .Z(new_n808));
  AOI22_X1  g607(.A1(new_n807), .A2(G106gat), .B1(new_n778), .B2(new_n808), .ZN(new_n809));
  OAI22_X1  g608(.A1(new_n805), .A2(new_n806), .B1(new_n809), .B2(new_n802), .ZN(G1339gat));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n679), .A2(new_n811), .A3(new_n566), .A4(new_n623), .ZN(new_n812));
  OAI21_X1  g611(.A(KEYINPUT115), .B1(new_n651), .B2(new_n565), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n550), .B1(new_n549), .B2(new_n551), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n540), .A2(new_n541), .A3(new_n515), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT117), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n817), .A2(new_n818), .A3(new_n510), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n510), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT117), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n564), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n639), .A2(new_n637), .A3(new_n640), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT116), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n823), .B(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n641), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n627), .B1(new_n644), .B2(KEYINPUT54), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n646), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n829), .B1(new_n825), .B2(new_n827), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n834), .B1(new_n835), .B2(KEYINPUT55), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n822), .A2(new_n833), .A3(new_n836), .A4(new_n715), .ZN(new_n837));
  AOI22_X1  g636(.A1(new_n831), .A2(new_n832), .B1(new_n560), .B2(new_n564), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n836), .A2(new_n838), .B1(new_n678), .B2(new_n822), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n837), .B1(new_n839), .B2(new_n715), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n814), .B1(new_n840), .B2(new_n591), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(new_n736), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n842), .A2(new_n695), .A3(new_n483), .A4(new_n661), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n843), .A2(new_n333), .A3(new_n566), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n678), .A2(new_n822), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n833), .A2(new_n836), .A3(new_n565), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n715), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n837), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n591), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n812), .A2(new_n813), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n851), .A2(new_n695), .A3(new_n501), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT118), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n662), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n841), .A2(new_n493), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(KEYINPUT118), .A3(new_n501), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n565), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n844), .B1(new_n859), .B2(new_n333), .ZN(G1340gat));
  NOR3_X1   g659(.A1(new_n843), .A2(new_n336), .A3(new_n679), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n858), .A2(new_n678), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n861), .B1(new_n862), .B2(new_n336), .ZN(G1341gat));
  OAI21_X1  g662(.A(G127gat), .B1(new_n843), .B2(new_n591), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n767), .A2(new_n327), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n864), .B1(new_n857), .B2(new_n865), .ZN(G1342gat));
  NOR2_X1   g665(.A1(new_n687), .A2(G134gat), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  OR3_X1    g667(.A1(new_n857), .A2(KEYINPUT56), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(G134gat), .B1(new_n843), .B2(new_n687), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT56), .B1(new_n857), .B2(new_n868), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(G1343gat));
  NAND2_X1  g671(.A1(new_n668), .A2(new_n736), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n873), .A2(new_n662), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n855), .A2(new_n874), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n875), .A2(G141gat), .A3(new_n566), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT58), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n661), .A2(new_n695), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n879), .A2(new_n487), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT57), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n882), .B1(new_n841), .B2(new_n414), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n851), .A2(KEYINPUT57), .A3(new_n736), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n885), .A2(new_n565), .ZN(new_n886));
  INV_X1    g685(.A(G141gat), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n877), .B(new_n878), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n887), .B1(new_n885), .B2(new_n565), .ZN(new_n889));
  OAI21_X1  g688(.A(KEYINPUT58), .B1(new_n889), .B2(new_n876), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n890), .ZN(G1344gat));
  INV_X1    g690(.A(new_n875), .ZN(new_n892));
  INV_X1    g691(.A(G148gat), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(new_n893), .A3(new_n678), .ZN(new_n894));
  XNOR2_X1  g693(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n880), .A2(new_n678), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n653), .A2(new_n566), .A3(new_n654), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n897), .B1(new_n840), .B2(new_n591), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n882), .B1(new_n898), .B2(new_n414), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n896), .B1(new_n899), .B2(new_n884), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT120), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n893), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(new_n897), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n849), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT57), .B1(new_n904), .B2(new_n736), .ZN(new_n905));
  AOI211_X1 g704(.A(new_n882), .B(new_n414), .C1(new_n849), .C2(new_n850), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(KEYINPUT120), .B1(new_n907), .B2(new_n896), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n895), .B1(new_n902), .B2(new_n908), .ZN(new_n909));
  AOI211_X1 g708(.A(KEYINPUT59), .B(new_n893), .C1(new_n885), .C2(new_n678), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n894), .B1(new_n909), .B2(new_n910), .ZN(G1345gat));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n767), .A2(new_n319), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n875), .A2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n885), .A2(new_n767), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n912), .B(new_n915), .C1(new_n916), .C2(new_n319), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n319), .B1(new_n885), .B2(new_n767), .ZN(new_n918));
  OAI21_X1  g717(.A(KEYINPUT121), .B1(new_n918), .B2(new_n914), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(G1346gat));
  NAND3_X1  g719(.A1(new_n892), .A2(new_n320), .A3(new_n715), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n885), .A2(new_n715), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(KEYINPUT122), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(G162gat), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n922), .A2(KEYINPUT122), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n921), .B1(new_n924), .B2(new_n925), .ZN(G1347gat));
  NOR2_X1   g725(.A1(new_n661), .A2(new_n695), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n483), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT124), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n842), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(G169gat), .B1(new_n930), .B2(new_n566), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n851), .A2(new_n493), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n662), .A2(new_n501), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n566), .A2(G169gat), .ZN(new_n935));
  AOI21_X1  g734(.A(KEYINPUT123), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT123), .ZN(new_n937));
  INV_X1    g736(.A(new_n935), .ZN(new_n938));
  NOR4_X1   g737(.A1(new_n932), .A2(new_n937), .A3(new_n933), .A4(new_n938), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n931), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT125), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT125), .ZN(new_n942));
  OAI211_X1 g741(.A(new_n931), .B(new_n942), .C1(new_n936), .C2(new_n939), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(G1348gat));
  OAI21_X1  g743(.A(G176gat), .B1(new_n930), .B2(new_n679), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n934), .A2(new_n224), .A3(new_n678), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1349gat));
  OAI21_X1  g746(.A(G183gat), .B1(new_n930), .B2(new_n591), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n934), .A2(new_n236), .A3(new_n767), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g750(.A1(new_n934), .A2(new_n237), .A3(new_n715), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n851), .A2(new_n929), .A3(new_n414), .A4(new_n715), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT61), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n953), .A2(new_n954), .A3(G190gat), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n954), .B1(new_n953), .B2(G190gat), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n952), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT126), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n957), .B(new_n958), .ZN(G1351gat));
  NOR2_X1   g758(.A1(new_n873), .A2(new_n661), .ZN(new_n960));
  XOR2_X1   g759(.A(new_n960), .B(KEYINPUT127), .Z(new_n961));
  NOR2_X1   g760(.A1(new_n961), .A2(new_n932), .ZN(new_n962));
  AOI21_X1  g761(.A(G197gat), .B1(new_n962), .B2(new_n565), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n899), .A2(new_n884), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n487), .A2(new_n695), .A3(new_n661), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n565), .A2(G197gat), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n963), .B1(new_n966), .B2(new_n967), .ZN(G1352gat));
  NOR4_X1   g767(.A1(new_n961), .A2(new_n932), .A3(G204gat), .A4(new_n679), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n969), .B(KEYINPUT62), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n966), .A2(new_n678), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(G204gat), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n970), .A2(new_n972), .ZN(G1353gat));
  NAND3_X1  g772(.A1(new_n962), .A2(new_n208), .A3(new_n767), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n964), .A2(new_n767), .A3(new_n965), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n975), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n976));
  AOI21_X1  g775(.A(KEYINPUT63), .B1(new_n975), .B2(G211gat), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n974), .B1(new_n976), .B2(new_n977), .ZN(G1354gat));
  NAND3_X1  g777(.A1(new_n962), .A2(new_n209), .A3(new_n715), .ZN(new_n979));
  AND2_X1   g778(.A1(new_n966), .A2(new_n715), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n979), .B1(new_n980), .B2(new_n209), .ZN(G1355gat));
endmodule


