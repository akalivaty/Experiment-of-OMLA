//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 1 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 0 0 0 1 0 1 1 1 0 1 1 1 0 1 0 1 0 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n775, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n851, new_n852, new_n854, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964;
  NOR2_X1   g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT80), .ZN(new_n204));
  NAND2_X1  g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n205), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT80), .B1(new_n207), .B2(new_n202), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT2), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n206), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  XOR2_X1   g009(.A(G155gat), .B(G162gat), .Z(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n203), .A2(new_n205), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT81), .B(G162gat), .ZN(new_n215));
  INV_X1    g014(.A(G155gat), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT2), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n212), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G120gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G113gat), .ZN(new_n221));
  INV_X1    g020(.A(G113gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G120gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G127gat), .ZN(new_n227));
  INV_X1    g026(.A(G134gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G127gat), .A2(G134gat), .ZN(new_n230));
  AOI22_X1  g029(.A1(new_n229), .A2(new_n230), .B1(KEYINPUT70), .B2(new_n225), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n226), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n225), .A2(KEYINPUT70), .ZN(new_n233));
  INV_X1    g032(.A(new_n230), .ZN(new_n234));
  NOR2_X1   g033(.A1(G127gat), .A2(G134gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n236), .A2(new_n225), .A3(new_n224), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n232), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n219), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G225gat), .A2(G233gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n238), .A2(new_n212), .A3(new_n218), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  AND3_X1   g042(.A1(new_n243), .A2(KEYINPUT86), .A3(KEYINPUT39), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n238), .B1(new_n219), .B2(KEYINPUT3), .ZN(new_n245));
  AOI22_X1  g044(.A1(new_n210), .A2(new_n211), .B1(new_n214), .B2(new_n217), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n242), .A2(KEYINPUT4), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT4), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n238), .A2(new_n212), .A3(new_n251), .A4(new_n218), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n241), .B1(new_n249), .B2(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT86), .B1(new_n243), .B2(KEYINPUT39), .ZN(new_n255));
  NOR3_X1   g054(.A1(new_n244), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  AOI211_X1 g056(.A(KEYINPUT39), .B(new_n241), .C1(new_n249), .C2(new_n253), .ZN(new_n258));
  XNOR2_X1  g057(.A(G1gat), .B(G29gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(KEYINPUT0), .ZN(new_n260));
  XNOR2_X1  g059(.A(G57gat), .B(G85gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(KEYINPUT84), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NOR3_X1   g063(.A1(new_n258), .A2(new_n264), .A3(KEYINPUT85), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT85), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT39), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n254), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n266), .B1(new_n268), .B2(new_n263), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n257), .B1(new_n265), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT87), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT40), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT85), .B1(new_n258), .B2(new_n264), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n268), .A2(new_n266), .A3(new_n263), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n256), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT87), .B1(new_n276), .B2(KEYINPUT40), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G8gat), .B(G36gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(G64gat), .B(G92gat), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n279), .B(new_n280), .Z(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G197gat), .B(G204gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(KEYINPUT76), .B(G211gat), .ZN(new_n284));
  INV_X1    g083(.A(G218gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n283), .B1(new_n286), .B2(KEYINPUT22), .ZN(new_n287));
  XNOR2_X1  g086(.A(G211gat), .B(G218gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  OR2_X1    g089(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n291), .A2(KEYINPUT27), .A3(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n294));
  INV_X1    g093(.A(G183gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n293), .B(new_n294), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(KEYINPUT27), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT27), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G183gat), .ZN(new_n300));
  INV_X1    g099(.A(G190gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n298), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  AOI22_X1  g101(.A1(new_n302), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n297), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT64), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT64), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n307), .A2(G169gat), .A3(G176gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT69), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT68), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT68), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n313), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n309), .A2(new_n310), .A3(new_n312), .A4(new_n314), .ZN(new_n315));
  OR3_X1    g114(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n309), .A2(new_n312), .A3(new_n314), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT69), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n304), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n291), .A2(new_n301), .A3(new_n292), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT66), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G183gat), .A2(G190gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT24), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT24), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n326), .A2(G183gat), .A3(G190gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n291), .A2(KEYINPUT66), .A3(new_n301), .A4(new_n292), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n323), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT23), .ZN(new_n331));
  INV_X1    g130(.A(G169gat), .ZN(new_n332));
  INV_X1    g131(.A(G176gat), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AND3_X1   g135(.A1(new_n336), .A2(new_n309), .A3(KEYINPUT25), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n295), .A2(new_n301), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n328), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n339), .A2(new_n309), .A3(new_n336), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT25), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n330), .A2(new_n337), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n320), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(G226gat), .A2(G233gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT77), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n346), .B1(new_n320), .B2(new_n342), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT29), .ZN(new_n348));
  INV_X1    g147(.A(new_n311), .ZN(new_n349));
  AOI22_X1  g148(.A1(new_n349), .A2(new_n313), .B1(new_n306), .B2(new_n308), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n310), .B1(new_n350), .B2(new_n312), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n315), .A2(new_n316), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n297), .B(new_n303), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n330), .A2(new_n337), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n340), .A2(new_n341), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n353), .A2(new_n356), .A3(KEYINPUT77), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n347), .A2(new_n348), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(new_n344), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n345), .B1(new_n359), .B2(KEYINPUT78), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT78), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n358), .A2(new_n361), .A3(new_n344), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n290), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n344), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n347), .A2(new_n364), .A3(new_n357), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n344), .B1(new_n343), .B2(KEYINPUT29), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT79), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n347), .A2(new_n357), .A3(KEYINPUT79), .A4(new_n364), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n289), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n282), .B1(new_n363), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n370), .ZN(new_n372));
  AND3_X1   g171(.A1(new_n358), .A2(new_n361), .A3(new_n344), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n361), .B1(new_n358), .B2(new_n344), .ZN(new_n374));
  NOR3_X1   g173(.A1(new_n373), .A2(new_n374), .A3(new_n345), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n372), .B(new_n281), .C1(new_n375), .C2(new_n290), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n371), .A2(new_n376), .A3(KEYINPUT30), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n359), .A2(KEYINPUT78), .ZN(new_n378));
  INV_X1    g177(.A(new_n345), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n378), .A2(new_n362), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n370), .B1(new_n380), .B2(new_n289), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT30), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n381), .A2(new_n382), .A3(new_n281), .ZN(new_n383));
  INV_X1    g182(.A(new_n241), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n384), .B1(new_n245), .B2(new_n248), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n252), .A2(KEYINPUT82), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT82), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n246), .A2(new_n387), .A3(new_n251), .A4(new_n238), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n386), .A2(new_n388), .A3(new_n250), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT5), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n240), .A2(new_n242), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n391), .B1(new_n392), .B2(new_n384), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT5), .B1(new_n250), .B2(new_n252), .ZN(new_n394));
  AOI22_X1  g193(.A1(new_n390), .A2(new_n393), .B1(new_n385), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT88), .B1(new_n395), .B2(new_n263), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT88), .ZN(new_n397));
  INV_X1    g196(.A(new_n242), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n238), .B1(new_n212), .B2(new_n218), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n384), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT5), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n401), .B1(new_n385), .B2(new_n389), .ZN(new_n402));
  AND2_X1   g201(.A1(new_n385), .A2(new_n394), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n397), .B(new_n264), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n276), .A2(KEYINPUT40), .B1(new_n396), .B2(new_n404), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n278), .A2(new_n377), .A3(new_n383), .A4(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n248), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n289), .B1(new_n407), .B2(KEYINPUT29), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT3), .B1(new_n290), .B2(new_n348), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n408), .B1(new_n409), .B2(new_n246), .ZN(new_n410));
  XNOR2_X1  g209(.A(G78gat), .B(G106gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(G228gat), .A2(G233gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(G22gat), .ZN(new_n414));
  XOR2_X1   g213(.A(KEYINPUT31), .B(G50gat), .Z(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n412), .B(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n406), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT37), .B1(new_n363), .B2(new_n370), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n282), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT90), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT37), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n422), .B(new_n372), .C1(new_n375), .C2(new_n290), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT89), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n381), .A2(KEYINPUT89), .A3(new_n422), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT90), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n428), .B(new_n282), .C1(new_n381), .C2(new_n422), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n421), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT38), .ZN(new_n431));
  OAI211_X1 g230(.A(KEYINPUT6), .B(new_n262), .C1(new_n402), .C2(new_n403), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n396), .A2(new_n404), .ZN(new_n434));
  INV_X1    g233(.A(new_n262), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT6), .B1(new_n395), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n433), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(new_n376), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n380), .A2(new_n290), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n368), .A2(new_n369), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n422), .B1(new_n440), .B2(new_n289), .ZN(new_n441));
  AOI211_X1 g240(.A(KEYINPUT38), .B(new_n281), .C1(new_n439), .C2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n438), .B1(new_n427), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n418), .B1(new_n431), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT71), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n238), .B1(new_n320), .B2(new_n342), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n353), .A2(new_n356), .A3(new_n239), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(G227gat), .ZN(new_n449));
  INV_X1    g248(.A(G233gat), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n445), .B1(new_n448), .B2(new_n452), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n446), .A2(new_n447), .A3(KEYINPUT71), .A4(new_n451), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT33), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n453), .A2(new_n454), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT32), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT73), .ZN(new_n459));
  XNOR2_X1  g258(.A(G15gat), .B(G43gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n460), .B(KEYINPUT72), .ZN(new_n461));
  XNOR2_X1  g260(.A(G71gat), .B(G99gat), .ZN(new_n462));
  XOR2_X1   g261(.A(new_n461), .B(new_n462), .Z(new_n463));
  NAND4_X1  g262(.A1(new_n456), .A2(new_n458), .A3(new_n459), .A4(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT75), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT32), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n466), .B1(new_n453), .B2(new_n454), .ZN(new_n467));
  INV_X1    g266(.A(new_n463), .ZN(new_n468));
  NOR3_X1   g267(.A1(new_n455), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n463), .A2(KEYINPUT33), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n457), .A2(KEYINPUT32), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT73), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n464), .B(new_n465), .C1(new_n469), .C2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT34), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n448), .A2(new_n474), .A3(new_n452), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT74), .ZN(new_n476));
  OR2_X1    g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n448), .A2(new_n452), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT34), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n475), .A2(new_n476), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n477), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n473), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n456), .A2(new_n458), .A3(new_n463), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n483), .A2(KEYINPUT73), .A3(new_n471), .ZN(new_n484));
  INV_X1    g283(.A(new_n481), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n484), .A2(new_n465), .A3(new_n464), .A4(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n482), .A2(new_n486), .A3(KEYINPUT36), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n464), .B1(new_n469), .B2(new_n472), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(new_n485), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT36), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n464), .B(new_n481), .C1(new_n469), .C2(new_n472), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT83), .B1(new_n395), .B2(new_n435), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT83), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n494), .B(new_n262), .C1(new_n402), .C2(new_n403), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n493), .A2(new_n436), .A3(new_n495), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n496), .A2(new_n432), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n497), .B1(new_n377), .B2(new_n383), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n487), .B(new_n492), .C1(new_n417), .C2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT91), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n377), .A2(new_n383), .ZN(new_n501));
  INV_X1    g300(.A(new_n437), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AOI211_X1 g302(.A(KEYINPUT91), .B(new_n437), .C1(new_n377), .C2(new_n383), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT35), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n489), .A2(new_n505), .A3(new_n417), .A4(new_n491), .ZN(new_n506));
  NOR3_X1   g305(.A1(new_n503), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n417), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n508), .B1(new_n482), .B2(new_n486), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n505), .B1(new_n509), .B2(new_n498), .ZN(new_n510));
  OAI22_X1  g309(.A1(new_n444), .A2(new_n499), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(G8gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(G15gat), .B(G22gat), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT16), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n513), .B1(new_n514), .B2(G1gat), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n512), .B1(new_n515), .B2(KEYINPUT95), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n515), .B1(G1gat), .B2(new_n513), .ZN(new_n517));
  OR2_X1    g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n517), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(G29gat), .A2(G36gat), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT14), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n522), .B(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(G29gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(KEYINPUT94), .B(G36gat), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT15), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n524), .B(KEYINPUT15), .C1(new_n525), .C2(new_n526), .ZN(new_n530));
  XNOR2_X1  g329(.A(G43gat), .B(G50gat), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  OR2_X1    g331(.A1(new_n530), .A2(new_n531), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n534), .A2(KEYINPUT17), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT17), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n536), .B1(new_n532), .B2(new_n533), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n521), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(G229gat), .A2(G233gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n534), .A2(new_n520), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT96), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT18), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n543), .B1(new_n542), .B2(new_n541), .ZN(new_n544));
  INV_X1    g343(.A(new_n540), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n534), .B(KEYINPUT17), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n545), .B1(new_n546), .B2(new_n521), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n547), .A2(KEYINPUT97), .A3(KEYINPUT18), .A4(new_n539), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT97), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT18), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n549), .B1(new_n541), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n534), .B(new_n520), .ZN(new_n553));
  XNOR2_X1  g352(.A(KEYINPUT98), .B(KEYINPUT13), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(new_n539), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n544), .A2(new_n552), .A3(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G113gat), .B(G141gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(G169gat), .B(G197gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(KEYINPUT93), .B(KEYINPUT12), .Z(new_n563));
  XOR2_X1   g362(.A(new_n562), .B(new_n563), .Z(new_n564));
  NAND2_X1  g363(.A1(new_n557), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n564), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n544), .A2(new_n552), .A3(new_n566), .A4(new_n556), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n565), .A2(KEYINPUT99), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT99), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n557), .A2(new_n569), .A3(new_n564), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  AND2_X1   g371(.A1(G71gat), .A2(G78gat), .ZN(new_n573));
  NOR2_X1   g372(.A1(G71gat), .A2(G78gat), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  XOR2_X1   g374(.A(G57gat), .B(G64gat), .Z(new_n576));
  AOI21_X1  g375(.A(new_n575), .B1(new_n576), .B2(KEYINPUT100), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n576), .B1(KEYINPUT9), .B2(new_n573), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI221_X1 g378(.A(new_n576), .B1(KEYINPUT9), .B2(new_n573), .C1(new_n575), .C2(KEYINPUT100), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n520), .B1(KEYINPUT21), .B2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT102), .B(KEYINPUT20), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n581), .A2(KEYINPUT21), .ZN(new_n586));
  NAND2_X1  g385(.A1(G231gat), .A2(G233gat), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n586), .B(new_n587), .Z(new_n588));
  XNOR2_X1  g387(.A(KEYINPUT101), .B(KEYINPUT19), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n588), .A2(new_n589), .ZN(new_n591));
  XNOR2_X1  g390(.A(G127gat), .B(G155gat), .ZN(new_n592));
  OR3_X1    g391(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n592), .B1(new_n590), .B2(new_n591), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G183gat), .B(G211gat), .Z(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n595), .A2(new_n596), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n585), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n599), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n601), .A2(new_n584), .A3(new_n597), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G232gat), .A2(G233gat), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n604), .B(KEYINPUT103), .Z(new_n605));
  INV_X1    g404(.A(KEYINPUT41), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G85gat), .A2(G92gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT7), .ZN(new_n609));
  OR2_X1    g408(.A1(G99gat), .A2(G106gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(G99gat), .A2(G106gat), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(G85gat), .ZN(new_n613));
  INV_X1    g412(.A(G92gat), .ZN(new_n614));
  AOI22_X1  g413(.A1(KEYINPUT8), .A2(new_n611), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n609), .A2(new_n612), .A3(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n616), .B(KEYINPUT104), .Z(new_n617));
  NAND2_X1  g416(.A1(new_n609), .A2(new_n615), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n618), .A2(new_n611), .A3(new_n610), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(KEYINPUT105), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n619), .A2(KEYINPUT105), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n617), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n607), .B1(new_n623), .B2(new_n534), .ZN(new_n624));
  XNOR2_X1  g423(.A(G190gat), .B(G218gat), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n535), .A2(new_n537), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n624), .B(new_n626), .C1(new_n627), .C2(new_n623), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT106), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n605), .A2(new_n606), .ZN(new_n631));
  XOR2_X1   g430(.A(G134gat), .B(G162gat), .Z(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n624), .B1(new_n627), .B2(new_n623), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n625), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n628), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n634), .A2(new_n637), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n603), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(G230gat), .A2(G233gat), .ZN(new_n644));
  AND3_X1   g443(.A1(new_n581), .A2(new_n616), .A3(new_n619), .ZN(new_n645));
  INV_X1    g444(.A(new_n581), .ZN(new_n646));
  AOI211_X1 g445(.A(KEYINPUT10), .B(new_n645), .C1(new_n622), .C2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n581), .A2(KEYINPUT10), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n622), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n644), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n645), .B1(new_n622), .B2(new_n646), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n650), .B1(new_n644), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(G120gat), .B(G148gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(G176gat), .B(G204gat), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n653), .B(new_n654), .Z(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT107), .ZN(new_n658));
  OAI211_X1 g457(.A(new_n650), .B(new_n655), .C1(new_n644), .C2(new_n651), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n652), .A2(KEYINPUT107), .A3(new_n656), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AND4_X1   g461(.A1(new_n511), .A2(new_n572), .A3(new_n643), .A4(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(new_n497), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(G1gat), .ZN(G1324gat));
  INV_X1    g464(.A(new_n501), .ZN(new_n666));
  XOR2_X1   g465(.A(KEYINPUT16), .B(G8gat), .Z(new_n667));
  AND3_X1   g466(.A1(new_n663), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n512), .B1(new_n663), .B2(new_n666), .ZN(new_n669));
  OAI21_X1  g468(.A(KEYINPUT42), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n670), .B1(KEYINPUT42), .B2(new_n668), .ZN(G1325gat));
  AND2_X1   g470(.A1(new_n489), .A2(new_n491), .ZN(new_n672));
  AOI21_X1  g471(.A(G15gat), .B1(new_n663), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n487), .A2(new_n492), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(G15gat), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n675), .B(KEYINPUT108), .Z(new_n676));
  AOI21_X1  g475(.A(new_n673), .B1(new_n663), .B2(new_n676), .ZN(G1326gat));
  NAND2_X1  g476(.A1(new_n663), .A2(new_n508), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT43), .B(G22gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1327gat));
  NAND2_X1  g479(.A1(new_n511), .A2(new_n642), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n572), .A2(new_n603), .A3(new_n662), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n683), .A2(new_n525), .A3(new_n497), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT45), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n406), .A2(new_n417), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT38), .ZN(new_n687));
  INV_X1    g486(.A(new_n429), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n428), .B1(new_n419), .B2(new_n282), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n687), .B1(new_n690), .B2(new_n427), .ZN(new_n691));
  INV_X1    g490(.A(new_n443), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n686), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n498), .A2(new_n417), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n674), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n501), .A2(new_n502), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(KEYINPUT91), .ZN(new_n697));
  INV_X1    g496(.A(new_n506), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n501), .A2(new_n502), .A3(new_n500), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n482), .A2(new_n486), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n701), .A2(new_n498), .A3(new_n417), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(KEYINPUT35), .ZN(new_n703));
  AOI22_X1  g502(.A1(new_n693), .A2(new_n695), .B1(new_n700), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT44), .B1(new_n704), .B2(new_n641), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT110), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n706), .B1(new_n639), .B2(new_n640), .ZN(new_n707));
  INV_X1    g506(.A(new_n640), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n708), .A2(KEYINPUT110), .A3(new_n638), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g509(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n711));
  NAND3_X1  g510(.A1(new_n511), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n682), .B1(new_n705), .B2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n497), .ZN(new_n715));
  OAI21_X1  g514(.A(G29gat), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n685), .A2(new_n716), .ZN(G1328gat));
  NAND3_X1  g516(.A1(new_n683), .A2(new_n666), .A3(new_n526), .ZN(new_n718));
  XOR2_X1   g517(.A(new_n718), .B(KEYINPUT46), .Z(new_n719));
  NOR2_X1   g518(.A1(new_n714), .A2(new_n501), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n719), .B1(new_n526), .B2(new_n720), .ZN(G1329gat));
  INV_X1    g520(.A(new_n674), .ZN(new_n722));
  OAI21_X1  g521(.A(G43gat), .B1(new_n714), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(G43gat), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n683), .A2(new_n724), .A3(new_n672), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(KEYINPUT47), .B1(new_n725), .B2(KEYINPUT111), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1330gat));
  NOR2_X1   g527(.A1(new_n417), .A2(G50gat), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n681), .A2(new_n682), .A3(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT112), .ZN(new_n733));
  AOI21_X1  g532(.A(KEYINPUT48), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT113), .ZN(new_n736));
  INV_X1    g535(.A(new_n682), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n738), .B1(new_n511), .B2(new_n642), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n710), .A2(new_n711), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n693), .A2(new_n695), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n700), .A2(new_n703), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n508), .B(new_n737), .C1(new_n739), .C2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(G50gat), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n736), .B1(new_n745), .B2(new_n732), .ZN(new_n746));
  AOI211_X1 g545(.A(KEYINPUT113), .B(new_n731), .C1(new_n744), .C2(G50gat), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n735), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(G50gat), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n749), .B1(new_n713), .B2(new_n508), .ZN(new_n750));
  OAI21_X1  g549(.A(KEYINPUT113), .B1(new_n750), .B2(new_n731), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n745), .A2(new_n732), .A3(new_n736), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n751), .A2(new_n734), .A3(new_n752), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n748), .A2(new_n753), .ZN(G1331gat));
  INV_X1    g553(.A(new_n662), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n643), .A2(new_n571), .A3(new_n755), .ZN(new_n756));
  OR3_X1    g555(.A1(new_n704), .A2(KEYINPUT114), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(KEYINPUT114), .B1(new_n704), .B2(new_n756), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n497), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g561(.A1(new_n759), .A2(new_n501), .ZN(new_n763));
  NOR2_X1   g562(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n764));
  AND2_X1   g563(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(new_n763), .B2(new_n764), .ZN(G1333gat));
  XOR2_X1   g566(.A(new_n672), .B(KEYINPUT115), .Z(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n759), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n674), .A2(G71gat), .ZN(new_n771));
  OAI22_X1  g570(.A1(new_n770), .A2(G71gat), .B1(new_n759), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(KEYINPUT116), .B(KEYINPUT50), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n772), .B(new_n773), .ZN(G1334gat));
  NAND2_X1  g573(.A1(new_n760), .A2(new_n508), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(G78gat), .ZN(G1335gat));
  INV_X1    g575(.A(new_n603), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n777), .A2(new_n572), .A3(new_n662), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n778), .B1(new_n739), .B2(new_n743), .ZN(new_n779));
  OAI21_X1  g578(.A(G85gat), .B1(new_n779), .B2(new_n715), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n511), .A2(new_n571), .A3(new_n642), .A4(new_n603), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT51), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n755), .A2(new_n613), .A3(new_n497), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n780), .B1(new_n782), .B2(new_n783), .ZN(G1336gat));
  OAI21_X1  g583(.A(G92gat), .B1(new_n779), .B2(new_n501), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n501), .A2(new_n662), .A3(G92gat), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n785), .B(new_n786), .C1(new_n782), .C2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT118), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n781), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT51), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n781), .A2(new_n791), .A3(KEYINPUT51), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n794), .A2(new_n795), .A3(new_n787), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n785), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n790), .B1(new_n797), .B2(KEYINPUT52), .ZN(new_n798));
  AOI211_X1 g597(.A(KEYINPUT118), .B(new_n786), .C1(new_n796), .C2(new_n785), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n789), .B1(new_n798), .B2(new_n799), .ZN(G1337gat));
  OAI21_X1  g599(.A(G99gat), .B1(new_n779), .B2(new_n722), .ZN(new_n801));
  INV_X1    g600(.A(G99gat), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n672), .A2(new_n802), .A3(new_n755), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n801), .B1(new_n782), .B2(new_n803), .ZN(G1338gat));
  OAI21_X1  g603(.A(G106gat), .B1(new_n779), .B2(new_n417), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n662), .A2(G106gat), .A3(new_n417), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n805), .B(new_n806), .C1(new_n782), .C2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n794), .A2(new_n795), .A3(new_n807), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n810), .A2(new_n805), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n809), .B1(new_n811), .B2(new_n806), .ZN(G1339gat));
  INV_X1    g611(.A(KEYINPUT119), .ZN(new_n813));
  INV_X1    g612(.A(new_n644), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT10), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n651), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n649), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n814), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n655), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n816), .A2(new_n814), .A3(new_n817), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n650), .A2(new_n821), .A3(KEYINPUT54), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n820), .A2(KEYINPUT55), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n659), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT55), .B1(new_n820), .B2(new_n822), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n813), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n825), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n827), .A2(KEYINPUT119), .A3(new_n659), .A4(new_n823), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n568), .A2(new_n826), .A3(new_n570), .A4(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n547), .A2(new_n539), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n553), .A2(new_n555), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n562), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n567), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n755), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n710), .B1(new_n829), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n709), .A2(new_n707), .A3(new_n833), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n826), .A2(new_n828), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n603), .B1(new_n835), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n643), .A2(new_n571), .A3(new_n662), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n715), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n841), .A2(new_n501), .A3(new_n509), .ZN(new_n842));
  AOI21_X1  g641(.A(G113gat), .B1(new_n842), .B2(new_n572), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n508), .B1(new_n839), .B2(new_n840), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n844), .A2(new_n497), .A3(new_n501), .A4(new_n672), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n845), .A2(new_n222), .A3(new_n571), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n843), .A2(new_n846), .ZN(G1340gat));
  AOI21_X1  g646(.A(G120gat), .B1(new_n842), .B2(new_n755), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n845), .A2(new_n220), .A3(new_n662), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(G1341gat));
  NAND3_X1  g649(.A1(new_n842), .A2(new_n227), .A3(new_n777), .ZN(new_n851));
  OAI21_X1  g650(.A(G127gat), .B1(new_n845), .B2(new_n603), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(G1342gat));
  NAND3_X1  g652(.A1(new_n842), .A2(new_n228), .A3(new_n642), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n854), .A2(KEYINPUT56), .ZN(new_n855));
  OAI21_X1  g654(.A(G134gat), .B1(new_n845), .B2(new_n641), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(KEYINPUT56), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(G1343gat));
  NOR3_X1   g657(.A1(new_n674), .A2(new_n666), .A3(new_n417), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n841), .A2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n571), .A2(G141gat), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(KEYINPUT120), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n839), .A2(new_n840), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n508), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(KEYINPUT57), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n674), .A2(new_n715), .A3(new_n666), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n824), .A2(new_n825), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n568), .A2(new_n570), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n642), .B1(new_n870), .B2(new_n834), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n603), .B1(new_n871), .B2(new_n838), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n417), .B1(new_n872), .B2(new_n840), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT57), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n868), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n867), .A2(new_n875), .A3(new_n571), .ZN(new_n876));
  INV_X1    g675(.A(G141gat), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n864), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n878), .B(KEYINPUT58), .ZN(G1344gat));
  NOR3_X1   g678(.A1(new_n860), .A2(G148gat), .A3(new_n662), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n880), .B(KEYINPUT121), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n868), .A2(new_n755), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n642), .A2(new_n833), .A3(new_n869), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n603), .B1(new_n871), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n417), .B1(new_n884), .B2(new_n840), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(KEYINPUT57), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n417), .B1(new_n839), .B2(new_n840), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT57), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n886), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  AOI211_X1 g689(.A(new_n874), .B(new_n417), .C1(new_n839), .C2(new_n840), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(KEYINPUT122), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n882), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n894));
  INV_X1    g693(.A(G148gat), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n867), .A2(new_n875), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n895), .B1(new_n896), .B2(new_n755), .ZN(new_n897));
  OAI221_X1 g696(.A(new_n881), .B1(new_n893), .B2(new_n894), .C1(KEYINPUT59), .C2(new_n897), .ZN(G1345gat));
  AOI21_X1  g697(.A(G155gat), .B1(new_n861), .B2(new_n777), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n603), .A2(new_n216), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT123), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n899), .B1(new_n896), .B2(new_n901), .ZN(G1346gat));
  INV_X1    g701(.A(new_n710), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n903), .A2(new_n215), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n861), .A2(new_n642), .ZN(new_n905));
  AOI22_X1  g704(.A1(new_n896), .A2(new_n904), .B1(new_n905), .B2(new_n215), .ZN(G1347gat));
  NOR2_X1   g705(.A1(new_n501), .A2(new_n497), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n865), .A2(new_n509), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(G169gat), .B1(new_n908), .B2(new_n572), .ZN(new_n909));
  INV_X1    g708(.A(new_n907), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n769), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n844), .A2(new_n911), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n912), .A2(new_n332), .A3(new_n571), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n909), .A2(new_n913), .ZN(G1348gat));
  NAND4_X1  g713(.A1(new_n844), .A2(G176gat), .A3(new_n755), .A4(new_n911), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n915), .A2(KEYINPUT124), .ZN(new_n916));
  AOI21_X1  g715(.A(G176gat), .B1(new_n908), .B2(new_n755), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n915), .A2(KEYINPUT124), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(G1349gat));
  NAND2_X1  g718(.A1(new_n291), .A2(new_n292), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n920), .B1(new_n912), .B2(new_n603), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n777), .A2(new_n298), .A3(new_n300), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n908), .A2(new_n922), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n923), .A2(KEYINPUT125), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n923), .A2(KEYINPUT125), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n921), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(KEYINPUT60), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT60), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n928), .B(new_n921), .C1(new_n924), .C2(new_n925), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n929), .ZN(G1350gat));
  NAND3_X1  g729(.A1(new_n908), .A2(new_n301), .A3(new_n710), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n844), .A2(new_n642), .A3(new_n911), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n933));
  AND3_X1   g732(.A1(new_n932), .A2(new_n933), .A3(G190gat), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n933), .B1(new_n932), .B2(G190gat), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n931), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT126), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n936), .B(new_n937), .ZN(G1351gat));
  NOR2_X1   g737(.A1(new_n674), .A2(new_n910), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n888), .A2(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(G197gat), .B1(new_n941), .B2(new_n572), .ZN(new_n942));
  INV_X1    g741(.A(new_n939), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n943), .B1(new_n890), .B2(new_n892), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n572), .A2(G197gat), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(G1352gat));
  NAND2_X1  g745(.A1(new_n944), .A2(new_n755), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(G204gat), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n940), .A2(G204gat), .A3(new_n662), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT62), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(G1353gat));
  OAI22_X1  g750(.A1(new_n891), .A2(KEYINPUT122), .B1(KEYINPUT57), .B2(new_n885), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n889), .A2(new_n887), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n777), .B(new_n939), .C1(new_n952), .C2(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(G211gat), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(KEYINPUT63), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT63), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n954), .A2(new_n957), .A3(G211gat), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n941), .A2(new_n284), .A3(new_n777), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT127), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n959), .B(new_n960), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n956), .A2(new_n958), .A3(new_n961), .ZN(G1354gat));
  NAND3_X1  g761(.A1(new_n941), .A2(new_n285), .A3(new_n710), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n944), .A2(new_n642), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n963), .B1(new_n964), .B2(new_n285), .ZN(G1355gat));
endmodule


