

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740;

  XNOR2_X1 U363 ( .A(n369), .B(n457), .ZN(n564) );
  AND2_X1 U364 ( .A1(n605), .A2(n604), .ZN(n340) );
  AND2_X1 U365 ( .A1(n591), .A2(n590), .ZN(n341) );
  AND2_X1 U366 ( .A1(n593), .A2(n592), .ZN(n342) );
  XNOR2_X2 U367 ( .A(n345), .B(n344), .ZN(n686) );
  XNOR2_X2 U368 ( .A(n543), .B(n542), .ZN(n575) );
  XNOR2_X2 U369 ( .A(n466), .B(n434), .ZN(n729) );
  XNOR2_X2 U370 ( .A(n446), .B(KEYINPUT10), .ZN(n466) );
  INV_X1 U371 ( .A(G953), .ZN(n723) );
  NAND2_X1 U372 ( .A1(n589), .A2(n363), .ZN(n594) );
  NAND2_X1 U373 ( .A1(n346), .A2(n343), .ZN(n345) );
  XNOR2_X1 U374 ( .A(n485), .B(n421), .ZN(n728) );
  INV_X1 U375 ( .A(KEYINPUT33), .ZN(n344) );
  INV_X1 U376 ( .A(KEYINPUT45), .ZN(n354) );
  XNOR2_X1 U377 ( .A(n355), .B(n354), .ZN(n716) );
  NAND2_X1 U378 ( .A1(n340), .A2(n353), .ZN(n355) );
  NAND2_X1 U379 ( .A1(n351), .A2(n350), .ZN(n353) );
  INV_X1 U380 ( .A(n342), .ZN(n352) );
  XNOR2_X1 U381 ( .A(n598), .B(n347), .ZN(n346) );
  INV_X1 U382 ( .A(n582), .ZN(n343) );
  XNOR2_X1 U383 ( .A(n443), .B(G134), .ZN(n485) );
  INV_X1 U384 ( .A(KEYINPUT102), .ZN(n347) );
  XNOR2_X1 U385 ( .A(G143), .B(G128), .ZN(n443) );
  INV_X1 U386 ( .A(KEYINPUT1), .ZN(n348) );
  INV_X1 U387 ( .A(n686), .ZN(n371) );
  INV_X1 U388 ( .A(n580), .ZN(n579) );
  XNOR2_X1 U389 ( .A(n516), .B(n348), .ZN(n580) );
  XNOR2_X2 U390 ( .A(n349), .B(n439), .ZN(n516) );
  NAND2_X1 U391 ( .A1(n642), .A2(n454), .ZN(n349) );
  NAND2_X1 U392 ( .A1(n594), .A2(n342), .ZN(n350) );
  NAND2_X1 U393 ( .A1(n341), .A2(n352), .ZN(n351) );
  INV_X1 U394 ( .A(n377), .ZN(n356) );
  XNOR2_X1 U395 ( .A(n438), .B(n379), .ZN(n357) );
  XNOR2_X1 U396 ( .A(n438), .B(n379), .ZN(n642) );
  INV_X1 U397 ( .A(n739), .ZN(n388) );
  XNOR2_X1 U398 ( .A(n426), .B(n366), .ZN(n442) );
  XNOR2_X1 U399 ( .A(G116), .B(G113), .ZN(n426) );
  XNOR2_X1 U400 ( .A(KEYINPUT3), .B(G119), .ZN(n366) );
  NOR2_X1 U401 ( .A1(n730), .A2(n361), .ZN(n376) );
  XOR2_X1 U402 ( .A(G137), .B(G140), .Z(n434) );
  XNOR2_X1 U403 ( .A(n367), .B(n437), .ZN(n441) );
  XNOR2_X1 U404 ( .A(n436), .B(G110), .ZN(n367) );
  XNOR2_X1 U405 ( .A(G101), .B(G107), .ZN(n436) );
  NAND2_X1 U406 ( .A1(n647), .A2(n390), .ZN(n386) );
  OR2_X1 U407 ( .A1(n610), .A2(n607), .ZN(n369) );
  XNOR2_X1 U408 ( .A(n514), .B(n513), .ZN(n364) );
  INV_X1 U409 ( .A(G101), .ZN(n423) );
  XNOR2_X1 U410 ( .A(G128), .B(G119), .ZN(n396) );
  XOR2_X1 U411 ( .A(G140), .B(G113), .Z(n392) );
  INV_X1 U412 ( .A(KEYINPUT83), .ZN(n527) );
  NAND2_X1 U413 ( .A1(n581), .A2(n580), .ZN(n598) );
  XNOR2_X1 U414 ( .A(n475), .B(G475), .ZN(n476) );
  INV_X1 U415 ( .A(KEYINPUT13), .ZN(n475) );
  INV_X1 U416 ( .A(G902), .ZN(n454) );
  XNOR2_X1 U417 ( .A(G116), .B(G107), .ZN(n481) );
  XNOR2_X1 U418 ( .A(n442), .B(n358), .ZN(n365) );
  NAND2_X1 U419 ( .A1(n375), .A2(n374), .ZN(n373) );
  NAND2_X1 U420 ( .A1(n377), .A2(n376), .ZN(n374) );
  NAND2_X1 U421 ( .A1(n378), .A2(n362), .ZN(n375) );
  XNOR2_X1 U422 ( .A(n650), .B(n552), .ZN(n574) );
  INV_X1 U423 ( .A(KEYINPUT35), .ZN(n372) );
  XNOR2_X1 U424 ( .A(n368), .B(n360), .ZN(n507) );
  NOR2_X1 U425 ( .A1(n564), .A2(n459), .ZN(n368) );
  XNOR2_X1 U426 ( .A(n381), .B(n434), .ZN(n380) );
  XNOR2_X1 U427 ( .A(n435), .B(n433), .ZN(n381) );
  NOR2_X1 U428 ( .A1(n723), .A2(G952), .ZN(n645) );
  NAND2_X1 U429 ( .A1(n385), .A2(n382), .ZN(n740) );
  NAND2_X1 U430 ( .A1(n384), .A2(n383), .ZN(n382) );
  AND2_X1 U431 ( .A1(n387), .A2(n386), .ZN(n385) );
  XNOR2_X1 U432 ( .A(n534), .B(n533), .ZN(n592) );
  AND2_X1 U433 ( .A1(n359), .A2(n599), .ZN(n651) );
  XOR2_X1 U434 ( .A(KEYINPUT16), .B(G122), .Z(n358) );
  AND2_X1 U435 ( .A1(n596), .A2(n597), .ZN(n359) );
  XOR2_X1 U436 ( .A(n460), .B(KEYINPUT19), .Z(n360) );
  NAND2_X1 U437 ( .A1(n607), .A2(n606), .ZN(n361) );
  XNOR2_X1 U438 ( .A(n441), .B(n365), .ZN(n722) );
  AND2_X1 U439 ( .A1(n607), .A2(KEYINPUT2), .ZN(n362) );
  NOR2_X1 U440 ( .A1(KEYINPUT44), .A2(KEYINPUT87), .ZN(n363) );
  NAND2_X1 U441 ( .A1(n364), .A2(n579), .ZN(n535) );
  NAND2_X1 U442 ( .A1(n364), .A2(n532), .ZN(n534) );
  AND2_X1 U443 ( .A1(n364), .A2(n518), .ZN(n602) );
  NAND2_X1 U444 ( .A1(n371), .A2(n599), .ZN(n584) );
  XNOR2_X2 U445 ( .A(n508), .B(n370), .ZN(n599) );
  INV_X1 U446 ( .A(KEYINPUT0), .ZN(n370) );
  INV_X1 U447 ( .A(n589), .ZN(n629) );
  XNOR2_X2 U448 ( .A(n588), .B(n372), .ZN(n589) );
  XNOR2_X2 U449 ( .A(n373), .B(KEYINPUT64), .ZN(n630) );
  OR2_X2 U450 ( .A1(n730), .A2(n716), .ZN(n378) );
  INV_X1 U451 ( .A(n716), .ZN(n377) );
  INV_X1 U452 ( .A(n378), .ZN(n706) );
  XNOR2_X1 U453 ( .A(n441), .B(n380), .ZN(n379) );
  XNOR2_X2 U454 ( .A(n728), .B(G146), .ZN(n438) );
  NAND2_X1 U455 ( .A1(n706), .A2(n606), .ZN(n710) );
  NAND2_X1 U456 ( .A1(n575), .A2(n390), .ZN(n387) );
  INV_X1 U457 ( .A(n740), .ZN(n389) );
  NOR2_X1 U458 ( .A1(n647), .A2(n390), .ZN(n383) );
  INV_X1 U459 ( .A(n575), .ZN(n384) );
  NAND2_X1 U460 ( .A1(n389), .A2(n388), .ZN(n549) );
  INV_X1 U461 ( .A(KEYINPUT40), .ZN(n390) );
  XNOR2_X1 U462 ( .A(n406), .B(n405), .ZN(n631) );
  NAND2_X1 U463 ( .A1(n631), .A2(n454), .ZN(n413) );
  XOR2_X1 U464 ( .A(KEYINPUT94), .B(KEYINPUT12), .Z(n391) );
  INV_X1 U465 ( .A(KEYINPUT67), .ZN(n491) );
  INV_X1 U466 ( .A(KEYINPUT80), .ZN(n433) );
  INV_X1 U467 ( .A(n671), .ZN(n581) );
  INV_X1 U468 ( .A(KEYINPUT105), .ZN(n494) );
  INV_X1 U469 ( .A(KEYINPUT99), .ZN(n552) );
  XNOR2_X1 U470 ( .A(n477), .B(n476), .ZN(n509) );
  OR2_X1 U471 ( .A1(n551), .A2(n550), .ZN(n650) );
  INV_X1 U472 ( .A(n650), .ZN(n662) );
  BUF_X1 U473 ( .A(n631), .Z(n632) );
  XNOR2_X1 U474 ( .A(KEYINPUT15), .B(G902), .ZN(n452) );
  NAND2_X1 U475 ( .A1(G234), .A2(n452), .ZN(n393) );
  XNOR2_X1 U476 ( .A(KEYINPUT20), .B(n393), .ZN(n407) );
  NAND2_X1 U477 ( .A1(n407), .A2(G221), .ZN(n395) );
  XOR2_X1 U478 ( .A(KEYINPUT21), .B(KEYINPUT90), .Z(n394) );
  XNOR2_X1 U479 ( .A(n395), .B(n394), .ZN(n674) );
  XNOR2_X2 U480 ( .A(G146), .B(G125), .ZN(n446) );
  XOR2_X1 U481 ( .A(KEYINPUT24), .B(G110), .Z(n397) );
  XNOR2_X1 U482 ( .A(n397), .B(n396), .ZN(n398) );
  OR2_X2 U483 ( .A1(n729), .A2(n398), .ZN(n400) );
  NAND2_X1 U484 ( .A1(n729), .A2(n398), .ZN(n399) );
  NAND2_X1 U485 ( .A1(n400), .A2(n399), .ZN(n406) );
  NAND2_X1 U486 ( .A1(n723), .A2(G234), .ZN(n402) );
  XNOR2_X1 U487 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n401) );
  XNOR2_X1 U488 ( .A(n402), .B(n401), .ZN(n483) );
  NAND2_X1 U489 ( .A1(n483), .A2(G221), .ZN(n404) );
  XNOR2_X1 U490 ( .A(KEYINPUT71), .B(KEYINPUT23), .ZN(n403) );
  XNOR2_X1 U491 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U492 ( .A(KEYINPUT79), .B(KEYINPUT25), .Z(n409) );
  NAND2_X1 U493 ( .A1(n407), .A2(G217), .ZN(n408) );
  XNOR2_X1 U494 ( .A(n409), .B(n408), .ZN(n411) );
  INV_X1 U495 ( .A(KEYINPUT78), .ZN(n410) );
  XNOR2_X1 U496 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X2 U497 ( .A(n413), .B(n412), .ZN(n490) );
  BUF_X1 U498 ( .A(n490), .Z(n536) );
  NAND2_X1 U499 ( .A1(G234), .A2(G237), .ZN(n414) );
  XOR2_X1 U500 ( .A(n414), .B(KEYINPUT14), .Z(n417) );
  INV_X1 U501 ( .A(n417), .ZN(n415) );
  NAND2_X1 U502 ( .A1(G952), .A2(n415), .ZN(n701) );
  NOR2_X1 U503 ( .A1(n701), .A2(G953), .ZN(n501) );
  NAND2_X1 U504 ( .A1(G953), .A2(G902), .ZN(n416) );
  NOR2_X1 U505 ( .A1(n417), .A2(n416), .ZN(n502) );
  XOR2_X1 U506 ( .A(n502), .B(KEYINPUT104), .Z(n418) );
  NOR2_X1 U507 ( .A1(G900), .A2(n418), .ZN(n419) );
  NOR2_X1 U508 ( .A1(n501), .A2(n419), .ZN(n496) );
  NOR2_X1 U509 ( .A1(n536), .A2(n496), .ZN(n420) );
  NAND2_X1 U510 ( .A1(n674), .A2(n420), .ZN(n520) );
  XOR2_X1 U511 ( .A(KEYINPUT4), .B(G131), .Z(n421) );
  XOR2_X1 U512 ( .A(G137), .B(KEYINPUT5), .Z(n425) );
  NOR2_X1 U513 ( .A1(G953), .A2(G237), .ZN(n463) );
  NAND2_X1 U514 ( .A1(G210), .A2(n463), .ZN(n422) );
  XNOR2_X1 U515 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U516 ( .A(n425), .B(n424), .ZN(n427) );
  XNOR2_X1 U517 ( .A(n427), .B(n442), .ZN(n428) );
  XNOR2_X1 U518 ( .A(n438), .B(n428), .ZN(n623) );
  NAND2_X1 U519 ( .A1(n623), .A2(n454), .ZN(n431) );
  INV_X1 U520 ( .A(KEYINPUT72), .ZN(n429) );
  XNOR2_X1 U521 ( .A(n429), .B(G472), .ZN(n430) );
  XNOR2_X2 U522 ( .A(n431), .B(n430), .ZN(n597) );
  OR2_X1 U523 ( .A1(n520), .A2(n597), .ZN(n432) );
  XNOR2_X1 U524 ( .A(n432), .B(KEYINPUT28), .ZN(n440) );
  NAND2_X1 U525 ( .A1(G227), .A2(n723), .ZN(n435) );
  XNOR2_X1 U526 ( .A(G104), .B(KEYINPUT77), .ZN(n437) );
  XOR2_X1 U527 ( .A(KEYINPUT70), .B(G469), .Z(n439) );
  NOR2_X1 U528 ( .A1(n440), .A2(n516), .ZN(n545) );
  NAND2_X1 U529 ( .A1(n723), .A2(G224), .ZN(n444) );
  XNOR2_X1 U530 ( .A(n444), .B(KEYINPUT4), .ZN(n445) );
  XNOR2_X1 U531 ( .A(n443), .B(n445), .ZN(n450) );
  BUF_X1 U532 ( .A(n446), .Z(n447) );
  XNOR2_X1 U533 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n448) );
  XNOR2_X1 U534 ( .A(n447), .B(n448), .ZN(n449) );
  XNOR2_X1 U535 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U536 ( .A(n722), .B(n451), .ZN(n610) );
  INV_X1 U537 ( .A(n452), .ZN(n607) );
  INV_X1 U538 ( .A(G237), .ZN(n453) );
  NAND2_X1 U539 ( .A1(n454), .A2(n453), .ZN(n458) );
  NAND2_X1 U540 ( .A1(n458), .A2(G210), .ZN(n456) );
  XNOR2_X1 U541 ( .A(KEYINPUT84), .B(KEYINPUT88), .ZN(n455) );
  XNOR2_X1 U542 ( .A(n456), .B(n455), .ZN(n457) );
  NAND2_X1 U543 ( .A1(n458), .A2(G214), .ZN(n689) );
  INV_X1 U544 ( .A(n689), .ZN(n459) );
  INV_X1 U545 ( .A(KEYINPUT65), .ZN(n460) );
  NAND2_X1 U546 ( .A1(n545), .A2(n507), .ZN(n655) );
  XOR2_X1 U547 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n462) );
  XNOR2_X1 U548 ( .A(KEYINPUT95), .B(KEYINPUT11), .ZN(n461) );
  XNOR2_X1 U549 ( .A(n462), .B(n461), .ZN(n465) );
  NAND2_X1 U550 ( .A1(G214), .A2(n463), .ZN(n464) );
  XNOR2_X1 U551 ( .A(n465), .B(n464), .ZN(n468) );
  BUF_X1 U552 ( .A(n466), .Z(n467) );
  XNOR2_X1 U553 ( .A(n468), .B(n467), .ZN(n474) );
  XNOR2_X1 U554 ( .A(G143), .B(G131), .ZN(n469) );
  XNOR2_X1 U555 ( .A(n392), .B(n469), .ZN(n472) );
  XNOR2_X1 U556 ( .A(G104), .B(G122), .ZN(n470) );
  XNOR2_X1 U557 ( .A(n391), .B(n470), .ZN(n471) );
  XNOR2_X1 U558 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U559 ( .A(n474), .B(n473), .ZN(n616) );
  NOR2_X1 U560 ( .A1(n616), .A2(G902), .ZN(n477) );
  XOR2_X1 U561 ( .A(n509), .B(KEYINPUT96), .Z(n551) );
  XOR2_X1 U562 ( .A(KEYINPUT98), .B(KEYINPUT7), .Z(n479) );
  XNOR2_X1 U563 ( .A(G122), .B(KEYINPUT9), .ZN(n478) );
  XNOR2_X1 U564 ( .A(n479), .B(n478), .ZN(n480) );
  XOR2_X1 U565 ( .A(n480), .B(KEYINPUT97), .Z(n482) );
  XNOR2_X1 U566 ( .A(n482), .B(n481), .ZN(n487) );
  NAND2_X1 U567 ( .A1(n483), .A2(G217), .ZN(n484) );
  XNOR2_X1 U568 ( .A(n485), .B(n484), .ZN(n486) );
  XOR2_X1 U569 ( .A(n487), .B(n486), .Z(n635) );
  NOR2_X1 U570 ( .A1(n635), .A2(G902), .ZN(n488) );
  XNOR2_X1 U571 ( .A(n488), .B(G478), .ZN(n550) );
  NAND2_X1 U572 ( .A1(n551), .A2(n550), .ZN(n647) );
  NOR2_X1 U573 ( .A1(n655), .A2(n647), .ZN(n489) );
  XOR2_X1 U574 ( .A(G146), .B(n489), .Z(G48) );
  NAND2_X1 U575 ( .A1(n490), .A2(n674), .ZN(n492) );
  XNOR2_X2 U576 ( .A(n492), .B(n491), .ZN(n671) );
  NOR2_X1 U577 ( .A1(n671), .A2(n516), .ZN(n493) );
  XNOR2_X1 U578 ( .A(n493), .B(KEYINPUT91), .ZN(n595) );
  XNOR2_X1 U579 ( .A(n595), .B(n494), .ZN(n495) );
  NOR2_X1 U580 ( .A1(n496), .A2(n495), .ZN(n541) );
  INV_X1 U581 ( .A(n597), .ZN(n680) );
  NAND2_X1 U582 ( .A1(n689), .A2(n680), .ZN(n497) );
  XOR2_X1 U583 ( .A(KEYINPUT30), .B(n497), .Z(n539) );
  AND2_X1 U584 ( .A1(n541), .A2(n539), .ZN(n500) );
  NOR2_X1 U585 ( .A1(n550), .A2(n509), .ZN(n498) );
  XNOR2_X1 U586 ( .A(n498), .B(KEYINPUT103), .ZN(n585) );
  NOR2_X1 U587 ( .A1(n585), .A2(n564), .ZN(n499) );
  NAND2_X1 U588 ( .A1(n500), .A2(n499), .ZN(n561) );
  XNOR2_X1 U589 ( .A(n561), .B(G143), .ZN(G45) );
  INV_X1 U590 ( .A(n501), .ZN(n505) );
  INV_X1 U591 ( .A(G898), .ZN(n719) );
  AND2_X1 U592 ( .A1(n719), .A2(n502), .ZN(n503) );
  XNOR2_X1 U593 ( .A(n503), .B(KEYINPUT89), .ZN(n504) );
  NAND2_X1 U594 ( .A1(n505), .A2(n504), .ZN(n506) );
  NAND2_X1 U595 ( .A1(n507), .A2(n506), .ZN(n508) );
  NAND2_X1 U596 ( .A1(n509), .A2(n550), .ZN(n692) );
  INV_X1 U597 ( .A(n674), .ZN(n510) );
  NOR2_X1 U598 ( .A1(n692), .A2(n510), .ZN(n511) );
  NAND2_X1 U599 ( .A1(n599), .A2(n511), .ZN(n514) );
  XNOR2_X1 U600 ( .A(KEYINPUT74), .B(KEYINPUT22), .ZN(n512) );
  XNOR2_X1 U601 ( .A(n512), .B(KEYINPUT73), .ZN(n513) );
  INV_X1 U602 ( .A(KEYINPUT6), .ZN(n515) );
  XNOR2_X1 U603 ( .A(n597), .B(n515), .ZN(n582) );
  XNOR2_X1 U604 ( .A(n536), .B(KEYINPUT100), .ZN(n673) );
  NAND2_X1 U605 ( .A1(n579), .A2(n673), .ZN(n517) );
  NOR2_X1 U606 ( .A1(n343), .A2(n517), .ZN(n518) );
  XNOR2_X1 U607 ( .A(G101), .B(KEYINPUT109), .ZN(n519) );
  XNOR2_X1 U608 ( .A(n602), .B(n519), .ZN(G3) );
  NOR2_X1 U609 ( .A1(n647), .A2(n520), .ZN(n521) );
  NAND2_X1 U610 ( .A1(n521), .A2(n689), .ZN(n522) );
  OR2_X1 U611 ( .A1(n522), .A2(n582), .ZN(n565) );
  INV_X1 U612 ( .A(n579), .ZN(n568) );
  NOR2_X1 U613 ( .A1(n565), .A2(n568), .ZN(n524) );
  INV_X1 U614 ( .A(KEYINPUT43), .ZN(n523) );
  XNOR2_X1 U615 ( .A(n524), .B(n523), .ZN(n525) );
  NAND2_X1 U616 ( .A1(n525), .A2(n564), .ZN(n576) );
  XOR2_X1 U617 ( .A(G140), .B(KEYINPUT115), .Z(n526) );
  XNOR2_X1 U618 ( .A(n576), .B(n526), .ZN(G42) );
  XNOR2_X1 U619 ( .A(n582), .B(n527), .ZN(n529) );
  INV_X1 U620 ( .A(n673), .ZN(n528) );
  NAND2_X1 U621 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U622 ( .A1(n530), .A2(n579), .ZN(n531) );
  XNOR2_X1 U623 ( .A(n531), .B(KEYINPUT82), .ZN(n532) );
  XOR2_X1 U624 ( .A(KEYINPUT81), .B(KEYINPUT32), .Z(n533) );
  XNOR2_X1 U625 ( .A(n592), .B(G119), .ZN(G21) );
  XNOR2_X1 U626 ( .A(n535), .B(KEYINPUT101), .ZN(n538) );
  NOR2_X1 U627 ( .A1(n680), .A2(n536), .ZN(n537) );
  NAND2_X1 U628 ( .A1(n538), .A2(n537), .ZN(n593) );
  XNOR2_X1 U629 ( .A(n593), .B(G110), .ZN(G12) );
  XNOR2_X1 U630 ( .A(n564), .B(KEYINPUT38), .ZN(n690) );
  AND2_X1 U631 ( .A1(n539), .A2(n690), .ZN(n540) );
  NAND2_X1 U632 ( .A1(n541), .A2(n540), .ZN(n543) );
  XOR2_X1 U633 ( .A(KEYINPUT86), .B(KEYINPUT39), .Z(n542) );
  XOR2_X1 U634 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n548) );
  NAND2_X1 U635 ( .A1(n690), .A2(n689), .ZN(n687) );
  NOR2_X1 U636 ( .A1(n692), .A2(n687), .ZN(n544) );
  XNOR2_X1 U637 ( .A(KEYINPUT41), .B(n544), .ZN(n703) );
  INV_X1 U638 ( .A(n703), .ZN(n546) );
  NAND2_X1 U639 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U640 ( .A(n548), .B(n547), .ZN(n739) );
  XNOR2_X1 U641 ( .A(n549), .B(KEYINPUT46), .ZN(n572) );
  AND2_X1 U642 ( .A1(n647), .A2(n574), .ZN(n688) );
  NOR2_X2 U643 ( .A1(n655), .A2(n688), .ZN(n558) );
  INV_X1 U644 ( .A(n558), .ZN(n555) );
  INV_X1 U645 ( .A(KEYINPUT76), .ZN(n553) );
  NOR2_X1 U646 ( .A1(n553), .A2(KEYINPUT47), .ZN(n554) );
  NAND2_X1 U647 ( .A1(n555), .A2(n554), .ZN(n560) );
  XNOR2_X1 U648 ( .A(KEYINPUT68), .B(KEYINPUT76), .ZN(n556) );
  XNOR2_X1 U649 ( .A(n556), .B(KEYINPUT47), .ZN(n557) );
  NAND2_X1 U650 ( .A1(n558), .A2(n557), .ZN(n559) );
  NAND2_X1 U651 ( .A1(n560), .A2(n559), .ZN(n562) );
  NAND2_X1 U652 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U653 ( .A(n563), .B(KEYINPUT75), .ZN(n570) );
  XNOR2_X1 U654 ( .A(KEYINPUT107), .B(KEYINPUT36), .ZN(n567) );
  NOR2_X1 U655 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U656 ( .A(n567), .B(n566), .Z(n569) );
  NAND2_X1 U657 ( .A1(n569), .A2(n568), .ZN(n668) );
  NAND2_X1 U658 ( .A1(n570), .A2(n668), .ZN(n571) );
  NOR2_X2 U659 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U660 ( .A(n573), .B(KEYINPUT48), .ZN(n578) );
  OR2_X1 U661 ( .A1(n575), .A2(n574), .ZN(n669) );
  AND2_X1 U662 ( .A1(n669), .A2(n576), .ZN(n577) );
  NAND2_X1 U663 ( .A1(n578), .A2(n577), .ZN(n730) );
  INV_X1 U664 ( .A(KEYINPUT34), .ZN(n583) );
  XNOR2_X1 U665 ( .A(n584), .B(n583), .ZN(n587) );
  INV_X1 U666 ( .A(n585), .ZN(n586) );
  NAND2_X1 U667 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U668 ( .A1(n589), .A2(KEYINPUT87), .ZN(n591) );
  INV_X1 U669 ( .A(KEYINPUT44), .ZN(n590) );
  NAND2_X1 U670 ( .A1(n629), .A2(KEYINPUT44), .ZN(n605) );
  INV_X1 U671 ( .A(n595), .ZN(n596) );
  NOR2_X1 U672 ( .A1(n598), .A2(n597), .ZN(n683) );
  NAND2_X1 U673 ( .A1(n683), .A2(n599), .ZN(n600) );
  XNOR2_X1 U674 ( .A(n600), .B(KEYINPUT31), .ZN(n663) );
  NOR2_X1 U675 ( .A1(n651), .A2(n663), .ZN(n601) );
  NOR2_X1 U676 ( .A1(n601), .A2(n688), .ZN(n603) );
  NOR2_X1 U677 ( .A1(n603), .A2(n602), .ZN(n604) );
  INV_X1 U678 ( .A(KEYINPUT2), .ZN(n606) );
  NAND2_X1 U679 ( .A1(n630), .A2(G210), .ZN(n612) );
  XNOR2_X1 U680 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n608) );
  XOR2_X1 U681 ( .A(n608), .B(KEYINPUT55), .Z(n609) );
  XNOR2_X1 U682 ( .A(n610), .B(n609), .ZN(n611) );
  XNOR2_X1 U683 ( .A(n612), .B(n611), .ZN(n613) );
  NOR2_X2 U684 ( .A1(n613), .A2(n645), .ZN(n614) );
  XNOR2_X1 U685 ( .A(n614), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U686 ( .A1(n630), .A2(G475), .ZN(n618) );
  XOR2_X1 U687 ( .A(KEYINPUT122), .B(KEYINPUT59), .Z(n615) );
  XNOR2_X1 U688 ( .A(n616), .B(n615), .ZN(n617) );
  XNOR2_X1 U689 ( .A(n618), .B(n617), .ZN(n619) );
  NOR2_X2 U690 ( .A1(n619), .A2(n645), .ZN(n622) );
  XNOR2_X1 U691 ( .A(KEYINPUT123), .B(KEYINPUT60), .ZN(n620) );
  XOR2_X1 U692 ( .A(n620), .B(KEYINPUT66), .Z(n621) );
  XNOR2_X1 U693 ( .A(n622), .B(n621), .ZN(G60) );
  NAND2_X1 U694 ( .A1(n630), .A2(G472), .ZN(n625) );
  XOR2_X1 U695 ( .A(KEYINPUT62), .B(n623), .Z(n624) );
  XNOR2_X1 U696 ( .A(n625), .B(n624), .ZN(n626) );
  NOR2_X2 U697 ( .A1(n626), .A2(n645), .ZN(n628) );
  XOR2_X1 U698 ( .A(KEYINPUT108), .B(KEYINPUT63), .Z(n627) );
  XNOR2_X1 U699 ( .A(n628), .B(n627), .ZN(G57) );
  XOR2_X1 U700 ( .A(n629), .B(G122), .Z(G24) );
  BUF_X2 U701 ( .A(n630), .Z(n639) );
  NAND2_X1 U702 ( .A1(n639), .A2(G217), .ZN(n633) );
  XOR2_X1 U703 ( .A(n633), .B(n632), .Z(n634) );
  NOR2_X1 U704 ( .A1(n634), .A2(n645), .ZN(G66) );
  NAND2_X1 U705 ( .A1(n639), .A2(G478), .ZN(n637) );
  XNOR2_X1 U706 ( .A(n635), .B(KEYINPUT124), .ZN(n636) );
  XNOR2_X1 U707 ( .A(n637), .B(n636), .ZN(n638) );
  NOR2_X1 U708 ( .A1(n638), .A2(n645), .ZN(G63) );
  NAND2_X1 U709 ( .A1(n639), .A2(G469), .ZN(n644) );
  XOR2_X1 U710 ( .A(KEYINPUT121), .B(KEYINPUT57), .Z(n640) );
  XNOR2_X1 U711 ( .A(n640), .B(KEYINPUT58), .ZN(n641) );
  XNOR2_X1 U712 ( .A(n357), .B(n641), .ZN(n643) );
  XNOR2_X1 U713 ( .A(n644), .B(n643), .ZN(n646) );
  NOR2_X1 U714 ( .A1(n646), .A2(n645), .ZN(G54) );
  INV_X1 U715 ( .A(n647), .ZN(n659) );
  NAND2_X1 U716 ( .A1(n651), .A2(n659), .ZN(n648) );
  XNOR2_X1 U717 ( .A(n648), .B(KEYINPUT110), .ZN(n649) );
  XNOR2_X1 U718 ( .A(G104), .B(n649), .ZN(G6) );
  XOR2_X1 U719 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n653) );
  NAND2_X1 U720 ( .A1(n651), .A2(n662), .ZN(n652) );
  XNOR2_X1 U721 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U722 ( .A(G107), .B(n654), .ZN(G9) );
  NOR2_X1 U723 ( .A1(n655), .A2(n650), .ZN(n657) );
  XNOR2_X1 U724 ( .A(KEYINPUT29), .B(KEYINPUT111), .ZN(n656) );
  XNOR2_X1 U725 ( .A(n657), .B(n656), .ZN(n658) );
  XOR2_X1 U726 ( .A(G128), .B(n658), .Z(G30) );
  NAND2_X1 U727 ( .A1(n663), .A2(n659), .ZN(n660) );
  XNOR2_X1 U728 ( .A(n660), .B(KEYINPUT112), .ZN(n661) );
  XNOR2_X1 U729 ( .A(G113), .B(n661), .ZN(G15) );
  XOR2_X1 U730 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n665) );
  NAND2_X1 U731 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U732 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U733 ( .A(G116), .B(n666), .ZN(G18) );
  XOR2_X1 U734 ( .A(G125), .B(KEYINPUT37), .Z(n667) );
  XNOR2_X1 U735 ( .A(n668), .B(n667), .ZN(G27) );
  INV_X1 U736 ( .A(n669), .ZN(n670) );
  XOR2_X1 U737 ( .A(G134), .B(n670), .Z(G36) );
  NAND2_X1 U738 ( .A1(n579), .A2(n671), .ZN(n672) );
  XNOR2_X1 U739 ( .A(KEYINPUT50), .B(n672), .ZN(n678) );
  NOR2_X1 U740 ( .A1(n674), .A2(n673), .ZN(n676) );
  XNOR2_X1 U741 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n675) );
  XNOR2_X1 U742 ( .A(n676), .B(n675), .ZN(n677) );
  NAND2_X1 U743 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U744 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U745 ( .A(KEYINPUT117), .B(n681), .Z(n682) );
  NOR2_X1 U746 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U747 ( .A(KEYINPUT51), .B(n684), .Z(n685) );
  NOR2_X1 U748 ( .A1(n703), .A2(n685), .ZN(n697) );
  NOR2_X1 U749 ( .A1(n688), .A2(n687), .ZN(n694) );
  NOR2_X1 U750 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U751 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U752 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U753 ( .A1(n686), .A2(n695), .ZN(n696) );
  NOR2_X1 U754 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U755 ( .A(n698), .B(KEYINPUT52), .ZN(n699) );
  XNOR2_X1 U756 ( .A(KEYINPUT118), .B(n699), .ZN(n700) );
  NOR2_X1 U757 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U758 ( .A(n702), .B(KEYINPUT119), .ZN(n705) );
  OR2_X1 U759 ( .A1(n686), .A2(n703), .ZN(n704) );
  NAND2_X1 U760 ( .A1(n705), .A2(n704), .ZN(n713) );
  OR2_X1 U761 ( .A1(n706), .A2(KEYINPUT85), .ZN(n707) );
  NAND2_X1 U762 ( .A1(n707), .A2(KEYINPUT2), .ZN(n709) );
  OR2_X1 U763 ( .A1(KEYINPUT2), .A2(KEYINPUT85), .ZN(n708) );
  NAND2_X1 U764 ( .A1(n709), .A2(n708), .ZN(n711) );
  NAND2_X1 U765 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U766 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U767 ( .A1(n723), .A2(n714), .ZN(n715) );
  XOR2_X1 U768 ( .A(KEYINPUT53), .B(n715), .Z(G75) );
  NOR2_X1 U769 ( .A1(n356), .A2(G953), .ZN(n721) );
  NAND2_X1 U770 ( .A1(G953), .A2(G224), .ZN(n717) );
  XOR2_X1 U771 ( .A(KEYINPUT61), .B(n717), .Z(n718) );
  NOR2_X1 U772 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U773 ( .A1(n721), .A2(n720), .ZN(n727) );
  XOR2_X1 U774 ( .A(KEYINPUT125), .B(n722), .Z(n725) );
  NOR2_X1 U775 ( .A1(n723), .A2(G898), .ZN(n724) );
  NOR2_X1 U776 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U777 ( .A(n727), .B(n726), .Z(G69) );
  XOR2_X1 U778 ( .A(n728), .B(n729), .Z(n732) );
  XOR2_X1 U779 ( .A(n730), .B(n732), .Z(n731) );
  NOR2_X1 U780 ( .A1(n731), .A2(G953), .ZN(n737) );
  XNOR2_X1 U781 ( .A(G227), .B(n732), .ZN(n733) );
  NAND2_X1 U782 ( .A1(n733), .A2(G900), .ZN(n734) );
  NAND2_X1 U783 ( .A1(n734), .A2(G953), .ZN(n735) );
  XOR2_X1 U784 ( .A(KEYINPUT126), .B(n735), .Z(n736) );
  NOR2_X1 U785 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U786 ( .A(KEYINPUT127), .B(n738), .ZN(G72) );
  XOR2_X1 U787 ( .A(G137), .B(n739), .Z(G39) );
  XOR2_X1 U788 ( .A(n740), .B(G131), .Z(G33) );
endmodule

