//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0 0 1 0 1 0 1 0 0 1 0 1 1 0 0 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 0 1 0 1 0 1 1 1 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n570, new_n572, new_n573, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n633, new_n636, new_n638, new_n639, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1201, new_n1202;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT67), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n465));
  XNOR2_X1  g040(.A(new_n464), .B(new_n465), .ZN(new_n466));
  AND3_X1   g041(.A1(KEYINPUT66), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(KEYINPUT3), .B1(KEYINPUT66), .B2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G137), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT3), .B(G2104), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n472), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n471), .B1(new_n461), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n466), .A2(new_n474), .ZN(G160));
  OAI21_X1  g050(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(G112), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(G2105), .ZN(new_n478));
  OAI21_X1  g053(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT69), .ZN(new_n482));
  AOI211_X1 g057(.A(new_n478), .B(new_n482), .C1(G136), .C2(new_n470), .ZN(G162));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n484));
  AND4_X1   g059(.A1(new_n484), .A2(new_n472), .A3(G138), .A4(new_n461), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n470), .A2(G138), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(KEYINPUT4), .ZN(new_n487));
  XNOR2_X1  g062(.A(KEYINPUT70), .B(G114), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G126), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(new_n479), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n487), .A2(new_n492), .ZN(G164));
  INV_X1    g068(.A(KEYINPUT72), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT5), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n494), .B1(new_n495), .B2(G543), .ZN(new_n496));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n497), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT71), .A2(G651), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT6), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(KEYINPUT71), .A2(KEYINPUT6), .A3(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n495), .A2(G543), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n499), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT73), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n497), .A2(KEYINPUT5), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n509), .B1(new_n496), .B2(new_n498), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n510), .A2(KEYINPUT73), .A3(new_n504), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n508), .A2(G88), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n504), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G50), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT74), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT74), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n512), .A2(new_n518), .A3(new_n515), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  OAI21_X1  g096(.A(KEYINPUT75), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  AND3_X1   g098(.A1(new_n497), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n524));
  AOI21_X1  g099(.A(KEYINPUT72), .B1(new_n497), .B2(KEYINPUT5), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n505), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G62), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n523), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT75), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n528), .A2(new_n529), .A3(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n522), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n517), .A2(new_n519), .A3(new_n531), .ZN(G303));
  INV_X1    g107(.A(G303), .ZN(G166));
  AND4_X1   g108(.A1(KEYINPUT73), .A2(new_n499), .A3(new_n504), .A4(new_n505), .ZN(new_n534));
  AOI21_X1  g109(.A(KEYINPUT73), .B1(new_n510), .B2(new_n504), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G89), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT7), .ZN(new_n538));
  NAND2_X1  g113(.A1(G76), .A2(G543), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n539), .B2(new_n521), .ZN(new_n540));
  XNOR2_X1  g115(.A(KEYINPUT76), .B(G51), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n513), .B2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(G63), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n526), .A2(new_n543), .B1(new_n538), .B2(new_n539), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n542), .B1(G651), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n537), .A2(new_n545), .ZN(G286));
  INV_X1    g121(.A(G286), .ZN(G168));
  NAND2_X1  g122(.A1(G77), .A2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G64), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n526), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G651), .ZN(new_n551));
  INV_X1    g126(.A(G52), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n508), .A2(new_n511), .ZN(new_n553));
  INV_X1    g128(.A(G90), .ZN(new_n554));
  OAI221_X1 g129(.A(new_n551), .B1(new_n552), .B2(new_n513), .C1(new_n553), .C2(new_n554), .ZN(G301));
  INV_X1    g130(.A(G301), .ZN(G171));
  NAND3_X1  g131(.A1(new_n508), .A2(G81), .A3(new_n511), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT77), .ZN(new_n558));
  NAND2_X1  g133(.A1(G68), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n560), .B1(new_n510), .B2(G56), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n558), .B1(new_n561), .B2(new_n521), .ZN(new_n562));
  OAI211_X1 g137(.A(G56), .B(new_n505), .C1(new_n524), .C2(new_n525), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(new_n559), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n564), .A2(KEYINPUT77), .A3(G651), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n514), .A2(G43), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n557), .A2(new_n562), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G860), .ZN(G153));
  AND3_X1   g144(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G36), .ZN(G176));
  NAND2_X1  g146(.A1(G1), .A2(G3), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT8), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n570), .A2(new_n573), .ZN(G188));
  OAI211_X1 g149(.A(G65), .B(new_n505), .C1(new_n524), .C2(new_n525), .ZN(new_n575));
  NAND2_X1  g150(.A1(G78), .A2(G543), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n503), .ZN(new_n578));
  AOI21_X1  g153(.A(KEYINPUT6), .B1(KEYINPUT71), .B2(G651), .ZN(new_n579));
  OAI211_X1 g154(.A(G53), .B(G543), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(KEYINPUT9), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT9), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n504), .A2(new_n582), .A3(G53), .A4(G543), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n577), .A2(G651), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n508), .A2(G91), .A3(new_n511), .ZN(new_n585));
  AND2_X1   g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G299));
  OAI21_X1  g162(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n588), .B(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n536), .A2(G87), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n514), .A2(G49), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(G288));
  AOI22_X1  g168(.A1(new_n536), .A2(G86), .B1(G48), .B2(new_n514), .ZN(new_n594));
  OAI211_X1 g169(.A(G61), .B(new_n505), .C1(new_n524), .C2(new_n525), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n595), .A2(KEYINPUT79), .B1(G73), .B2(G543), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT79), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n510), .A2(new_n597), .A3(G61), .ZN(new_n598));
  AOI211_X1 g173(.A(KEYINPUT80), .B(new_n521), .C1(new_n596), .C2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT80), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n595), .A2(KEYINPUT79), .ZN(new_n601));
  NAND2_X1  g176(.A1(G73), .A2(G543), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n601), .A2(new_n598), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n600), .B1(new_n603), .B2(G651), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n594), .B1(new_n599), .B2(new_n604), .ZN(G305));
  NAND2_X1  g180(.A1(new_n536), .A2(G85), .ZN(new_n606));
  NAND2_X1  g181(.A1(G72), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G60), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n526), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n609), .A2(G651), .B1(G47), .B2(new_n514), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n606), .A2(new_n610), .ZN(G290));
  NAND2_X1  g186(.A1(G301), .A2(G868), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT81), .ZN(new_n613));
  AND2_X1   g188(.A1(new_n514), .A2(G54), .ZN(new_n614));
  AND2_X1   g189(.A1(KEYINPUT82), .A2(G66), .ZN(new_n615));
  NOR2_X1   g190(.A1(KEYINPUT82), .A2(G66), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n510), .A2(new_n617), .B1(G79), .B2(G543), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT83), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n521), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(G79), .A2(G543), .ZN(new_n621));
  INV_X1    g196(.A(new_n617), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n526), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(KEYINPUT83), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n614), .B1(new_n620), .B2(new_n624), .ZN(new_n625));
  AOI21_X1  g200(.A(KEYINPUT10), .B1(new_n536), .B2(G92), .ZN(new_n626));
  NAND4_X1  g201(.A1(new_n508), .A2(KEYINPUT10), .A3(G92), .A4(new_n511), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n625), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n613), .B1(G868), .B2(new_n630), .ZN(G284));
  OAI21_X1  g206(.A(new_n613), .B1(G868), .B2(new_n630), .ZN(G321));
  NAND2_X1  g207(.A1(G286), .A2(G868), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(G868), .B2(new_n586), .ZN(G297));
  OAI21_X1  g209(.A(new_n633), .B1(G868), .B2(new_n586), .ZN(G280));
  INV_X1    g210(.A(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n630), .B1(new_n636), .B2(G860), .ZN(G148));
  NAND2_X1  g212(.A1(new_n630), .A2(new_n636), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(G868), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(G868), .B2(new_n568), .ZN(G323));
  XNOR2_X1  g215(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g216(.A1(new_n463), .A2(new_n472), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT13), .B(G2100), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n470), .A2(G135), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n480), .A2(G123), .ZN(new_n648));
  OR2_X1    g223(.A1(G99), .A2(G2105), .ZN(new_n649));
  OAI211_X1 g224(.A(new_n649), .B(G2104), .C1(G111), .C2(new_n461), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n647), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n651), .A2(G2096), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(G2096), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n646), .A2(new_n652), .A3(new_n653), .ZN(G156));
  INV_X1    g229(.A(KEYINPUT14), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2427), .B(G2438), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2430), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT15), .B(G2435), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n659), .B1(new_n658), .B2(new_n657), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2451), .B(G2454), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT16), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1341), .B(G1348), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n660), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2443), .B(G2446), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  AND3_X1   g243(.A1(new_n667), .A2(G14), .A3(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT85), .Z(G401));
  XOR2_X1   g245(.A(G2084), .B(G2090), .Z(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2072), .B(G2078), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n672), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT87), .ZN(new_n676));
  INV_X1    g251(.A(new_n673), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n674), .B(KEYINPUT17), .Z(new_n678));
  OAI21_X1  g253(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n678), .A2(new_n677), .A3(new_n671), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n671), .A2(new_n673), .A3(new_n674), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT86), .B(KEYINPUT18), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n679), .A2(new_n680), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G2096), .B(G2100), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(G227));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT19), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G1956), .B(G2474), .Z(new_n690));
  XOR2_X1   g265(.A(G1961), .B(G1966), .Z(new_n691));
  AND2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT20), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n690), .A2(new_n691), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  MUX2_X1   g272(.A(new_n697), .B(new_n696), .S(new_n689), .Z(new_n698));
  NOR2_X1   g273(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1991), .B(G1996), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1981), .B(G1986), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(G229));
  INV_X1    g280(.A(G29), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G35), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G162), .B2(new_n706), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT29), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n709), .A2(G2090), .ZN(new_n710));
  INV_X1    g285(.A(G16), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G20), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT23), .Z(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(G299), .B2(G16), .ZN(new_n714));
  INV_X1    g289(.A(G1956), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n568), .A2(new_n711), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n711), .B2(G19), .ZN(new_n718));
  INV_X1    g293(.A(G1341), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR3_X1   g295(.A1(new_n710), .A2(new_n716), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(G160), .A2(G29), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT95), .B(KEYINPUT24), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(G34), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n722), .B1(G29), .B2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(G2084), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n711), .A2(G5), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G171), .B2(new_n711), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n706), .A2(G32), .ZN(new_n730));
  NAND3_X1  g305(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT26), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n731), .A2(new_n732), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n463), .A2(G105), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n470), .A2(G141), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n480), .A2(G129), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT96), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n738), .A2(new_n739), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n730), .B1(new_n742), .B2(G29), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT27), .B(G1996), .ZN(new_n744));
  OAI221_X1 g319(.A(new_n727), .B1(G1961), .B2(new_n729), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n721), .B1(KEYINPUT99), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(G27), .A2(G29), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G164), .B2(G29), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT100), .B(G2078), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT31), .B(G11), .Z(new_n751));
  NOR2_X1   g326(.A1(new_n651), .A2(new_n706), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT98), .B(G28), .Z(new_n753));
  OR2_X1    g328(.A1(new_n753), .A2(KEYINPUT30), .ZN(new_n754));
  AOI21_X1  g329(.A(G29), .B1(new_n753), .B2(KEYINPUT30), .ZN(new_n755));
  AOI211_X1 g330(.A(new_n751), .B(new_n752), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n750), .B(new_n756), .C1(new_n725), .C2(new_n726), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n748), .A2(new_n749), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n706), .A2(G33), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n472), .A2(G127), .ZN(new_n760));
  NAND2_X1  g335(.A1(G115), .A2(G2104), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT94), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n461), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n763), .B2(new_n762), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT93), .B(KEYINPUT25), .ZN(new_n766));
  AND3_X1   g341(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n766), .A2(new_n767), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n768), .A2(new_n769), .B1(new_n470), .B2(G139), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n765), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n759), .B1(new_n771), .B2(new_n706), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n758), .B1(G2072), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G2072), .B2(new_n772), .ZN(new_n774));
  AOI211_X1 g349(.A(new_n757), .B(new_n774), .C1(new_n743), .C2(new_n744), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n709), .A2(G2090), .B1(new_n719), .B2(new_n718), .ZN(new_n776));
  NAND2_X1  g351(.A1(G168), .A2(G16), .ZN(new_n777));
  NOR2_X1   g352(.A1(G16), .A2(G21), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n777), .B1(KEYINPUT97), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(KEYINPUT97), .B2(new_n777), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1966), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n706), .A2(G26), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT28), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n470), .A2(G140), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n480), .A2(G128), .ZN(new_n785));
  OR2_X1    g360(.A1(G104), .A2(G2105), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n786), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n784), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n783), .B1(new_n788), .B2(G29), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT92), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G2067), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G1961), .B2(new_n729), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n775), .A2(new_n776), .A3(new_n781), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n745), .A2(KEYINPUT99), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n711), .A2(G4), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n630), .B2(new_n711), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT91), .B(G1348), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n794), .A2(new_n798), .ZN(new_n799));
  NOR3_X1   g374(.A1(new_n746), .A2(new_n793), .A3(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT36), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n706), .A2(G25), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n470), .A2(G131), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n480), .A2(G119), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n461), .A2(G107), .ZN(new_n806));
  OAI21_X1  g381(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n804), .B(new_n805), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT88), .Z(new_n809));
  OAI21_X1  g384(.A(new_n803), .B1(new_n809), .B2(new_n706), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT35), .B(G1991), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n711), .A2(G24), .ZN(new_n813));
  INV_X1    g388(.A(G290), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n813), .B1(new_n814), .B2(new_n711), .ZN(new_n815));
  INV_X1    g390(.A(G1986), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n812), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n711), .A2(G23), .ZN(new_n819));
  AND3_X1   g394(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(new_n820), .B2(new_n711), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT33), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G1976), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n711), .A2(G6), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n514), .A2(G48), .ZN(new_n825));
  INV_X1    g400(.A(G86), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n553), .B2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n604), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n521), .B1(new_n596), .B2(new_n598), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(new_n600), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n827), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n824), .B1(new_n831), .B2(new_n711), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT32), .B(G1981), .Z(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(G16), .A2(G22), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(G166), .B2(G16), .ZN(new_n836));
  INV_X1    g411(.A(G1971), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n823), .A2(new_n834), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(KEYINPUT90), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT90), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n823), .A2(new_n841), .A3(new_n834), .A4(new_n838), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(KEYINPUT89), .B(KEYINPUT34), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n818), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n844), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n840), .A2(new_n842), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n802), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n845), .A2(new_n802), .A3(new_n847), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n801), .B1(new_n849), .B2(new_n850), .ZN(G311));
  INV_X1    g426(.A(new_n850), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n800), .B1(new_n852), .B2(new_n848), .ZN(G150));
  NAND2_X1  g428(.A1(new_n630), .A2(G559), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT38), .ZN(new_n855));
  AOI22_X1  g430(.A1(new_n536), .A2(G81), .B1(G43), .B2(new_n514), .ZN(new_n856));
  AOI21_X1  g431(.A(KEYINPUT77), .B1(new_n564), .B2(G651), .ZN(new_n857));
  AOI211_X1 g432(.A(new_n558), .B(new_n521), .C1(new_n563), .C2(new_n559), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n508), .A2(G93), .A3(new_n511), .ZN(new_n860));
  NAND2_X1  g435(.A1(G80), .A2(G543), .ZN(new_n861));
  INV_X1    g436(.A(G67), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n861), .B1(new_n526), .B2(new_n862), .ZN(new_n863));
  AOI22_X1  g438(.A1(new_n863), .A2(G651), .B1(G55), .B2(new_n514), .ZN(new_n864));
  AOI22_X1  g439(.A1(new_n856), .A2(new_n859), .B1(new_n860), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n860), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n567), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n855), .B(new_n868), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n869), .A2(KEYINPUT39), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(KEYINPUT39), .ZN(new_n871));
  NOR3_X1   g446(.A1(new_n870), .A2(new_n871), .A3(G860), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n866), .A2(G860), .ZN(new_n873));
  XOR2_X1   g448(.A(KEYINPUT101), .B(KEYINPUT37), .Z(new_n874));
  XOR2_X1   g449(.A(new_n873), .B(new_n874), .Z(new_n875));
  OR2_X1    g450(.A1(new_n872), .A2(new_n875), .ZN(G145));
  NAND2_X1  g451(.A1(new_n470), .A2(G142), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n480), .A2(G130), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n461), .A2(G118), .ZN(new_n879));
  OAI21_X1  g454(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n877), .B(new_n878), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n808), .B(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(G164), .B(KEYINPUT102), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n771), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n883), .A2(new_n771), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n882), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n886), .ZN(new_n888));
  INV_X1    g463(.A(new_n882), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n888), .A2(new_n884), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n742), .A2(new_n788), .ZN(new_n892));
  INV_X1    g467(.A(new_n788), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n893), .B1(new_n740), .B2(new_n741), .ZN(new_n894));
  OR3_X1    g469(.A1(new_n892), .A2(new_n644), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n644), .B1(new_n892), .B2(new_n894), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n891), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(G160), .B(new_n651), .ZN(new_n899));
  XOR2_X1   g474(.A(new_n899), .B(G162), .Z(new_n900));
  NAND4_X1  g475(.A1(new_n887), .A2(new_n890), .A3(new_n895), .A4(new_n896), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n898), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(G37), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n900), .B1(new_n898), .B2(new_n901), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n905), .A2(KEYINPUT103), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT103), .ZN(new_n907));
  AOI211_X1 g482(.A(new_n907), .B(new_n900), .C1(new_n898), .C2(new_n901), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n904), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g485(.A1(new_n831), .A2(G303), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n519), .A2(new_n531), .ZN(new_n912));
  NAND3_X1  g487(.A1(G305), .A2(new_n912), .A3(new_n517), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n606), .A2(KEYINPUT105), .A3(new_n610), .ZN(new_n915));
  AOI21_X1  g490(.A(KEYINPUT105), .B1(new_n606), .B2(new_n610), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n820), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT105), .ZN(new_n918));
  NAND2_X1  g493(.A1(G290), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n606), .A2(KEYINPUT105), .A3(new_n610), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n919), .A2(G288), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n917), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n914), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n911), .A2(new_n913), .A3(new_n917), .A4(new_n921), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n925), .A2(KEYINPUT106), .ZN(new_n926));
  XOR2_X1   g501(.A(new_n926), .B(KEYINPUT42), .Z(new_n927));
  XOR2_X1   g502(.A(new_n638), .B(new_n868), .Z(new_n928));
  XNOR2_X1  g503(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n508), .A2(G92), .A3(new_n511), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT10), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n627), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n934), .A2(new_n586), .A3(new_n625), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n586), .B1(new_n934), .B2(new_n625), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n930), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n629), .A2(G299), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT41), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n934), .A2(new_n586), .A3(new_n625), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n928), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n935), .A2(new_n936), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n943), .B1(new_n945), .B2(new_n928), .ZN(new_n946));
  XOR2_X1   g521(.A(new_n927), .B(new_n946), .Z(new_n947));
  MUX2_X1   g522(.A(new_n866), .B(new_n947), .S(G868), .Z(G295));
  MUX2_X1   g523(.A(new_n866), .B(new_n947), .S(G868), .Z(G331));
  OAI21_X1  g524(.A(G171), .B1(new_n865), .B2(new_n867), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n856), .A2(new_n859), .A3(new_n860), .A4(new_n864), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n567), .A2(new_n866), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(G301), .A3(new_n952), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n950), .A2(G168), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(G168), .B1(new_n950), .B2(new_n953), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n944), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n951), .A2(G301), .A3(new_n952), .ZN(new_n957));
  AOI21_X1  g532(.A(G301), .B1(new_n951), .B2(new_n952), .ZN(new_n958));
  OAI21_X1  g533(.A(G286), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n950), .A2(G168), .A3(new_n953), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n959), .A2(new_n942), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n956), .A2(new_n925), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n903), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n925), .B1(new_n956), .B2(new_n961), .ZN(new_n964));
  OR3_X1    g539(.A1(new_n963), .A2(KEYINPUT43), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n925), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n939), .B1(new_n935), .B2(new_n936), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n938), .A2(new_n940), .A3(new_n930), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n954), .A2(new_n969), .A3(new_n955), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n945), .B1(new_n959), .B2(new_n960), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n966), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT109), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n959), .A2(new_n960), .A3(new_n968), .A4(new_n967), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n956), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n976), .A2(KEYINPUT109), .A3(new_n966), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n963), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT43), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n965), .B(KEYINPUT44), .C1(new_n978), .C2(new_n979), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n962), .A2(new_n903), .ZN(new_n981));
  AOI21_X1  g556(.A(KEYINPUT109), .B1(new_n976), .B2(new_n966), .ZN(new_n982));
  AOI211_X1 g557(.A(new_n973), .B(new_n925), .C1(new_n956), .C2(new_n975), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n981), .B(new_n979), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT110), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n974), .A2(new_n977), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n987), .A2(KEYINPUT110), .A3(new_n979), .A4(new_n981), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT43), .B1(new_n963), .B2(new_n964), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(KEYINPUT108), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT108), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n991), .B(KEYINPUT43), .C1(new_n963), .C2(new_n964), .ZN(new_n992));
  AOI22_X1  g567(.A1(new_n986), .A2(new_n988), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  XOR2_X1   g568(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n994));
  OAI21_X1  g569(.A(new_n980), .B1(new_n993), .B2(new_n994), .ZN(G397));
  INV_X1    g570(.A(G1384), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n996), .B1(new_n487), .B2(new_n492), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT45), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G40), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n466), .A2(new_n1001), .A3(new_n474), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G1996), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  XOR2_X1   g580(.A(new_n1005), .B(KEYINPUT111), .Z(new_n1006));
  NOR2_X1   g581(.A1(new_n1006), .A2(new_n742), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n788), .A2(G2067), .ZN(new_n1008));
  INV_X1    g583(.A(G2067), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n893), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1003), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1003), .A2(new_n742), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1011), .B1(new_n1012), .B2(new_n1004), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1007), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1003), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n808), .B(new_n811), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1014), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n814), .A2(new_n816), .ZN(new_n1018));
  NAND2_X1  g593(.A1(G290), .A2(G1986), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1015), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT63), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1023), .B(new_n996), .C1(new_n487), .C2(new_n492), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n1024), .B(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n997), .A2(KEYINPUT50), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n1002), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G2090), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1026), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  OAI211_X1 g605(.A(KEYINPUT45), .B(new_n996), .C1(new_n487), .C2(new_n492), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1002), .A2(new_n999), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n837), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1030), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1030), .A2(KEYINPUT115), .A3(new_n1033), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1036), .A2(G8), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(G303), .A2(G8), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n1040));
  XNOR2_X1  g615(.A(new_n1039), .B(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1038), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G8), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1002), .A2(new_n1027), .A3(new_n1029), .A4(new_n1024), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1044), .B1(new_n1033), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1041), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT112), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1041), .A2(new_n1046), .A3(KEYINPUT112), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n997), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1044), .B1(new_n1002), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G1976), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1053), .B1(new_n1054), .B2(G288), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT52), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1057), .B1(new_n820), .B2(G1976), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1056), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G1981), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n831), .A2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(G1981), .B1(new_n827), .B2(new_n829), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(KEYINPUT49), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT49), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1053), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1059), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1043), .A2(new_n1051), .A3(new_n1067), .ZN(new_n1068));
  AND3_X1   g643(.A1(new_n1002), .A2(new_n1027), .A3(new_n1024), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(new_n726), .ZN(new_n1070));
  INV_X1    g645(.A(G1966), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1032), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1044), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(G168), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1022), .B1(new_n1068), .B2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1041), .A2(new_n1046), .ZN(new_n1076));
  NOR3_X1   g651(.A1(new_n1074), .A2(new_n1076), .A3(new_n1022), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1077), .A2(new_n1051), .A3(new_n1067), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT116), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1077), .A2(new_n1051), .A3(new_n1080), .A4(new_n1067), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1075), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  OR2_X1    g657(.A1(new_n1069), .A2(G1961), .ZN(new_n1083));
  INV_X1    g658(.A(G2078), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1002), .A2(new_n999), .A3(new_n1084), .A4(new_n1031), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1085), .A2(KEYINPUT124), .A3(KEYINPUT53), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT53), .B1(new_n1085), .B2(KEYINPUT124), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1083), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(G171), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1068), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(G8), .ZN(new_n1092));
  NAND2_X1  g667(.A1(G286), .A2(G8), .ZN(new_n1093));
  XOR2_X1   g668(.A(new_n1093), .B(KEYINPUT122), .Z(new_n1094));
  INV_X1    g669(.A(KEYINPUT123), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT51), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1092), .B(new_n1094), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1094), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(new_n1091), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n1073), .B2(new_n1098), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT51), .B1(new_n1073), .B2(KEYINPUT123), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1097), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT62), .ZN(new_n1103));
  OR2_X1    g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1090), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  AOI211_X1 g681(.A(G1976), .B(G288), .C1(new_n1066), .C2(new_n1063), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1061), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1053), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1067), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  OR2_X1    g686(.A1(new_n1111), .A2(KEYINPUT113), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(KEYINPUT113), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1082), .A2(new_n1106), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1043), .A2(new_n1051), .A3(new_n1067), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1083), .B(G301), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT54), .B1(new_n1089), .B2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1102), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1089), .A2(KEYINPUT54), .A3(new_n1116), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n1119), .A2(KEYINPUT125), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1119), .A2(KEYINPUT125), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1115), .B(new_n1118), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT61), .ZN(new_n1123));
  XNOR2_X1  g698(.A(new_n586), .B(KEYINPUT57), .ZN(new_n1124));
  AOI21_X1  g699(.A(G1956), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT117), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n1125), .B(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1032), .ZN(new_n1128));
  XNOR2_X1  g703(.A(KEYINPUT56), .B(G2072), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1124), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1126), .B1(new_n1132), .B2(new_n715), .ZN(new_n1133));
  AOI211_X1 g708(.A(KEYINPUT117), .B(G1956), .C1(new_n1026), .C2(new_n1028), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1130), .B(new_n1124), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1123), .B1(new_n1131), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT121), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1002), .A2(new_n1027), .A3(new_n1024), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(new_n797), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1002), .A2(new_n1009), .A3(new_n1052), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT60), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1142), .A2(new_n1143), .A3(new_n630), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1140), .A2(new_n629), .A3(new_n1141), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n629), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT60), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT59), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1002), .A2(new_n999), .A3(new_n1004), .A4(new_n1031), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT119), .ZN(new_n1150));
  OR2_X1    g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1002), .A2(new_n1052), .ZN(new_n1152));
  XNOR2_X1  g727(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1153), .B(new_n719), .ZN(new_n1154));
  AOI22_X1  g729(.A1(new_n1149), .A2(new_n1150), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1151), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1148), .B1(new_n1156), .B2(new_n568), .ZN(new_n1157));
  AOI211_X1 g732(.A(KEYINPUT59), .B(new_n567), .C1(new_n1151), .C2(new_n1155), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1144), .B(new_n1147), .C1(new_n1157), .C2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1130), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT118), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  OAI211_X1 g737(.A(KEYINPUT118), .B(new_n1130), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1124), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n1135), .A2(KEYINPUT61), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1159), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT121), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1168), .B(new_n1123), .C1(new_n1131), .C2(new_n1136), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1138), .A2(new_n1167), .A3(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1165), .B1(new_n629), .B2(new_n1142), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(new_n1135), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1122), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1021), .B1(new_n1114), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n809), .A2(new_n811), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n1007), .A2(new_n1013), .A3(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1003), .B1(new_n1176), .B2(new_n1008), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1178), .B(KEYINPUT48), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1006), .B(KEYINPUT46), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT47), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1182));
  XOR2_X1   g757(.A(new_n1182), .B(KEYINPUT126), .Z(new_n1183));
  NAND3_X1  g758(.A1(new_n1180), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1184), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1181), .B1(new_n1180), .B2(new_n1183), .ZN(new_n1186));
  OAI221_X1 g761(.A(new_n1177), .B1(new_n1017), .B2(new_n1179), .C1(new_n1185), .C2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1174), .A2(new_n1188), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g764(.A(KEYINPUT127), .ZN(new_n1191));
  NAND2_X1  g765(.A1(new_n986), .A2(new_n988), .ZN(new_n1192));
  NAND2_X1  g766(.A1(new_n990), .A2(new_n992), .ZN(new_n1193));
  NAND2_X1  g767(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NOR4_X1   g768(.A1(G229), .A2(new_n459), .A3(new_n669), .A4(G227), .ZN(new_n1195));
  AND2_X1   g769(.A1(new_n909), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g770(.A(new_n1191), .B1(new_n1194), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g771(.A1(new_n909), .A2(new_n1195), .ZN(new_n1198));
  NOR3_X1   g772(.A1(new_n993), .A2(KEYINPUT127), .A3(new_n1198), .ZN(new_n1199));
  NOR2_X1   g773(.A1(new_n1197), .A2(new_n1199), .ZN(G308));
  NAND3_X1  g774(.A1(new_n1194), .A2(new_n1191), .A3(new_n1196), .ZN(new_n1201));
  OAI21_X1  g775(.A(KEYINPUT127), .B1(new_n993), .B2(new_n1198), .ZN(new_n1202));
  NAND2_X1  g776(.A1(new_n1201), .A2(new_n1202), .ZN(G225));
endmodule


