//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 1 1 0 1 1 1 1 0 1 0 1 1 0 0 1 1 0 1 1 1 0 0 1 0 1 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 0 0 1 0 1 1 1 1 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n541, new_n542,
    new_n544, new_n545, new_n546, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n559,
    new_n560, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n625,
    new_n627, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT66), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT67), .Z(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT68), .Z(G217));
  NOR4_X1   g026(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  OR2_X1    g030(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT69), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  AOI22_X1  g033(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n462), .A2(new_n464), .A3(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n460), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G101), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT3), .B(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n469), .B1(new_n470), .B2(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(KEYINPUT70), .B1(new_n471), .B2(G2105), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n462), .A2(new_n464), .A3(G137), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(new_n468), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT70), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n474), .A2(new_n475), .A3(new_n460), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n467), .B1(new_n472), .B2(new_n476), .ZN(G160));
  NAND2_X1  g052(.A1(new_n462), .A2(new_n464), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(new_n460), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n478), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  NAND4_X1  g061(.A1(new_n462), .A2(new_n464), .A3(G126), .A4(G2105), .ZN(new_n487));
  OR2_X1    g062(.A1(G102), .A2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n488), .A2(new_n490), .A3(G2104), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT71), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n462), .A2(new_n464), .A3(G138), .A4(new_n460), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n470), .A2(KEYINPUT4), .A3(G138), .A4(new_n460), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n487), .A2(new_n498), .A3(new_n491), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n493), .A2(new_n496), .A3(new_n497), .A4(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  AND2_X1   g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  OAI211_X1 g078(.A(G50), .B(G543), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G543), .ZN(new_n508));
  OAI211_X1 g083(.A(new_n506), .B(new_n508), .C1(new_n502), .C2(new_n503), .ZN(new_n509));
  XOR2_X1   g084(.A(KEYINPUT72), .B(G88), .Z(new_n510));
  OAI21_X1  g085(.A(new_n504), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n506), .A2(new_n508), .A3(G62), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n511), .A2(new_n515), .ZN(G166));
  OR2_X1    g091(.A1(new_n502), .A2(new_n503), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n506), .A2(new_n508), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n517), .A2(G51), .A3(G543), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XOR2_X1   g098(.A(new_n523), .B(KEYINPUT7), .Z(new_n524));
  NOR3_X1   g099(.A1(new_n520), .A2(new_n522), .A3(new_n524), .ZN(G168));
  NAND2_X1  g100(.A1(new_n517), .A2(G543), .ZN(new_n526));
  INV_X1    g101(.A(G52), .ZN(new_n527));
  INV_X1    g102(.A(G90), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n526), .A2(new_n527), .B1(new_n528), .B2(new_n509), .ZN(new_n529));
  XNOR2_X1  g104(.A(KEYINPUT5), .B(G543), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n530), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n531), .A2(new_n512), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n529), .A2(new_n532), .ZN(G171));
  XOR2_X1   g108(.A(KEYINPUT73), .B(G43), .Z(new_n534));
  INV_X1    g109(.A(G81), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n526), .A2(new_n534), .B1(new_n535), .B2(new_n509), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n530), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n512), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G860), .ZN(G153));
  AND3_X1   g115(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G36), .ZN(new_n542));
  XOR2_X1   g117(.A(new_n542), .B(KEYINPUT74), .Z(G176));
  NAND2_X1  g118(.A1(G1), .A2(G3), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT75), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n541), .A2(new_n546), .ZN(G188));
  OAI211_X1 g122(.A(G53), .B(G543), .C1(new_n502), .C2(new_n503), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT9), .ZN(new_n549));
  INV_X1    g124(.A(new_n509), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G91), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT76), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n506), .A2(new_n508), .A3(G65), .ZN(new_n553));
  NAND2_X1  g128(.A1(G78), .A2(G543), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n552), .B1(new_n555), .B2(G651), .ZN(new_n556));
  AOI211_X1 g131(.A(KEYINPUT76), .B(new_n512), .C1(new_n553), .C2(new_n554), .ZN(new_n557));
  OAI211_X1 g132(.A(new_n549), .B(new_n551), .C1(new_n556), .C2(new_n557), .ZN(G299));
  OR3_X1    g133(.A1(new_n529), .A2(new_n532), .A3(KEYINPUT77), .ZN(new_n559));
  OAI21_X1  g134(.A(KEYINPUT77), .B1(new_n529), .B2(new_n532), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(G301));
  OR3_X1    g136(.A1(new_n520), .A2(new_n522), .A3(new_n524), .ZN(G286));
  NAND2_X1  g137(.A1(new_n513), .A2(new_n514), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G651), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT78), .ZN(new_n565));
  XNOR2_X1  g140(.A(KEYINPUT72), .B(G88), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n517), .A2(new_n530), .A3(new_n566), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n564), .A2(new_n565), .A3(new_n504), .A4(new_n567), .ZN(new_n568));
  OAI21_X1  g143(.A(KEYINPUT78), .B1(new_n511), .B2(new_n515), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(G303));
  OAI21_X1  g145(.A(G651), .B1(new_n530), .B2(G74), .ZN(new_n571));
  INV_X1    g146(.A(G87), .ZN(new_n572));
  INV_X1    g147(.A(G49), .ZN(new_n573));
  OAI221_X1 g148(.A(new_n571), .B1(new_n572), .B2(new_n509), .C1(new_n526), .C2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT79), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n574), .B(new_n575), .ZN(G288));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G61), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n519), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G651), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(G48), .ZN(new_n582));
  INV_X1    g157(.A(G86), .ZN(new_n583));
  OAI22_X1  g158(.A1(new_n526), .A2(new_n582), .B1(new_n583), .B2(new_n509), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT80), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g162(.A(KEYINPUT80), .B1(new_n584), .B2(new_n581), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(G305));
  INV_X1    g164(.A(G47), .ZN(new_n590));
  INV_X1    g165(.A(G85), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n526), .A2(new_n590), .B1(new_n591), .B2(new_n509), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n530), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n593), .A2(new_n512), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G290));
  INV_X1    g171(.A(G301), .ZN(new_n597));
  INV_X1    g172(.A(G868), .ZN(new_n598));
  OR3_X1    g173(.A1(new_n597), .A2(KEYINPUT81), .A3(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(KEYINPUT81), .B1(new_n597), .B2(new_n598), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  INV_X1    g176(.A(G79), .ZN(new_n602));
  OAI22_X1  g177(.A1(new_n519), .A2(new_n601), .B1(new_n602), .B2(new_n505), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT82), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI221_X1 g180(.A(KEYINPUT82), .B1(new_n602), .B2(new_n505), .C1(new_n519), .C2(new_n601), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n605), .A2(G651), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n517), .A2(G54), .A3(G543), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n550), .A2(KEYINPUT10), .A3(G92), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  INV_X1    g185(.A(G92), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n509), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n607), .A2(new_n608), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(KEYINPUT83), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT83), .ZN(new_n616));
  NAND4_X1  g191(.A1(new_n607), .A2(new_n613), .A3(new_n616), .A4(new_n608), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n599), .B(new_n600), .C1(G868), .C2(new_n619), .ZN(G284));
  OAI211_X1 g195(.A(new_n599), .B(new_n600), .C1(G868), .C2(new_n619), .ZN(G321));
  NAND2_X1  g196(.A1(G299), .A2(new_n598), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(new_n598), .B2(G168), .ZN(G297));
  OAI21_X1  g198(.A(new_n622), .B1(new_n598), .B2(G168), .ZN(G280));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n619), .B1(new_n625), .B2(G860), .ZN(G148));
  NOR2_X1   g201(.A1(new_n618), .A2(G559), .ZN(new_n627));
  OR3_X1    g202(.A1(new_n627), .A2(KEYINPUT84), .A3(new_n598), .ZN(new_n628));
  OAI21_X1  g203(.A(KEYINPUT84), .B1(new_n627), .B2(new_n598), .ZN(new_n629));
  OAI211_X1 g204(.A(new_n628), .B(new_n629), .C1(G868), .C2(new_n539), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g206(.A1(new_n470), .A2(new_n460), .ZN(new_n632));
  OR3_X1    g207(.A1(new_n632), .A2(KEYINPUT12), .A3(new_n461), .ZN(new_n633));
  OAI21_X1  g208(.A(KEYINPUT12), .B1(new_n632), .B2(new_n461), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2100), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n481), .A2(G135), .ZN(new_n638));
  OR2_X1    g213(.A1(G99), .A2(G2105), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n639), .B(G2104), .C1(G111), .C2(new_n460), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n641), .B1(G123), .B2(new_n479), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2096), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n637), .A2(new_n643), .ZN(G156));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT86), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2427), .B(G2430), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(KEYINPUT14), .ZN(new_n650));
  XOR2_X1   g225(.A(KEYINPUT85), .B(KEYINPUT16), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2451), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2454), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n650), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2443), .B(G2446), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(G14), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(G401));
  XOR2_X1   g235(.A(G2072), .B(G2078), .Z(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n661), .B1(new_n664), .B2(KEYINPUT18), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2096), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(G2100), .Z(new_n667));
  AND2_X1   g242(.A1(new_n664), .A2(KEYINPUT17), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n662), .A2(new_n663), .ZN(new_n669));
  AOI21_X1  g244(.A(KEYINPUT18), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n667), .B(new_n670), .ZN(G227));
  XNOR2_X1  g246(.A(G1991), .B(G1996), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT88), .Z(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT87), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT19), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  AND2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT20), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n679), .A2(new_n680), .ZN(new_n684));
  AOI22_X1  g259(.A1(new_n682), .A2(new_n683), .B1(new_n678), .B2(new_n684), .ZN(new_n685));
  OR3_X1    g260(.A1(new_n678), .A2(new_n681), .A3(new_n684), .ZN(new_n686));
  OAI211_X1 g261(.A(new_n685), .B(new_n686), .C1(new_n683), .C2(new_n682), .ZN(new_n687));
  XOR2_X1   g262(.A(G1981), .B(G1986), .Z(new_n688));
  OR2_X1    g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n687), .A2(new_n688), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n689), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n691), .B1(new_n689), .B2(new_n692), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n674), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n695), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n697), .A2(new_n673), .A3(new_n693), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n698), .ZN(G229));
  NAND2_X1  g274(.A1(new_n479), .A2(G119), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n481), .A2(G131), .ZN(new_n701));
  OR2_X1    g276(.A1(G95), .A2(G2105), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n702), .B(G2104), .C1(G107), .C2(new_n460), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n700), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT89), .B(G29), .ZN(new_n705));
  MUX2_X1   g280(.A(G25), .B(new_n704), .S(new_n705), .Z(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT35), .B(G1991), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT90), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n706), .B(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G24), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(new_n595), .B2(new_n710), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n712), .A2(G1986), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n712), .A2(G1986), .ZN(new_n714));
  NOR3_X1   g289(.A1(new_n709), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n710), .B1(new_n587), .B2(new_n588), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n710), .A2(G6), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT32), .B(G1981), .Z(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  OR3_X1    g294(.A1(new_n716), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n716), .B2(new_n717), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n710), .A2(G22), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G166), .B2(new_n710), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(G1971), .Z(new_n725));
  INV_X1    g300(.A(new_n574), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G16), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G16), .B2(G23), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT33), .B(G1976), .Z(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n727), .B(new_n729), .C1(G16), .C2(G23), .ZN(new_n732));
  AND3_X1   g307(.A1(new_n725), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  AND3_X1   g308(.A1(new_n722), .A2(KEYINPUT34), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(KEYINPUT34), .B1(new_n722), .B2(new_n733), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n715), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(KEYINPUT36), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT36), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n738), .B(new_n715), .C1(new_n734), .C2(new_n735), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(G171), .A2(G16), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G5), .B2(G16), .ZN(new_n742));
  INV_X1    g317(.A(G1961), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OR2_X1    g319(.A1(G29), .A2(G32), .ZN(new_n745));
  NAND3_X1  g320(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT26), .Z(new_n747));
  AOI22_X1  g322(.A1(new_n470), .A2(G141), .B1(G105), .B2(G2104), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n479), .A2(G129), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n749), .A2(KEYINPUT94), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n749), .A2(KEYINPUT94), .ZN(new_n751));
  OAI221_X1 g326(.A(new_n747), .B1(G2105), .B2(new_n748), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G29), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n745), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT27), .B(G1996), .Z(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n744), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT97), .ZN(new_n758));
  NAND2_X1  g333(.A1(G160), .A2(G29), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT24), .B(G34), .Z(new_n760));
  OAI21_X1  g335(.A(new_n759), .B1(new_n705), .B2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G2084), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OR3_X1    g338(.A1(new_n757), .A2(new_n758), .A3(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(G16), .A2(G21), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G168), .B2(G16), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT95), .B(G1966), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n539), .A2(new_n710), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n710), .A2(G19), .ZN(new_n770));
  OAI21_X1  g345(.A(G1341), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OR3_X1    g346(.A1(new_n769), .A2(G1341), .A3(new_n770), .ZN(new_n772));
  XOR2_X1   g347(.A(KEYINPUT31), .B(G11), .Z(new_n773));
  INV_X1    g348(.A(KEYINPUT30), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n774), .A2(G28), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n774), .A2(G28), .ZN(new_n776));
  NOR3_X1   g351(.A1(new_n775), .A2(new_n776), .A3(G29), .ZN(new_n777));
  AOI211_X1 g352(.A(new_n773), .B(new_n777), .C1(new_n642), .C2(new_n705), .ZN(new_n778));
  AND4_X1   g353(.A1(new_n768), .A2(new_n771), .A3(new_n772), .A4(new_n778), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT91), .B(G1348), .Z(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n619), .A2(new_n710), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n710), .A2(G4), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(new_n705), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(G27), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G164), .B2(new_n785), .ZN(new_n787));
  MUX2_X1   g362(.A(new_n786), .B(new_n787), .S(KEYINPUT98), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n788), .A2(G2078), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n764), .A2(new_n779), .A3(new_n784), .A4(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(G35), .ZN(new_n791));
  OAI21_X1  g366(.A(KEYINPUT99), .B1(new_n705), .B2(new_n791), .ZN(new_n792));
  OR3_X1    g367(.A1(new_n705), .A2(KEYINPUT99), .A3(new_n791), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n792), .B(new_n793), .C1(G162), .C2(new_n785), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT29), .B(G2090), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n790), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n758), .B1(new_n757), .B2(new_n763), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n761), .A2(new_n762), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT93), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n788), .A2(G2078), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n754), .A2(new_n756), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n798), .A2(new_n800), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  NOR3_X1   g378(.A1(new_n782), .A2(new_n783), .A3(new_n781), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n479), .A2(G128), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n481), .A2(G140), .ZN(new_n806));
  OR2_X1    g381(.A1(G104), .A2(G2105), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n807), .B(G2104), .C1(G116), .C2(new_n460), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n805), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n785), .A2(G26), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n809), .A2(G29), .B1(KEYINPUT28), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(KEYINPUT28), .B2(new_n810), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G2067), .ZN(new_n813));
  NOR3_X1   g388(.A1(new_n803), .A2(new_n804), .A3(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT100), .B(KEYINPUT23), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n710), .A2(G20), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(G299), .B2(G16), .ZN(new_n818));
  INV_X1    g393(.A(G1956), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  AND3_X1   g396(.A1(new_n797), .A2(new_n814), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n742), .A2(new_n743), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT96), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT25), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(G139), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n829), .B2(new_n632), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n830), .A2(KEYINPUT92), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n830), .A2(KEYINPUT92), .ZN(new_n832));
  AOI22_X1  g407(.A1(new_n470), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n833));
  OAI22_X1  g408(.A1(new_n831), .A2(new_n832), .B1(new_n460), .B2(new_n833), .ZN(new_n834));
  MUX2_X1   g409(.A(G33), .B(new_n834), .S(G29), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(G2072), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n740), .A2(new_n822), .A3(new_n825), .A4(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(G311));
  NAND2_X1  g414(.A1(new_n838), .A2(KEYINPUT101), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n797), .A2(new_n814), .A3(new_n821), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(new_n737), .B2(new_n739), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT101), .ZN(new_n843));
  NAND4_X1  g418(.A1(new_n842), .A2(new_n843), .A3(new_n825), .A4(new_n837), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n840), .A2(new_n844), .ZN(G150));
  INV_X1    g420(.A(G55), .ZN(new_n846));
  INV_X1    g421(.A(G93), .ZN(new_n847));
  OAI22_X1  g422(.A1(new_n526), .A2(new_n846), .B1(new_n847), .B2(new_n509), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n530), .A2(G67), .ZN(new_n849));
  NAND2_X1  g424(.A1(G80), .A2(G543), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n512), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(G860), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT37), .Z(new_n855));
  NOR2_X1   g430(.A1(new_n618), .A2(new_n625), .ZN(new_n856));
  XOR2_X1   g431(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  OR3_X1    g433(.A1(new_n848), .A2(KEYINPUT102), .A3(new_n851), .ZN(new_n859));
  OAI21_X1  g434(.A(KEYINPUT102), .B1(new_n848), .B2(new_n851), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n539), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n859), .A2(new_n539), .A3(new_n860), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n858), .B(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n855), .B1(new_n865), .B2(G860), .ZN(G145));
  AND4_X1   g441(.A1(new_n496), .A2(new_n497), .A3(new_n487), .A4(new_n491), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n809), .B(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n752), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n834), .B(KEYINPUT104), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n479), .A2(G130), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n481), .A2(G142), .ZN(new_n873));
  NOR2_X1   g448(.A1(G106), .A2(G2105), .ZN(new_n874));
  OAI21_X1  g449(.A(G2104), .B1(new_n460), .B2(G118), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n872), .B(new_n873), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n635), .B(new_n876), .Z(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n704), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n878), .A2(KEYINPUT105), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n871), .B(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n485), .B(KEYINPUT103), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n881), .B(new_n642), .Z(new_n882));
  XOR2_X1   g457(.A(new_n882), .B(G160), .Z(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(G37), .B1(new_n880), .B2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n871), .B(new_n878), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(new_n883), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g464(.A1(new_n853), .A2(G868), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n614), .B(G299), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(KEYINPUT106), .ZN(new_n892));
  INV_X1    g467(.A(new_n863), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n893), .A2(new_n861), .ZN(new_n894));
  AND2_X1   g469(.A1(new_n894), .A2(new_n627), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n894), .A2(new_n627), .ZN(new_n896));
  OR3_X1    g471(.A1(new_n892), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n891), .B(KEYINPUT41), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n898), .B1(new_n895), .B2(new_n896), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(G305), .A2(KEYINPUT107), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT107), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n587), .A2(new_n903), .A3(new_n588), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n564), .A2(new_n504), .A3(new_n567), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n574), .B(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(G290), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n726), .A2(new_n906), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n574), .A2(G166), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n595), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n905), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n902), .A2(new_n908), .A3(new_n911), .A4(new_n904), .ZN(new_n914));
  AOI21_X1  g489(.A(KEYINPUT108), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n913), .A2(new_n914), .A3(KEYINPUT108), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT42), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n913), .A2(new_n914), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n901), .B(new_n919), .C1(KEYINPUT42), .C2(new_n920), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n918), .A2(KEYINPUT42), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n920), .A2(KEYINPUT42), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n900), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n921), .A2(new_n924), .A3(KEYINPUT109), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT109), .ZN(new_n926));
  OAI211_X1 g501(.A(new_n926), .B(new_n900), .C1(new_n922), .C2(new_n923), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n890), .B1(new_n928), .B2(G868), .ZN(G295));
  AOI21_X1  g504(.A(new_n890), .B1(new_n928), .B2(G868), .ZN(G331));
  AOI21_X1  g505(.A(G286), .B1(new_n559), .B2(new_n560), .ZN(new_n931));
  INV_X1    g506(.A(G171), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n932), .A2(G168), .ZN(new_n933));
  OAI22_X1  g508(.A1(new_n893), .A2(new_n861), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(G301), .A2(G168), .ZN(new_n935));
  INV_X1    g510(.A(new_n933), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n862), .A2(new_n935), .A3(new_n936), .A4(new_n863), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT110), .B1(new_n934), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT110), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n935), .A2(new_n936), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n939), .B1(new_n864), .B2(new_n940), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n938), .A2(new_n941), .A3(new_n891), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n934), .A2(new_n937), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n898), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n917), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n947), .A2(new_n915), .ZN(new_n948));
  AOI21_X1  g523(.A(G37), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n898), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n943), .A2(new_n939), .ZN(new_n951));
  INV_X1    g526(.A(new_n941), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n892), .A2(new_n943), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n918), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n949), .A2(KEYINPUT43), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT111), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n957), .B1(new_n942), .B2(new_n945), .ZN(new_n958));
  INV_X1    g533(.A(new_n891), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n951), .A2(new_n959), .A3(new_n952), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n960), .A2(KEYINPUT111), .A3(new_n944), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n958), .A2(new_n961), .A3(new_n918), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT43), .B1(new_n962), .B2(new_n949), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT44), .B1(new_n956), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT44), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT43), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n966), .B1(new_n962), .B2(new_n949), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n948), .A2(new_n944), .A3(new_n960), .ZN(new_n968));
  INV_X1    g543(.A(G37), .ZN(new_n969));
  AND4_X1   g544(.A1(new_n966), .A2(new_n955), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n965), .B1(new_n967), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n964), .A2(new_n971), .ZN(G397));
  NAND4_X1  g547(.A1(new_n496), .A2(new_n497), .A3(new_n487), .A4(new_n491), .ZN(new_n973));
  INV_X1    g548(.A(G1384), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT45), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n467), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n475), .B1(new_n474), .B2(new_n460), .ZN(new_n979));
  AOI211_X1 g554(.A(KEYINPUT70), .B(G2105), .C1(new_n473), .C2(new_n468), .ZN(new_n980));
  OAI211_X1 g555(.A(G40), .B(new_n978), .C1(new_n979), .C2(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n977), .A2(new_n981), .ZN(new_n982));
  OR2_X1    g557(.A1(new_n982), .A2(KEYINPUT112), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(KEYINPUT112), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OR2_X1    g560(.A1(new_n752), .A2(G1996), .ZN(new_n986));
  INV_X1    g561(.A(G2067), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n809), .B(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n752), .A2(G1996), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n986), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n704), .A2(new_n707), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n704), .A2(new_n707), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n990), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G1986), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n993), .B1(new_n994), .B2(new_n595), .ZN(new_n995));
  NOR2_X1   g570(.A1(G290), .A2(G1986), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n985), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n500), .A2(KEYINPUT45), .A3(new_n974), .ZN(new_n998));
  INV_X1    g573(.A(G40), .ZN(new_n999));
  AOI211_X1 g574(.A(new_n999), .B(new_n467), .C1(new_n472), .C2(new_n476), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n998), .A2(new_n1000), .A3(new_n977), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n767), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT119), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT50), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n973), .A2(new_n1005), .A3(new_n974), .ZN(new_n1006));
  NAND3_X1  g581(.A1(G160), .A2(new_n1006), .A3(G40), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n500), .A2(new_n974), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(KEYINPUT50), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1008), .A2(new_n762), .A3(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1001), .A2(KEYINPUT119), .A3(new_n767), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1004), .A2(G168), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(G8), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT51), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT62), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT51), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1004), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1017), .B1(new_n1018), .B2(G286), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1015), .B(new_n1016), .C1(new_n1014), .C2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g595(.A(KEYINPUT114), .B(KEYINPUT55), .Z(new_n1021));
  AOI21_X1  g596(.A(new_n1021), .B1(G303), .B2(G8), .ZN(new_n1022));
  INV_X1    g597(.A(G8), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT114), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1024), .A2(KEYINPUT55), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  AOI211_X1 g601(.A(new_n1023), .B(new_n1026), .C1(new_n568), .C2(new_n569), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1022), .A2(new_n1027), .ZN(new_n1028));
  XOR2_X1   g603(.A(KEYINPUT113), .B(G1971), .Z(new_n1029));
  NAND3_X1  g604(.A1(new_n973), .A2(KEYINPUT45), .A3(new_n974), .ZN(new_n1030));
  AND3_X1   g605(.A1(G160), .A2(new_n1030), .A3(G40), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1009), .A2(new_n976), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1029), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1005), .B1(new_n500), .B2(new_n974), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n1007), .A2(new_n1034), .A3(G2090), .ZN(new_n1035));
  OAI211_X1 g610(.A(G8), .B(new_n1028), .C1(new_n1033), .C2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G2090), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1008), .A2(new_n1039), .A3(new_n1010), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1029), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1000), .A2(new_n1030), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT45), .B1(new_n500), .B2(new_n974), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1041), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1040), .A2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1045), .A2(KEYINPUT115), .A3(G8), .A4(new_n1028), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1038), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n500), .A2(new_n1005), .A3(new_n974), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n975), .A2(KEYINPUT50), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1048), .A2(new_n1000), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n1039), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1005), .B1(new_n973), .B2(new_n974), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n981), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1049), .B1(new_n1054), .B2(new_n1048), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1044), .B1(new_n1052), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(G8), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1028), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  XOR2_X1   g634(.A(KEYINPUT116), .B(G1981), .Z(new_n1060));
  NAND2_X1  g635(.A1(new_n585), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G1981), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1061), .B1(new_n585), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT49), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n981), .A2(new_n975), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1066), .A2(new_n1023), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1061), .B(KEYINPUT49), .C1(new_n585), .C2(new_n1062), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1065), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G1976), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT52), .B1(G288), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n726), .A2(G1976), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(new_n1067), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1067), .A2(new_n1072), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT52), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1069), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G2078), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1031), .A2(new_n1078), .A3(new_n1032), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1010), .A2(new_n1000), .A3(new_n1006), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n1079), .A2(new_n1080), .B1(new_n1081), .B2(new_n743), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1078), .A2(KEYINPUT53), .ZN(new_n1083));
  OR2_X1    g658(.A1(new_n1001), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(G301), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  AND4_X1   g660(.A1(new_n1047), .A2(new_n1059), .A3(new_n1077), .A4(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT124), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1020), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1087), .B1(new_n1020), .B2(new_n1086), .ZN(new_n1089));
  OR2_X1    g664(.A1(new_n1019), .A2(new_n1014), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1016), .B1(new_n1090), .B2(new_n1015), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n1088), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1047), .A2(new_n1059), .A3(new_n1077), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT122), .B1(new_n1081), .B2(new_n743), .ZN(new_n1094));
  OAI211_X1 g669(.A(KEYINPUT122), .B(new_n743), .C1(new_n1007), .C2(new_n1034), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  AND4_X1   g672(.A1(KEYINPUT53), .A2(new_n1000), .A3(new_n977), .A4(new_n1030), .ZN(new_n1098));
  XNOR2_X1  g673(.A(KEYINPUT123), .B(G2078), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1080), .A2(new_n1079), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n932), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1081), .A2(new_n743), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1102), .A2(new_n1084), .A3(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1104), .A2(new_n597), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT54), .B1(new_n1101), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1097), .A2(G301), .A3(new_n1100), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1104), .A2(new_n597), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1093), .B1(new_n1106), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT61), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT56), .B(G2072), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1048), .A2(new_n1000), .A3(new_n1050), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1113), .A2(new_n1114), .B1(new_n819), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT57), .ZN(new_n1117));
  XNOR2_X1  g692(.A(G299), .B(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1112), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT121), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1115), .A2(new_n819), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1031), .A2(new_n1032), .A3(new_n1114), .ZN(new_n1122));
  AOI211_X1 g697(.A(new_n1120), .B(new_n1118), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1118), .ZN(new_n1125));
  AOI21_X1  g700(.A(KEYINPUT121), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1119), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1118), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1112), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1042), .A2(G1996), .A3(new_n1043), .ZN(new_n1131));
  XNOR2_X1  g706(.A(KEYINPUT58), .B(G1341), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1066), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n539), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT59), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT59), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1136), .B(new_n539), .C1(new_n1131), .C2(new_n1133), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(G1348), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1139), .B1(new_n1007), .B2(new_n1034), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1066), .A2(new_n987), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  OAI211_X1 g718(.A(KEYINPUT60), .B(new_n619), .C1(new_n1141), .C2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT60), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n618), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n615), .A2(KEYINPUT60), .A3(new_n617), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1146), .A2(new_n1142), .A3(new_n1140), .A4(new_n1147), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1144), .A2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1127), .A2(new_n1130), .A3(new_n1138), .A4(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n619), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1151), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1152), .B1(new_n1125), .B2(new_n1124), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1150), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1090), .A2(new_n1015), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1111), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1047), .A2(new_n1076), .ZN(new_n1157));
  XOR2_X1   g732(.A(new_n1067), .B(KEYINPUT117), .Z(new_n1158));
  INV_X1    g733(.A(G288), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1069), .A2(new_n1070), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1158), .B1(new_n1160), .B2(new_n1061), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1157), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT63), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1018), .A2(G8), .A3(G168), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1163), .B1(new_n1093), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1045), .A2(G8), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1163), .B1(new_n1167), .B2(new_n1058), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1164), .A2(new_n1047), .A3(new_n1077), .A4(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT120), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1076), .B1(new_n1038), .B2(new_n1046), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1172), .A2(KEYINPUT120), .A3(new_n1164), .A4(new_n1168), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1166), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1156), .A2(new_n1162), .A3(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n997), .B1(new_n1092), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(new_n985), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT46), .ZN(new_n1178));
  OR3_X1    g753(.A1(new_n1177), .A2(new_n1178), .A3(G1996), .ZN(new_n1179));
  INV_X1    g754(.A(new_n988), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n985), .B1(new_n752), .B2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1178), .B1(new_n1177), .B2(G1996), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1179), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT47), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n985), .A2(new_n996), .ZN(new_n1185));
  XOR2_X1   g760(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1186));
  XNOR2_X1  g761(.A(new_n1185), .B(new_n1186), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1187), .B1(new_n1177), .B2(new_n993), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n809), .A2(G2067), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n985), .A2(new_n990), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1189), .B1(new_n1190), .B2(new_n991), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n1191), .B(KEYINPUT125), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1192), .A2(new_n985), .ZN(new_n1193));
  AND3_X1   g768(.A1(new_n1184), .A2(new_n1188), .A3(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1176), .A2(new_n1194), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g770(.A(G319), .ZN(new_n1197));
  OR2_X1    g771(.A1(G227), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g772(.A(KEYINPUT127), .ZN(new_n1199));
  NAND2_X1  g773(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  OAI211_X1 g774(.A(new_n659), .B(new_n1200), .C1(new_n967), .C2(new_n970), .ZN(new_n1201));
  OR2_X1    g775(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1202));
  NAND4_X1  g776(.A1(new_n888), .A2(new_n698), .A3(new_n696), .A4(new_n1202), .ZN(new_n1203));
  NOR2_X1   g777(.A1(new_n1201), .A2(new_n1203), .ZN(G308));
  NAND3_X1  g778(.A1(new_n949), .A2(new_n966), .A3(new_n955), .ZN(new_n1205));
  AND2_X1   g779(.A1(new_n962), .A2(new_n949), .ZN(new_n1206));
  OAI21_X1  g780(.A(new_n1205), .B1(new_n1206), .B2(new_n966), .ZN(new_n1207));
  NAND3_X1  g781(.A1(new_n1202), .A2(new_n696), .A3(new_n698), .ZN(new_n1208));
  AOI21_X1  g782(.A(new_n1208), .B1(new_n885), .B2(new_n887), .ZN(new_n1209));
  NAND4_X1  g783(.A1(new_n1207), .A2(new_n659), .A3(new_n1209), .A4(new_n1200), .ZN(G225));
endmodule


