//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 1 1 0 1 1 1 0 0 0 1 0 0 0 0 0 0 0 1 0 0 1 0 1 0 1 0 0 1 1 0 1 0 0 1 0 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n809, new_n810, new_n811, new_n813, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n887, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n987, new_n988,
    new_n989, new_n990;
  XNOR2_X1  g000(.A(G64gat), .B(G92gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT80), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G8gat), .ZN(new_n204));
  INV_X1    g003(.A(G36gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G226gat), .A2(G233gat), .ZN(new_n207));
  XOR2_X1   g006(.A(new_n207), .B(KEYINPUT79), .Z(new_n208));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT69), .ZN(new_n212));
  NAND2_X1  g011(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n213), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT69), .B1(new_n215), .B2(new_n210), .ZN(new_n216));
  AOI21_X1  g015(.A(G190gat), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT28), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n209), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT68), .B(G183gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT27), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n211), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G190gat), .ZN(new_n223));
  AND3_X1   g022(.A1(new_n222), .A2(new_n218), .A3(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT26), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n229));
  AND3_X1   g028(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NOR3_X1   g029(.A1(new_n219), .A2(new_n224), .A3(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT65), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(new_n225), .B2(KEYINPUT23), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT23), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n234), .B(KEYINPUT65), .C1(G169gat), .C2(G176gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n225), .A2(KEYINPUT23), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(new_n237), .A3(new_n228), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(KEYINPUT66), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n236), .A2(new_n240), .A3(new_n237), .A4(new_n228), .ZN(new_n241));
  AND3_X1   g040(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(G183gat), .A2(G190gat), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT64), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT64), .ZN(new_n248));
  NOR4_X1   g047(.A1(new_n242), .A2(new_n243), .A3(new_n245), .A4(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n239), .A2(new_n241), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT25), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AND2_X1   g052(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n254));
  NOR2_X1   g053(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n223), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n252), .B1(new_n244), .B2(new_n256), .ZN(new_n257));
  XOR2_X1   g056(.A(new_n228), .B(KEYINPUT67), .Z(new_n258));
  NAND4_X1  g057(.A1(new_n257), .A2(new_n237), .A3(new_n236), .A4(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n231), .B1(new_n253), .B2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n208), .B1(new_n260), .B2(KEYINPUT29), .ZN(new_n261));
  INV_X1    g060(.A(G211gat), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT22), .ZN(new_n263));
  AND2_X1   g062(.A1(KEYINPUT77), .A2(G218gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(KEYINPUT77), .A2(G218gat), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G197gat), .B(G204gat), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n262), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(G204gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(G197gat), .ZN(new_n270));
  INV_X1    g069(.A(G197gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(G204gat), .ZN(new_n272));
  AND4_X1   g071(.A1(KEYINPUT22), .A2(new_n270), .A3(new_n272), .A4(new_n262), .ZN(new_n273));
  OAI21_X1  g072(.A(G218gat), .B1(new_n268), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT77), .ZN(new_n275));
  INV_X1    g074(.A(G218gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(KEYINPUT77), .A2(G218gat), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT22), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n270), .A2(new_n272), .ZN(new_n280));
  OAI21_X1  g079(.A(G211gat), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n267), .A2(KEYINPUT22), .A3(new_n262), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n281), .A2(new_n276), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n274), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT78), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n274), .A2(new_n283), .A3(KEYINPUT78), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n208), .ZN(new_n289));
  INV_X1    g088(.A(new_n259), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n290), .B1(new_n251), .B2(new_n252), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n289), .B1(new_n291), .B2(new_n231), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n261), .A2(new_n288), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n288), .B1(new_n261), .B2(new_n292), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n206), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n261), .A2(new_n292), .ZN(new_n296));
  INV_X1    g095(.A(new_n288), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n206), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n261), .A2(new_n288), .A3(new_n292), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n295), .A2(new_n301), .A3(KEYINPUT30), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT30), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n303), .B(new_n206), .C1(new_n293), .C2(new_n294), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT2), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT81), .ZN(new_n308));
  OR2_X1    g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(new_n306), .ZN(new_n310));
  INV_X1    g109(.A(G148gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G141gat), .ZN(new_n312));
  INV_X1    g111(.A(G141gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(G148gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT81), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n306), .A2(new_n316), .A3(KEYINPUT2), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n308), .A2(new_n310), .A3(new_n315), .A4(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G141gat), .B(G148gat), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n306), .B(new_n309), .C1(new_n319), .C2(KEYINPUT2), .ZN(new_n320));
  AND2_X1   g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT3), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT1), .ZN(new_n324));
  OR2_X1    g123(.A1(new_n324), .A2(KEYINPUT72), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(KEYINPUT72), .ZN(new_n326));
  OR2_X1    g125(.A1(G127gat), .A2(G134gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(G127gat), .A2(G134gat), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n325), .A2(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(G120gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(G113gat), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT71), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G113gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(G120gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n330), .A2(KEYINPUT71), .A3(G113gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n333), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n329), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n335), .A2(new_n331), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(new_n324), .ZN(new_n340));
  AND2_X1   g139(.A1(G127gat), .A2(G134gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(G127gat), .A2(G134gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT70), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT1), .B1(new_n335), .B2(new_n331), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n327), .A2(new_n328), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT70), .ZN(new_n347));
  NOR3_X1   g146(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n338), .B1(new_n344), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n318), .A2(new_n320), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT3), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n323), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT4), .ZN(new_n353));
  NAND2_X1  g152(.A1(G225gat), .A2(G233gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(KEYINPUT82), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n347), .B1(new_n345), .B2(new_n346), .ZN(new_n356));
  XNOR2_X1  g155(.A(G113gat), .B(G120gat), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n343), .B(KEYINPUT70), .C1(new_n357), .C2(KEYINPUT1), .ZN(new_n358));
  AOI22_X1  g157(.A1(new_n356), .A2(new_n358), .B1(new_n329), .B2(new_n337), .ZN(new_n359));
  AOI211_X1 g158(.A(new_n353), .B(new_n355), .C1(new_n359), .C2(new_n321), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n359), .A2(new_n353), .A3(new_n321), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n352), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT5), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n350), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n359), .A2(new_n321), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n364), .B1(new_n367), .B2(new_n355), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n361), .A2(KEYINPUT83), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n366), .A2(KEYINPUT4), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT83), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n359), .A2(new_n321), .A3(new_n372), .A4(new_n353), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n370), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n355), .A2(KEYINPUT5), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n374), .A2(new_n352), .A3(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT0), .B(G57gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(G85gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(G1gat), .B(G29gat), .ZN(new_n379));
  XOR2_X1   g178(.A(new_n378), .B(new_n379), .Z(new_n380));
  NAND3_X1  g179(.A1(new_n369), .A2(new_n376), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT84), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n369), .A2(new_n376), .A3(KEYINPUT84), .A4(new_n380), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT6), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n369), .A2(new_n376), .ZN(new_n387));
  XOR2_X1   g186(.A(new_n380), .B(KEYINPUT87), .Z(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n385), .A2(new_n386), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n380), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n387), .A2(KEYINPUT6), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n305), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT90), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(G227gat), .A2(G233gat), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n253), .A2(new_n259), .ZN(new_n400));
  INV_X1    g199(.A(new_n231), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n359), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NOR3_X1   g201(.A1(new_n291), .A2(new_n349), .A3(new_n231), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n399), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(KEYINPUT73), .B(G71gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n405), .B(G99gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(G15gat), .B(G43gat), .ZN(new_n407));
  XOR2_X1   g206(.A(new_n406), .B(new_n407), .Z(new_n408));
  OR2_X1    g207(.A1(new_n408), .A2(KEYINPUT74), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(KEYINPUT74), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(KEYINPUT33), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n404), .A2(KEYINPUT32), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n400), .A2(new_n359), .A3(new_n401), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n349), .B1(new_n291), .B2(new_n231), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT32), .ZN(new_n416));
  AOI22_X1  g215(.A1(new_n415), .A2(new_n399), .B1(new_n416), .B2(KEYINPUT33), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n412), .B1(new_n417), .B2(new_n408), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n413), .A2(new_n398), .A3(new_n414), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT34), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n419), .B(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT33), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n404), .B1(KEYINPUT32), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n408), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n419), .B(KEYINPUT34), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(new_n427), .A3(new_n412), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n422), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT86), .ZN(new_n430));
  INV_X1    g229(.A(G228gat), .ZN(new_n431));
  INV_X1    g230(.A(G233gat), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT29), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n323), .A2(new_n434), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n274), .A2(new_n283), .A3(KEYINPUT78), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT78), .B1(new_n274), .B2(new_n283), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n274), .A2(new_n283), .A3(new_n434), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n322), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n350), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n433), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n439), .A2(KEYINPUT85), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT85), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n274), .A2(new_n283), .A3(new_n444), .A4(new_n434), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n443), .A2(new_n322), .A3(new_n445), .ZN(new_n446));
  AOI22_X1  g245(.A1(new_n446), .A2(new_n350), .B1(new_n288), .B2(new_n435), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n442), .B1(new_n447), .B2(new_n433), .ZN(new_n448));
  INV_X1    g247(.A(G22gat), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n430), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(G78gat), .B(G106gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(KEYINPUT31), .B(G50gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n451), .B(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n446), .A2(new_n350), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n455), .A2(new_n433), .A3(new_n438), .ZN(new_n456));
  INV_X1    g255(.A(new_n442), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n456), .A2(new_n457), .A3(new_n449), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n449), .B1(new_n456), .B2(new_n457), .ZN(new_n459));
  OAI22_X1  g258(.A1(new_n450), .A2(new_n454), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n459), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n448), .A2(new_n449), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n461), .A2(new_n462), .A3(new_n430), .A4(new_n453), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT35), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n429), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n305), .A2(new_n394), .A3(KEYINPUT90), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n397), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT91), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n427), .A2(KEYINPUT75), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n471), .B(new_n418), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n464), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n387), .A2(new_n392), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n385), .A2(new_n386), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n393), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n305), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT35), .B1(new_n473), .B2(new_n477), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n397), .A2(new_n466), .A3(KEYINPUT91), .A4(new_n467), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n470), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n472), .A2(KEYINPUT36), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT76), .B1(new_n429), .B2(KEYINPUT36), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n472), .A2(KEYINPUT76), .A3(KEYINPUT36), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n305), .ZN(new_n486));
  INV_X1    g285(.A(new_n355), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n487), .B1(new_n374), .B2(new_n352), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n489), .B(KEYINPUT39), .C1(new_n355), .C2(new_n367), .ZN(new_n490));
  XOR2_X1   g289(.A(KEYINPUT88), .B(KEYINPUT39), .Z(new_n491));
  NAND2_X1  g290(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT89), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n492), .A2(new_n493), .A3(new_n388), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n493), .B1(new_n492), .B2(new_n388), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n490), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT40), .ZN(new_n497));
  OR2_X1    g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n497), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n486), .A2(new_n498), .A3(new_n390), .A4(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT38), .ZN(new_n501));
  NOR3_X1   g300(.A1(new_n293), .A2(new_n294), .A3(KEYINPUT37), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT37), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n503), .B1(new_n298), .B2(new_n300), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n501), .B(new_n299), .C1(new_n502), .C2(new_n504), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n505), .A2(new_n393), .A3(new_n295), .A4(new_n391), .ZN(new_n506));
  OR2_X1    g305(.A1(new_n502), .A2(new_n504), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n501), .B1(new_n507), .B2(new_n299), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n500), .B(new_n464), .C1(new_n506), .C2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n464), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n477), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n485), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n480), .A2(new_n512), .ZN(new_n513));
  XOR2_X1   g312(.A(G57gat), .B(G64gat), .Z(new_n514));
  INV_X1    g313(.A(G71gat), .ZN(new_n515));
  INV_X1    g314(.A(G78gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(G71gat), .A2(G78gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT9), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n514), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G57gat), .B(G64gat), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n518), .B(new_n517), .C1(new_n523), .C2(new_n520), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  OR2_X1    g324(.A1(new_n525), .A2(KEYINPUT21), .ZN(new_n526));
  XNOR2_X1  g325(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n527));
  XOR2_X1   g326(.A(new_n526), .B(new_n527), .Z(new_n528));
  XNOR2_X1  g327(.A(G127gat), .B(G155gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(new_n262), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n525), .A2(KEYINPUT98), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n522), .A2(new_n524), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT98), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT21), .ZN(new_n536));
  XNOR2_X1  g335(.A(G15gat), .B(G22gat), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n537), .A2(G1gat), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(G8gat), .ZN(new_n540));
  INV_X1    g339(.A(G1gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT16), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n539), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n540), .B1(new_n539), .B2(new_n543), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n536), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(G183gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT97), .ZN(new_n549));
  INV_X1    g348(.A(G183gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n547), .B(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT97), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(G231gat), .A2(G233gat), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n549), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n555), .B1(new_n549), .B2(new_n553), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n530), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n549), .A2(new_n553), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(new_n554), .ZN(new_n561));
  INV_X1    g360(.A(new_n530), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n561), .A2(new_n556), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n528), .B1(new_n559), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n559), .A2(new_n528), .A3(new_n563), .ZN(new_n566));
  NAND2_X1  g365(.A1(G99gat), .A2(G106gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT8), .ZN(new_n568));
  NAND2_X1  g367(.A1(G85gat), .A2(G92gat), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT7), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(G85gat), .ZN(new_n572));
  INV_X1    g371(.A(G92gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n568), .A2(new_n571), .A3(new_n574), .A4(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G99gat), .B(G106gat), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT99), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n571), .A2(new_n575), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT99), .ZN(new_n581));
  AOI22_X1  g380(.A1(KEYINPUT8), .A2(new_n567), .B1(new_n572), .B2(new_n573), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n580), .A2(new_n581), .A3(new_n577), .A4(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT100), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n576), .A2(new_n585), .A3(new_n578), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n585), .B1(new_n576), .B2(new_n578), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n584), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT101), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AND3_X1   g390(.A1(new_n576), .A2(new_n585), .A3(new_n578), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n592), .A2(new_n587), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n593), .A2(KEYINPUT101), .A3(new_n584), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT93), .B1(G29gat), .B2(G36gat), .ZN(new_n596));
  NOR3_X1   g395(.A1(KEYINPUT93), .A2(G29gat), .A3(G36gat), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT14), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI211_X1 g398(.A(KEYINPUT93), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(G29gat), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n602), .A2(new_n205), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G43gat), .B(G50gat), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n605), .A2(KEYINPUT15), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n603), .B1(new_n599), .B2(new_n600), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(KEYINPUT15), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n606), .A2(KEYINPUT15), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n595), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT17), .ZN(new_n615));
  AND4_X1   g414(.A1(new_n609), .A2(new_n601), .A3(new_n610), .A4(new_n604), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n609), .B1(new_n608), .B2(new_n610), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n607), .A2(KEYINPUT17), .A3(new_n611), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n613), .B(new_n614), .C1(new_n595), .C2(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(G134gat), .B(G162gat), .Z(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G190gat), .B(G218gat), .ZN(new_n624));
  AOI21_X1  g423(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n623), .B(new_n626), .Z(new_n627));
  NAND3_X1  g426(.A1(new_n565), .A2(new_n566), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G113gat), .B(G141gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(G169gat), .B(G197gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT12), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT96), .ZN(new_n637));
  OR2_X1    g436(.A1(new_n544), .A2(new_n545), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n637), .B1(new_n638), .B2(new_n612), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n546), .B1(new_n607), .B2(new_n611), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(G229gat), .A2(G233gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT13), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n639), .A2(new_n640), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n641), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT18), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n618), .A2(new_n619), .A3(new_n546), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n638), .A2(new_n612), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n648), .A2(new_n642), .A3(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT95), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n647), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT94), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n651), .B1(new_n650), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n646), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n654), .A2(KEYINPUT18), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n636), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n650), .A2(new_n651), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(KEYINPUT18), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n650), .A2(new_n653), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(KEYINPUT95), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n654), .A2(KEYINPUT18), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n662), .A2(new_n646), .A3(new_n663), .A4(new_n635), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n657), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(G120gat), .B(G148gat), .ZN(new_n667));
  INV_X1    g466(.A(G176gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(new_n269), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT10), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n672), .B1(new_n531), .B2(new_n534), .ZN(new_n673));
  AND4_X1   g472(.A1(KEYINPUT101), .A2(new_n584), .A3(new_n586), .A4(new_n588), .ZN(new_n674));
  AOI21_X1  g473(.A(KEYINPUT101), .B1(new_n593), .B2(new_n584), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n589), .A2(new_n532), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n576), .B1(KEYINPUT102), .B2(new_n577), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT102), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n580), .A2(new_n578), .A3(new_n679), .A4(new_n582), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n532), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n677), .A2(new_n672), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n676), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(G230gat), .A2(G233gat), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n671), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n685), .ZN(new_n687));
  AOI211_X1 g486(.A(KEYINPUT103), .B(new_n687), .C1(new_n676), .C2(new_n683), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n681), .B1(new_n589), .B2(new_n532), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n690), .A2(new_n685), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n670), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  AOI211_X1 g491(.A(new_n670), .B(new_n691), .C1(new_n684), .C2(new_n685), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n666), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n513), .A2(new_n629), .A3(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT104), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n697), .A2(new_n698), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n701), .A2(new_n476), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(new_n541), .ZN(G1324gat));
  OR3_X1    g502(.A1(new_n701), .A2(KEYINPUT105), .A3(new_n305), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT105), .B1(new_n701), .B2(new_n305), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT42), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n704), .B(new_n705), .C1(new_n706), .C2(G8gat), .ZN(new_n707));
  XNOR2_X1  g506(.A(KEYINPUT16), .B(G8gat), .ZN(new_n708));
  OR4_X1    g507(.A1(new_n706), .A2(new_n701), .A3(new_n305), .A4(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n706), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n707), .A2(new_n709), .A3(new_n710), .ZN(G1325gat));
  INV_X1    g510(.A(new_n701), .ZN(new_n712));
  AOI21_X1  g511(.A(G15gat), .B1(new_n712), .B2(new_n429), .ZN(new_n713));
  OR2_X1    g512(.A1(new_n485), .A2(KEYINPUT106), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n485), .A2(KEYINPUT106), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(G15gat), .ZN(new_n718));
  XOR2_X1   g517(.A(new_n718), .B(KEYINPUT107), .Z(new_n719));
  AOI21_X1  g518(.A(new_n713), .B1(new_n712), .B2(new_n719), .ZN(G1326gat));
  NOR2_X1   g519(.A1(new_n701), .A2(new_n464), .ZN(new_n721));
  XOR2_X1   g520(.A(KEYINPUT43), .B(G22gat), .Z(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(G1327gat));
  INV_X1    g522(.A(KEYINPUT111), .ZN(new_n724));
  INV_X1    g523(.A(new_n627), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n726), .A2(KEYINPUT109), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n513), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n729));
  INV_X1    g528(.A(new_n566), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n729), .B1(new_n730), .B2(new_n564), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n565), .A2(KEYINPUT108), .A3(new_n566), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n733), .A2(new_n696), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n627), .B1(new_n480), .B2(new_n512), .ZN(new_n735));
  XNOR2_X1  g534(.A(KEYINPUT109), .B(KEYINPUT44), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n728), .B(new_n734), .C1(new_n735), .C2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT110), .ZN(new_n739));
  OR3_X1    g538(.A1(new_n738), .A2(new_n739), .A3(new_n476), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(new_n738), .B2(new_n476), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n740), .A2(G29gat), .A3(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n730), .A2(new_n564), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  AND4_X1   g543(.A1(new_n744), .A2(new_n513), .A3(new_n725), .A4(new_n696), .ZN(new_n745));
  INV_X1    g544(.A(new_n476), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n745), .A2(new_n602), .A3(new_n746), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n747), .A2(KEYINPUT45), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n747), .A2(KEYINPUT45), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n724), .B1(new_n742), .B2(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n740), .A2(G29gat), .A3(new_n741), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n752), .B(KEYINPUT111), .C1(new_n748), .C2(new_n749), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(G1328gat));
  NAND3_X1  g553(.A1(new_n745), .A2(new_n205), .A3(new_n486), .ZN(new_n755));
  XOR2_X1   g554(.A(new_n755), .B(KEYINPUT46), .Z(new_n756));
  OAI21_X1  g555(.A(G36gat), .B1(new_n738), .B2(new_n305), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(G1329gat));
  INV_X1    g557(.A(G43gat), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n745), .A2(KEYINPUT112), .A3(new_n759), .A4(new_n429), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT112), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n735), .A2(new_n759), .A3(new_n744), .A4(new_n696), .ZN(new_n762));
  INV_X1    g561(.A(new_n429), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT47), .ZN(new_n766));
  OAI21_X1  g565(.A(G43gat), .B1(new_n738), .B2(new_n716), .ZN(new_n767));
  AND3_X1   g566(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n513), .A2(new_n725), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n736), .ZN(new_n770));
  INV_X1    g569(.A(new_n485), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n770), .A2(new_n771), .A3(new_n728), .A4(new_n734), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(G43gat), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n766), .B1(new_n765), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(KEYINPUT113), .B1(new_n768), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n777));
  AOI22_X1  g576(.A1(new_n764), .A2(new_n760), .B1(new_n772), .B2(G43gat), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n776), .B(new_n777), .C1(new_n766), .C2(new_n778), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n775), .A2(new_n779), .ZN(G1330gat));
  INV_X1    g579(.A(KEYINPUT115), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n770), .A2(new_n510), .A3(new_n728), .A4(new_n734), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(G50gat), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT114), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT48), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n781), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT114), .B1(new_n782), .B2(G50gat), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n788), .A2(KEYINPUT115), .A3(KEYINPUT48), .ZN(new_n789));
  INV_X1    g588(.A(new_n783), .ZN(new_n790));
  INV_X1    g589(.A(new_n745), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n791), .A2(G50gat), .A3(new_n464), .ZN(new_n792));
  OAI22_X1  g591(.A1(new_n787), .A2(new_n789), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n785), .A2(new_n781), .A3(new_n786), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n790), .A2(new_n792), .ZN(new_n795));
  OAI21_X1  g594(.A(KEYINPUT115), .B1(new_n788), .B2(KEYINPUT48), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n793), .A2(new_n797), .ZN(G1331gat));
  AOI211_X1 g597(.A(new_n628), .B(new_n665), .C1(new_n480), .C2(new_n512), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n695), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n800), .A2(new_n476), .ZN(new_n801));
  XNOR2_X1  g600(.A(KEYINPUT116), .B(G57gat), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n801), .B(new_n802), .ZN(G1332gat));
  NOR2_X1   g602(.A1(new_n800), .A2(new_n305), .ZN(new_n804));
  NOR2_X1   g603(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n805));
  AND2_X1   g604(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n807), .B1(new_n804), .B2(new_n805), .ZN(G1333gat));
  OAI21_X1  g607(.A(new_n515), .B1(new_n800), .B2(new_n763), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n799), .A2(G71gat), .A3(new_n695), .A4(new_n717), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g611(.A1(new_n800), .A2(new_n464), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(new_n516), .ZN(G1335gat));
  INV_X1    g613(.A(new_n695), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n815), .A2(new_n665), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n770), .A2(new_n744), .A3(new_n728), .A4(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n817), .A2(new_n572), .A3(new_n476), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n735), .A2(new_n744), .A3(new_n666), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(KEYINPUT51), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT51), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n735), .A2(new_n821), .A3(new_n744), .A4(new_n666), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n820), .A2(new_n746), .A3(new_n695), .A4(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n818), .B1(new_n572), .B2(new_n823), .ZN(G1336gat));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n825));
  OAI21_X1  g624(.A(G92gat), .B1(new_n817), .B2(new_n305), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT117), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n820), .A2(new_n573), .A3(new_n695), .A4(new_n822), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n826), .B1(new_n305), .B2(new_n829), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n828), .B(new_n830), .ZN(G1337gat));
  OAI21_X1  g630(.A(G99gat), .B1(new_n817), .B2(new_n716), .ZN(new_n832));
  INV_X1    g631(.A(G99gat), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n820), .A2(new_n833), .A3(new_n695), .A4(new_n822), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n832), .B1(new_n763), .B2(new_n834), .ZN(G1338gat));
  OAI21_X1  g634(.A(G106gat), .B1(new_n817), .B2(new_n464), .ZN(new_n836));
  AOI21_X1  g635(.A(KEYINPUT53), .B1(new_n836), .B2(KEYINPUT118), .ZN(new_n837));
  INV_X1    g636(.A(G106gat), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n820), .A2(new_n838), .A3(new_n695), .A4(new_n822), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n836), .B1(new_n464), .B2(new_n839), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n837), .A2(new_n840), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n841), .A2(new_n842), .ZN(G1339gat));
  NOR3_X1   g642(.A1(new_n628), .A2(new_n695), .A3(new_n665), .ZN(new_n844));
  INV_X1    g643(.A(new_n670), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n846));
  AOI22_X1  g645(.A1(new_n595), .A2(new_n673), .B1(new_n690), .B2(new_n672), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n846), .B1(new_n847), .B2(new_n687), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n684), .A2(new_n685), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n845), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n846), .B1(new_n686), .B2(new_n688), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT55), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n693), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n850), .A2(new_n851), .A3(KEYINPUT55), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n850), .A2(new_n851), .A3(KEYINPUT119), .A4(KEYINPUT55), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n854), .A2(new_n665), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n644), .B1(new_n641), .B2(new_n645), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n642), .B1(new_n648), .B2(new_n649), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n634), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n664), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n695), .ZN(new_n864));
  AOI21_X1  g663(.A(KEYINPUT120), .B1(new_n859), .B2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n859), .A2(KEYINPUT120), .A3(new_n864), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n627), .A3(new_n867), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n857), .A2(new_n858), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n725), .A2(new_n863), .A3(new_n854), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n844), .B1(new_n871), .B2(new_n733), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n763), .A2(new_n510), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n486), .A2(new_n476), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  XOR2_X1   g675(.A(new_n876), .B(KEYINPUT121), .Z(new_n877));
  OAI21_X1  g676(.A(G113gat), .B1(new_n877), .B2(new_n666), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n872), .A2(new_n473), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n875), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(new_n334), .A3(new_n665), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n878), .A2(new_n882), .ZN(G1340gat));
  OAI21_X1  g682(.A(G120gat), .B1(new_n877), .B2(new_n815), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n881), .A2(new_n330), .A3(new_n695), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(G1341gat));
  INV_X1    g685(.A(G127gat), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n877), .A2(new_n887), .A3(new_n733), .ZN(new_n888));
  AOI21_X1  g687(.A(G127gat), .B1(new_n881), .B2(new_n743), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n888), .A2(new_n889), .ZN(G1342gat));
  OAI21_X1  g689(.A(G134gat), .B1(new_n877), .B2(new_n627), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n880), .A2(G134gat), .A3(new_n627), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT56), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n893), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n891), .A2(new_n894), .A3(new_n895), .ZN(G1343gat));
  INV_X1    g695(.A(KEYINPUT122), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n859), .A2(KEYINPUT120), .A3(new_n864), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n898), .A2(new_n865), .A3(new_n725), .ZN(new_n899));
  INV_X1    g698(.A(new_n870), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n733), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n629), .A2(new_n815), .A3(new_n666), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n464), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n897), .B1(new_n903), .B2(KEYINPUT57), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n859), .A2(new_n864), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n627), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n743), .B1(new_n870), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n510), .B1(new_n844), .B2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT57), .ZN(new_n909));
  OR2_X1    g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI211_X1 g709(.A(KEYINPUT122), .B(new_n909), .C1(new_n872), .C2(new_n464), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n904), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(new_n875), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n771), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n912), .A2(new_n665), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(G141gat), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n717), .A2(new_n913), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n903), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n313), .A3(new_n665), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(KEYINPUT58), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT58), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n916), .A2(new_n923), .A3(new_n920), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(G1344gat));
  XNOR2_X1  g724(.A(KEYINPUT124), .B(KEYINPUT59), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n903), .A2(KEYINPUT57), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n908), .A2(new_n909), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n929), .A2(new_n695), .A3(new_n914), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n926), .B1(new_n930), .B2(new_n311), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n912), .A2(new_n695), .A3(new_n914), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT123), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n311), .A2(KEYINPUT59), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n933), .B1(new_n932), .B2(new_n934), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n931), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n919), .A2(new_n311), .A3(new_n695), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(G1345gat));
  NAND3_X1  g738(.A1(new_n912), .A2(G155gat), .A3(new_n914), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n940), .A2(new_n733), .ZN(new_n941));
  AOI21_X1  g740(.A(G155gat), .B1(new_n919), .B2(new_n743), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n941), .A2(new_n942), .ZN(G1346gat));
  AOI21_X1  g742(.A(G162gat), .B1(new_n919), .B2(new_n725), .ZN(new_n944));
  AND3_X1   g743(.A1(new_n912), .A2(new_n725), .A3(new_n914), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n944), .B1(new_n945), .B2(G162gat), .ZN(G1347gat));
  NOR2_X1   g745(.A1(new_n746), .A2(new_n305), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n873), .A2(new_n874), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g747(.A(G169gat), .B1(new_n948), .B2(new_n666), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n879), .A2(new_n947), .ZN(new_n950));
  OR2_X1    g749(.A1(new_n950), .A2(G169gat), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n949), .B1(new_n951), .B2(new_n666), .ZN(G1348gat));
  INV_X1    g751(.A(new_n950), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n953), .A2(new_n668), .A3(new_n695), .ZN(new_n954));
  OAI21_X1  g753(.A(G176gat), .B1(new_n948), .B2(new_n815), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  XOR2_X1   g755(.A(new_n956), .B(KEYINPUT125), .Z(G1349gat));
  AND2_X1   g756(.A1(new_n214), .A2(new_n216), .ZN(new_n958));
  OR2_X1    g757(.A1(new_n950), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n948), .A2(new_n733), .ZN(new_n960));
  OAI22_X1  g759(.A1(new_n959), .A2(new_n744), .B1(new_n220), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g761(.A(G190gat), .B1(new_n948), .B2(new_n627), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT61), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n953), .A2(new_n223), .A3(new_n725), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(G1351gat));
  NAND2_X1  g765(.A1(new_n716), .A2(new_n947), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(new_n903), .ZN(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g769(.A(G197gat), .B1(new_n970), .B2(new_n665), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n271), .B1(new_n927), .B2(new_n928), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n967), .B(KEYINPUT126), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n973), .A2(new_n666), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n971), .B1(new_n972), .B2(new_n974), .ZN(G1352gat));
  NAND3_X1  g774(.A1(new_n970), .A2(new_n269), .A3(new_n695), .ZN(new_n976));
  OR2_X1    g775(.A1(new_n976), .A2(KEYINPUT62), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(KEYINPUT62), .ZN(new_n978));
  INV_X1    g777(.A(new_n973), .ZN(new_n979));
  AND3_X1   g778(.A1(new_n979), .A2(new_n695), .A3(new_n929), .ZN(new_n980));
  OAI211_X1 g779(.A(new_n977), .B(new_n978), .C1(new_n980), .C2(new_n269), .ZN(G1353gat));
  NAND3_X1  g780(.A1(new_n970), .A2(new_n262), .A3(new_n743), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n929), .A2(new_n743), .A3(new_n968), .ZN(new_n983));
  AND3_X1   g782(.A1(new_n983), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n984));
  AOI21_X1  g783(.A(KEYINPUT63), .B1(new_n983), .B2(G211gat), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n982), .B1(new_n984), .B2(new_n985), .ZN(G1354gat));
  AOI21_X1  g785(.A(G218gat), .B1(new_n970), .B2(new_n725), .ZN(new_n987));
  OR2_X1    g786(.A1(new_n987), .A2(KEYINPUT127), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(KEYINPUT127), .ZN(new_n989));
  AND4_X1   g788(.A1(new_n725), .A2(new_n929), .A3(new_n277), .A4(new_n278), .ZN(new_n990));
  AOI22_X1  g789(.A1(new_n988), .A2(new_n989), .B1(new_n979), .B2(new_n990), .ZN(G1355gat));
endmodule


