//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 0 0 1 1 1 0 0 1 0 0 1 1 0 0 0 1 1 1 0 1 1 1 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1 0 1 1 1 0 0 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n770, new_n771,
    new_n772, new_n774, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924;
  INV_X1    g000(.A(KEYINPUT88), .ZN(new_n202));
  XNOR2_X1  g001(.A(G78gat), .B(G106gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n203), .B(KEYINPUT86), .Z(new_n204));
  INV_X1    g003(.A(KEYINPUT87), .ZN(new_n205));
  XNOR2_X1  g004(.A(G211gat), .B(G218gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G197gat), .B(G204gat), .ZN(new_n208));
  AOI21_X1  g007(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT72), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n209), .A2(KEYINPUT72), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n207), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n212), .ZN(new_n214));
  NAND4_X1  g013(.A1(new_n214), .A2(new_n206), .A3(new_n210), .A4(new_n208), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n215), .A3(KEYINPUT73), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT73), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n217), .B(new_n207), .C1(new_n211), .C2(new_n212), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G141gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G148gat), .ZN(new_n222));
  INV_X1    g021(.A(G148gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(G141gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT78), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT2), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT78), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n222), .A2(new_n224), .A3(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n226), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G162gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G155gat), .ZN(new_n232));
  INV_X1    g031(.A(G155gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G162gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n223), .A2(KEYINPUT79), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT79), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(G148gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n236), .A2(new_n238), .A3(G141gat), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n235), .B1(new_n239), .B2(new_n222), .ZN(new_n240));
  AND2_X1   g039(.A1(KEYINPUT80), .A2(G155gat), .ZN(new_n241));
  NOR2_X1   g040(.A1(KEYINPUT80), .A2(G155gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT2), .B1(new_n243), .B2(new_n231), .ZN(new_n244));
  AOI22_X1  g043(.A1(new_n230), .A2(new_n235), .B1(new_n240), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT29), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n205), .B1(new_n220), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT29), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n216), .A2(new_n249), .A3(new_n218), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(new_n246), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n229), .A2(new_n227), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n228), .B1(new_n222), .B2(new_n224), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n235), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n240), .A2(new_n244), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n251), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(G228gat), .ZN(new_n258));
  INV_X1    g057(.A(G233gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n249), .B1(new_n256), .B2(KEYINPUT3), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n261), .A2(KEYINPUT87), .A3(new_n219), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n248), .A2(new_n257), .A3(new_n260), .A4(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n220), .A2(new_n247), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n213), .A2(new_n215), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(new_n249), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n245), .B1(new_n266), .B2(new_n246), .ZN(new_n267));
  OAI22_X1  g066(.A1(new_n264), .A2(new_n267), .B1(new_n258), .B2(new_n259), .ZN(new_n268));
  INV_X1    g067(.A(G22gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n263), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n269), .B1(new_n263), .B2(new_n268), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n204), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n263), .A2(new_n268), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(G22gat), .ZN(new_n275));
  INV_X1    g074(.A(new_n204), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n275), .A2(new_n276), .A3(new_n270), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT31), .B(G50gat), .ZN(new_n278));
  AND3_X1   g077(.A1(new_n273), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n278), .B1(new_n273), .B2(new_n277), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  XOR2_X1   g080(.A(G8gat), .B(G36gat), .Z(new_n282));
  XNOR2_X1  g081(.A(new_n282), .B(KEYINPUT76), .ZN(new_n283));
  XNOR2_X1  g082(.A(G64gat), .B(G92gat), .ZN(new_n284));
  XOR2_X1   g083(.A(new_n283), .B(new_n284), .Z(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT75), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT74), .ZN(new_n288));
  NAND2_X1  g087(.A1(G226gat), .A2(G233gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT27), .B(G183gat), .ZN(new_n290));
  INV_X1    g089(.A(G190gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  XOR2_X1   g091(.A(KEYINPUT70), .B(KEYINPUT28), .Z(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(KEYINPUT70), .A2(KEYINPUT28), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n290), .A2(new_n291), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(G183gat), .A2(G190gat), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(G169gat), .A2(G176gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NOR3_X1   g100(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n298), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n297), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT25), .ZN(new_n305));
  INV_X1    g104(.A(G183gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(new_n291), .ZN(new_n307));
  NAND3_X1  g106(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n307), .B(new_n308), .C1(new_n309), .C2(KEYINPUT65), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n309), .A2(KEYINPUT65), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(G169gat), .ZN(new_n313));
  INV_X1    g112(.A(G176gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n313), .A2(new_n314), .A3(KEYINPUT23), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT23), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n316), .B1(G169gat), .B2(G176gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n315), .A2(new_n317), .A3(new_n300), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n305), .B1(new_n312), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n298), .A2(KEYINPUT68), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT68), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n321), .A2(G183gat), .A3(G190gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT24), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n320), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT69), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n307), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(G183gat), .A2(G190gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n327), .A2(KEYINPUT69), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n324), .B(new_n308), .C1(new_n326), .C2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT67), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n300), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n315), .A2(new_n331), .A3(new_n317), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT25), .B1(new_n300), .B2(new_n330), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI22_X1  g133(.A1(new_n319), .A2(KEYINPUT66), .B1(new_n329), .B2(new_n334), .ZN(new_n335));
  AND2_X1   g134(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n327), .B1(new_n336), .B2(G190gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n298), .A2(new_n323), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT65), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n309), .A2(KEYINPUT65), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n337), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n318), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT25), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT66), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n304), .B1(new_n335), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n289), .B1(new_n347), .B2(KEYINPUT29), .ZN(new_n348));
  OR2_X1    g147(.A1(new_n297), .A2(new_n303), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n329), .A2(new_n334), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n350), .B1(new_n344), .B2(new_n345), .ZN(new_n351));
  AOI211_X1 g150(.A(KEYINPUT66), .B(KEYINPUT25), .C1(new_n342), .C2(new_n343), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n349), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n289), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n288), .B1(new_n348), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n353), .A2(new_n249), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT74), .B1(new_n357), .B2(new_n289), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n287), .B(new_n219), .C1(new_n356), .C2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n319), .A2(KEYINPUT66), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(new_n346), .A3(new_n350), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT29), .B1(new_n361), .B2(new_n349), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n355), .B1(new_n362), .B2(new_n354), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n363), .A2(new_n219), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n359), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n354), .B1(new_n353), .B2(new_n249), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n289), .B1(new_n361), .B2(new_n349), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT74), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n288), .B1(new_n362), .B2(new_n354), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n220), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n371), .A2(new_n287), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n286), .B1(new_n366), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n364), .B1(new_n371), .B2(new_n287), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n358), .B1(new_n363), .B2(KEYINPUT74), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT75), .B1(new_n375), .B2(new_n220), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n374), .A2(new_n376), .A3(KEYINPUT30), .A4(new_n285), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G1gat), .B(G29gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n379), .B(KEYINPUT0), .ZN(new_n380));
  XNOR2_X1  g179(.A(G57gat), .B(G85gat), .ZN(new_n381));
  XOR2_X1   g180(.A(new_n380), .B(new_n381), .Z(new_n382));
  INV_X1    g181(.A(KEYINPUT83), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT82), .ZN(new_n384));
  INV_X1    g183(.A(G134gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(G127gat), .ZN(new_n386));
  INV_X1    g185(.A(G127gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(G134gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G113gat), .B(G120gat), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n389), .B1(new_n390), .B2(KEYINPUT1), .ZN(new_n391));
  INV_X1    g190(.A(G120gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(G113gat), .ZN(new_n393));
  INV_X1    g192(.A(G113gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(G120gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(G127gat), .B(G134gat), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT1), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n391), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n384), .B1(new_n245), .B2(new_n400), .ZN(new_n401));
  AND4_X1   g200(.A1(new_n384), .A2(new_n400), .A3(new_n255), .A4(new_n254), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT4), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n400), .A2(new_n254), .A3(new_n255), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT4), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n400), .B1(new_n256), .B2(KEYINPUT3), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n245), .A2(new_n246), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT5), .ZN(new_n411));
  NAND2_X1  g210(.A1(G225gat), .A2(G233gat), .ZN(new_n412));
  XOR2_X1   g211(.A(new_n412), .B(KEYINPUT81), .Z(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n410), .A2(new_n411), .A3(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n383), .B1(new_n407), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n406), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n404), .A2(KEYINPUT82), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n245), .A2(new_n384), .A3(new_n400), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n417), .B1(new_n420), .B2(KEYINPUT4), .ZN(new_n421));
  AOI211_X1 g220(.A(KEYINPUT5), .B(new_n413), .C1(new_n408), .C2(new_n409), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(new_n422), .A3(KEYINPUT83), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n416), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n418), .A2(new_n419), .A3(new_n405), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n245), .A2(KEYINPUT4), .A3(new_n400), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n425), .A2(new_n410), .A3(new_n426), .A4(new_n414), .ZN(new_n427));
  INV_X1    g226(.A(new_n400), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n256), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n418), .A2(new_n419), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n411), .B1(new_n430), .B2(new_n413), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n427), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n382), .B1(new_n424), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT85), .B1(new_n433), .B2(KEYINPUT6), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n416), .A2(new_n423), .B1(new_n427), .B2(new_n431), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT85), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT6), .ZN(new_n437));
  NOR4_X1   g236(.A1(new_n435), .A2(new_n436), .A3(new_n437), .A4(new_n382), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n424), .A2(new_n382), .A3(new_n432), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT84), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n424), .A2(new_n432), .ZN(new_n442));
  INV_X1    g241(.A(new_n382), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT84), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n435), .A2(new_n445), .A3(new_n382), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n441), .A2(new_n444), .A3(new_n437), .A4(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n378), .B1(new_n439), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n374), .A2(new_n376), .A3(new_n285), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT77), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT30), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n374), .A2(new_n376), .A3(KEYINPUT77), .A4(new_n285), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n281), .B1(new_n448), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT36), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n353), .A2(new_n428), .ZN(new_n457));
  NAND2_X1  g256(.A1(G227gat), .A2(G233gat), .ZN(new_n458));
  XOR2_X1   g257(.A(new_n458), .B(KEYINPUT64), .Z(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n361), .A2(new_n400), .A3(new_n349), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n457), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n462), .B(KEYINPUT34), .ZN(new_n463));
  XOR2_X1   g262(.A(G15gat), .B(G43gat), .Z(new_n464));
  XNOR2_X1  g263(.A(G71gat), .B(G99gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n464), .B(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n460), .B1(new_n457), .B2(new_n461), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n466), .B1(new_n467), .B2(KEYINPUT33), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT32), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n457), .A2(new_n461), .ZN(new_n472));
  AOI221_X4 g271(.A(new_n469), .B1(KEYINPUT33), .B2(new_n466), .C1(new_n472), .C2(new_n459), .ZN(new_n473));
  OAI211_X1 g272(.A(KEYINPUT71), .B(new_n463), .C1(new_n471), .C2(new_n473), .ZN(new_n474));
  OR2_X1    g273(.A1(new_n468), .A2(new_n470), .ZN(new_n475));
  INV_X1    g274(.A(new_n463), .ZN(new_n476));
  INV_X1    g275(.A(new_n473), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n463), .B1(new_n471), .B2(new_n473), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n456), .B(new_n474), .C1(new_n480), .C2(KEYINPUT71), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n478), .A2(KEYINPUT36), .A3(new_n479), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n202), .B1(new_n455), .B2(new_n484), .ZN(new_n485));
  XOR2_X1   g284(.A(KEYINPUT94), .B(KEYINPUT37), .Z(new_n486));
  NAND3_X1  g285(.A1(new_n374), .A2(new_n376), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT95), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT37), .B1(new_n366), .B2(new_n372), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT95), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n374), .A2(new_n376), .A3(new_n490), .A4(new_n486), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n488), .A2(new_n286), .A3(new_n489), .A4(new_n491), .ZN(new_n492));
  XOR2_X1   g291(.A(KEYINPUT93), .B(KEYINPUT38), .Z(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AND2_X1   g293(.A1(new_n451), .A2(new_n453), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n442), .A2(KEYINPUT6), .A3(new_n443), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n436), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n433), .A2(KEYINPUT85), .A3(KEYINPUT6), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n443), .B1(new_n435), .B2(KEYINPUT90), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n424), .A2(KEYINPUT90), .A3(new_n432), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT91), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT90), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n442), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT91), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n435), .A2(KEYINPUT90), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n504), .A2(new_n505), .A3(new_n443), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n502), .A2(new_n507), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n441), .A2(new_n437), .A3(new_n446), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n499), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n220), .B1(new_n356), .B2(new_n358), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT37), .ZN(new_n512));
  INV_X1    g311(.A(new_n363), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n512), .B1(new_n513), .B2(new_n219), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n493), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n488), .A2(new_n286), .A3(new_n491), .A4(new_n515), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n494), .A2(new_n495), .A3(new_n510), .A4(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n281), .ZN(new_n518));
  INV_X1    g317(.A(new_n378), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n454), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n414), .B1(new_n421), .B2(new_n410), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n418), .A2(new_n419), .A3(new_n414), .A4(new_n429), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(KEYINPUT89), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n522), .A2(KEYINPUT39), .A3(new_n524), .ZN(new_n525));
  AND2_X1   g324(.A1(KEYINPUT92), .A2(KEYINPUT40), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT39), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n443), .B1(new_n521), .B2(new_n528), .ZN(new_n529));
  AND3_X1   g328(.A1(new_n525), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n527), .B1(new_n525), .B2(new_n529), .ZN(new_n531));
  OAI22_X1  g330(.A1(new_n530), .A2(new_n531), .B1(KEYINPUT92), .B2(KEYINPUT40), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n532), .B1(new_n502), .B2(new_n507), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n518), .B1(new_n520), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n447), .A2(new_n498), .A3(new_n497), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n454), .A2(new_n519), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(new_n518), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n538), .A2(KEYINPUT88), .A3(new_n483), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n485), .A2(new_n535), .A3(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n474), .B1(new_n480), .B2(KEYINPUT71), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT35), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n541), .A2(new_n542), .A3(new_n281), .ZN(new_n543));
  OR3_X1    g342(.A1(new_n543), .A2(new_n520), .A3(new_n510), .ZN(new_n544));
  NOR3_X1   g343(.A1(new_n480), .A2(new_n279), .A3(new_n280), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n545), .A2(new_n454), .A3(new_n536), .A4(new_n519), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT35), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n540), .A2(KEYINPUT96), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(KEYINPUT96), .B1(new_n540), .B2(new_n548), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(KEYINPUT105), .B(G92gat), .ZN(new_n552));
  INV_X1    g351(.A(G85gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(G99gat), .ZN(new_n555));
  INV_X1    g354(.A(G106gat), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT8), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT106), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(G85gat), .A2(G92gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT7), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(G99gat), .B(G106gat), .Z(new_n564));
  OR2_X1    g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n564), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G57gat), .B(G64gat), .ZN(new_n568));
  AOI21_X1  g367(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n569));
  OR2_X1    g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G71gat), .B(G78gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n567), .A2(KEYINPUT10), .A3(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n573), .A2(KEYINPUT108), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n565), .A2(new_n566), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(new_n572), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT10), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n573), .A2(KEYINPUT108), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n574), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G230gat), .A2(G233gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n582), .B1(new_n581), .B2(new_n576), .ZN(new_n583));
  XNOR2_X1  g382(.A(G120gat), .B(G148gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(G176gat), .B(G204gat), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n584), .B(new_n585), .Z(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n583), .A2(new_n587), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(G29gat), .ZN(new_n592));
  INV_X1    g391(.A(G36gat), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n592), .A2(new_n593), .A3(KEYINPUT99), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT99), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n595), .B1(G29gat), .B2(G36gat), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n594), .A2(new_n596), .A3(KEYINPUT14), .ZN(new_n597));
  NAND2_X1  g396(.A1(G29gat), .A2(G36gat), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n597), .B(new_n598), .C1(KEYINPUT14), .C2(new_n596), .ZN(new_n599));
  XOR2_X1   g398(.A(G43gat), .B(G50gat), .Z(new_n600));
  AOI21_X1  g399(.A(new_n599), .B1(KEYINPUT100), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT15), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n602), .B1(new_n599), .B2(new_n600), .ZN(new_n603));
  OR2_X1    g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n601), .A2(KEYINPUT15), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT17), .ZN(new_n607));
  XNOR2_X1  g406(.A(G15gat), .B(G22gat), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT16), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n608), .B1(new_n609), .B2(G1gat), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n610), .B1(G1gat), .B2(new_n608), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(G8gat), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n604), .A2(new_n612), .A3(new_n605), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT101), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(G229gat), .A2(G233gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(KEYINPUT102), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n619), .A2(KEYINPUT18), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n612), .B1(new_n604), .B2(new_n605), .ZN(new_n621));
  OR2_X1    g420(.A1(new_n615), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n617), .B(KEYINPUT13), .Z(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n619), .A2(KEYINPUT18), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n620), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G113gat), .B(G141gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT97), .B(KEYINPUT11), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g428(.A(G169gat), .B(G197gat), .Z(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(KEYINPUT98), .B(KEYINPUT12), .Z(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n626), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n620), .A2(new_n633), .A3(new_n624), .A4(new_n625), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n607), .A2(new_n567), .ZN(new_n638));
  XNOR2_X1  g437(.A(G190gat), .B(G218gat), .ZN(new_n639));
  AND2_X1   g438(.A1(G232gat), .A2(G233gat), .ZN(new_n640));
  AOI22_X1  g439(.A1(new_n639), .A2(KEYINPUT107), .B1(KEYINPUT41), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n641), .B1(new_n575), .B2(new_n606), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n639), .A2(KEYINPUT107), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n640), .A2(KEYINPUT41), .ZN(new_n646));
  XNOR2_X1  g445(.A(G134gat), .B(G162gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n645), .B(new_n648), .Z(new_n649));
  NOR2_X1   g448(.A1(new_n572), .A2(KEYINPUT21), .ZN(new_n650));
  XOR2_X1   g449(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n612), .B1(KEYINPUT21), .B2(new_n572), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G127gat), .B(G155gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT104), .ZN(new_n656));
  NAND2_X1  g455(.A1(G231gat), .A2(G233gat), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n657), .B(KEYINPUT103), .Z(new_n658));
  XNOR2_X1  g457(.A(new_n656), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G183gat), .B(G211gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n654), .B(new_n661), .Z(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n649), .A2(new_n663), .ZN(new_n664));
  AND3_X1   g463(.A1(new_n591), .A2(new_n637), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n551), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n536), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g469(.A1(new_n667), .A2(new_n520), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n671), .A2(G8gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT16), .B(G8gat), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT42), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n675), .B1(KEYINPUT42), .B2(new_n674), .ZN(G1325gat));
  OAI21_X1  g475(.A(G15gat), .B1(new_n666), .B2(new_n483), .ZN(new_n677));
  INV_X1    g476(.A(G15gat), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n541), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n677), .B1(new_n666), .B2(new_n679), .ZN(G1326gat));
  NOR2_X1   g479(.A1(new_n666), .A2(new_n281), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT43), .B(G22gat), .Z(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1327gat));
  NAND2_X1  g482(.A1(new_n540), .A2(new_n548), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT96), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n540), .A2(KEYINPUT96), .A3(new_n548), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n686), .A2(new_n687), .A3(new_n649), .ZN(new_n688));
  INV_X1    g487(.A(new_n637), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n689), .A2(new_n662), .A3(new_n590), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n692), .A2(new_n592), .A3(new_n668), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT45), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT109), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n546), .A2(KEYINPUT35), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n543), .A2(new_n520), .A3(new_n510), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n695), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n544), .A2(KEYINPUT109), .A3(new_n547), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n455), .A2(new_n484), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n535), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n698), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703));
  AND3_X1   g502(.A1(new_n702), .A2(new_n703), .A3(new_n649), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n649), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n549), .A2(new_n550), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n705), .B1(new_n707), .B2(new_n703), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT110), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n708), .A2(new_n709), .A3(new_n690), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n704), .B1(new_n688), .B2(KEYINPUT44), .ZN(new_n711));
  OAI21_X1  g510(.A(KEYINPUT110), .B1(new_n711), .B2(new_n691), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n713), .A2(new_n536), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n694), .B1(new_n714), .B2(new_n592), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT111), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OAI211_X1 g516(.A(KEYINPUT111), .B(new_n694), .C1(new_n714), .C2(new_n592), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(G1328gat));
  NAND2_X1  g518(.A1(new_n707), .A2(new_n690), .ZN(new_n720));
  INV_X1    g519(.A(new_n520), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n720), .A2(G36gat), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT46), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT112), .B1(new_n713), .B2(new_n721), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(G36gat), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n713), .A2(KEYINPUT112), .A3(new_n721), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n723), .B1(new_n725), .B2(new_n726), .ZN(G1329gat));
  INV_X1    g526(.A(G43gat), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n692), .A2(new_n728), .A3(new_n541), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n711), .A2(new_n483), .A3(new_n691), .ZN(new_n730));
  OAI211_X1 g529(.A(KEYINPUT47), .B(new_n729), .C1(new_n730), .C2(new_n728), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n710), .A2(new_n712), .A3(new_n484), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT113), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n732), .A2(new_n733), .A3(G43gat), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n733), .B1(new_n732), .B2(G43gat), .ZN(new_n735));
  INV_X1    g534(.A(new_n729), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n731), .B1(new_n737), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g537(.A1(new_n711), .A2(new_n281), .A3(new_n691), .ZN(new_n739));
  INV_X1    g538(.A(G50gat), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n692), .A2(KEYINPUT116), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n692), .A2(KEYINPUT116), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n281), .A2(G50gat), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI221_X1 g543(.A(KEYINPUT48), .B1(new_n739), .B2(new_n740), .C1(new_n741), .C2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n710), .A2(new_n712), .A3(new_n518), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT115), .ZN(new_n747));
  AND3_X1   g546(.A1(new_n746), .A2(new_n747), .A3(G50gat), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n747), .B1(new_n746), .B2(G50gat), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT117), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n750), .B1(new_n744), .B2(new_n741), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT116), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n720), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n753), .A2(new_n742), .A3(KEYINPUT117), .A4(new_n743), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n748), .A2(new_n749), .A3(new_n755), .ZN(new_n756));
  XOR2_X1   g555(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n757));
  OAI21_X1  g556(.A(new_n745), .B1(new_n756), .B2(new_n757), .ZN(G1331gat));
  AND3_X1   g557(.A1(new_n689), .A2(new_n664), .A3(new_n590), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n702), .A2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(new_n668), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g562(.A1(new_n760), .A2(new_n721), .ZN(new_n764));
  NOR2_X1   g563(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n765));
  AND2_X1   g564(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(new_n764), .B2(new_n765), .ZN(G1333gat));
  INV_X1    g567(.A(G71gat), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n769), .B1(new_n761), .B2(new_n484), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n541), .A2(new_n769), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n770), .B1(new_n761), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g572(.A1(new_n761), .A2(new_n518), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g574(.A1(new_n637), .A2(new_n662), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n702), .A2(new_n649), .A3(new_n776), .ZN(new_n777));
  XOR2_X1   g576(.A(new_n777), .B(KEYINPUT51), .Z(new_n778));
  AND2_X1   g577(.A1(new_n778), .A2(new_n590), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n779), .A2(new_n553), .A3(new_n668), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n708), .A2(new_n590), .A3(new_n776), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n781), .A2(new_n668), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n780), .B1(new_n782), .B2(new_n553), .ZN(G1336gat));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n520), .ZN(new_n784));
  INV_X1    g583(.A(new_n552), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n721), .A2(G92gat), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT118), .ZN(new_n788));
  AOI22_X1  g587(.A1(new_n779), .A2(new_n787), .B1(new_n788), .B2(KEYINPUT52), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  OR2_X1    g589(.A1(new_n788), .A2(KEYINPUT52), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n790), .B(new_n791), .ZN(G1337gat));
  XOR2_X1   g591(.A(KEYINPUT119), .B(G99gat), .Z(new_n793));
  NAND4_X1  g592(.A1(new_n778), .A2(new_n541), .A3(new_n590), .A4(new_n793), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n781), .A2(new_n484), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n794), .B1(new_n795), .B2(new_n793), .ZN(G1338gat));
  NOR2_X1   g595(.A1(new_n281), .A2(G106gat), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n779), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT121), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n779), .A2(KEYINPUT121), .A3(new_n797), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n556), .B1(new_n781), .B2(new_n518), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n590), .A2(new_n797), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(KEYINPUT120), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n804), .B1(new_n778), .B2(new_n806), .ZN(new_n807));
  OAI22_X1  g606(.A1(new_n803), .A2(new_n804), .B1(new_n807), .B2(new_n801), .ZN(G1339gat));
  NAND2_X1  g607(.A1(new_n582), .A2(KEYINPUT54), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n580), .A2(new_n581), .ZN(new_n810));
  OR2_X1    g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n582), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n586), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n811), .A2(KEYINPUT55), .A3(new_n814), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n817), .A2(new_n637), .A3(new_n588), .A4(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n616), .A2(new_n617), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n622), .A2(new_n623), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n631), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n590), .A2(new_n636), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n649), .B1(new_n819), .B2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n817), .A2(new_n818), .A3(new_n588), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n649), .A2(new_n636), .A3(new_n822), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n663), .B1(new_n824), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n689), .A2(new_n664), .A3(new_n591), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AND4_X1   g629(.A1(new_n668), .A2(new_n830), .A3(new_n545), .A4(new_n721), .ZN(new_n831));
  AOI21_X1  g630(.A(G113gat), .B1(new_n831), .B2(new_n637), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n518), .A2(new_n536), .ZN(new_n833));
  AND4_X1   g632(.A1(new_n721), .A2(new_n830), .A3(new_n541), .A4(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n689), .A2(new_n394), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n832), .B1(new_n834), .B2(new_n835), .ZN(G1340gat));
  AOI21_X1  g635(.A(G120gat), .B1(new_n831), .B2(new_n590), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n591), .A2(new_n392), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n837), .B1(new_n834), .B2(new_n838), .ZN(G1341gat));
  NAND3_X1  g638(.A1(new_n831), .A2(new_n387), .A3(new_n662), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n834), .A2(new_n662), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n840), .B1(new_n841), .B2(new_n387), .ZN(G1342gat));
  AND2_X1   g641(.A1(new_n834), .A2(new_n649), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n843), .A2(new_n385), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n831), .A2(new_n385), .A3(new_n649), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n844), .B1(KEYINPUT56), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n846), .B1(KEYINPUT56), .B2(new_n845), .ZN(G1343gat));
  AOI21_X1  g646(.A(new_n281), .B1(new_n828), .B2(new_n829), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n484), .A2(new_n536), .A3(new_n520), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(new_n221), .A3(new_n637), .ZN(new_n851));
  NAND2_X1  g650(.A1(KEYINPUT122), .A2(KEYINPUT58), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n848), .A2(KEYINPUT57), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n848), .A2(KEYINPUT57), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n637), .B(new_n849), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n853), .B1(G141gat), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(KEYINPUT122), .A2(KEYINPUT58), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n857), .B(new_n858), .ZN(G1344gat));
  OAI211_X1 g658(.A(new_n590), .B(new_n849), .C1(new_n854), .C2(new_n855), .ZN(new_n860));
  AOI21_X1  g659(.A(KEYINPUT59), .B1(new_n236), .B2(new_n238), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(G148gat), .ZN(new_n863));
  AOI21_X1  g662(.A(KEYINPUT123), .B1(new_n863), .B2(KEYINPUT59), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT123), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n866));
  AOI211_X1 g665(.A(new_n865), .B(new_n866), .C1(new_n860), .C2(G148gat), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n862), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n850), .A2(new_n236), .A3(new_n238), .A4(new_n590), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(G1345gat));
  OR2_X1    g669(.A1(new_n854), .A2(new_n855), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n849), .ZN(new_n872));
  OAI22_X1  g671(.A1(new_n872), .A2(new_n663), .B1(new_n242), .B2(new_n241), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n850), .A2(new_n243), .A3(new_n662), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(G1346gat));
  OAI21_X1  g674(.A(G162gat), .B1(new_n872), .B2(new_n706), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n850), .A2(new_n231), .A3(new_n649), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1347gat));
  NOR3_X1   g677(.A1(new_n721), .A2(new_n668), .A3(new_n518), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n830), .A2(new_n879), .ZN(new_n880));
  AND3_X1   g679(.A1(new_n880), .A2(new_n479), .A3(new_n478), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(new_n313), .A3(new_n637), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n541), .ZN(new_n883));
  OAI21_X1  g682(.A(G169gat), .B1(new_n883), .B2(new_n689), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  XOR2_X1   g684(.A(new_n885), .B(KEYINPUT124), .Z(G1348gat));
  AND4_X1   g685(.A1(G176gat), .A2(new_n880), .A3(new_n541), .A4(new_n590), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n881), .A2(new_n590), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n314), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n889), .A2(KEYINPUT125), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(KEYINPUT125), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n887), .B1(new_n890), .B2(new_n891), .ZN(G1349gat));
  NAND3_X1  g691(.A1(new_n881), .A2(new_n290), .A3(new_n662), .ZN(new_n893));
  OAI21_X1  g692(.A(G183gat), .B1(new_n883), .B2(new_n663), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n896));
  XOR2_X1   g695(.A(new_n895), .B(new_n896), .Z(G1350gat));
  NAND3_X1  g696(.A1(new_n881), .A2(new_n291), .A3(new_n649), .ZN(new_n898));
  OAI21_X1  g697(.A(G190gat), .B1(new_n883), .B2(new_n706), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n899), .A2(KEYINPUT61), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n899), .A2(KEYINPUT61), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(G1351gat));
  NOR3_X1   g701(.A1(new_n484), .A2(new_n721), .A3(new_n668), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n848), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(G197gat), .B1(new_n904), .B2(new_n637), .ZN(new_n905));
  XOR2_X1   g704(.A(new_n903), .B(KEYINPUT127), .Z(new_n906));
  NAND2_X1  g705(.A1(new_n871), .A2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n637), .A2(G197gat), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n905), .B1(new_n908), .B2(new_n909), .ZN(G1352gat));
  INV_X1    g709(.A(G204gat), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n904), .A2(new_n911), .A3(new_n590), .ZN(new_n912));
  XOR2_X1   g711(.A(new_n912), .B(KEYINPUT62), .Z(new_n913));
  OAI21_X1  g712(.A(G204gat), .B1(new_n907), .B2(new_n591), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(G1353gat));
  INV_X1    g714(.A(G211gat), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n904), .A2(new_n916), .A3(new_n662), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n871), .A2(new_n662), .A3(new_n906), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n918), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n919));
  AOI21_X1  g718(.A(KEYINPUT63), .B1(new_n918), .B2(G211gat), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n917), .B1(new_n919), .B2(new_n920), .ZN(G1354gat));
  OAI21_X1  g720(.A(G218gat), .B1(new_n907), .B2(new_n706), .ZN(new_n922));
  INV_X1    g721(.A(G218gat), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n904), .A2(new_n923), .A3(new_n649), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(G1355gat));
endmodule


