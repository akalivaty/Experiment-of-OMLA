

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594;

  OR2_X1 U325 ( .A1(n371), .A2(n370), .ZN(n379) );
  XNOR2_X1 U326 ( .A(n436), .B(n315), .ZN(n316) );
  XNOR2_X1 U327 ( .A(G8GAT), .B(G183GAT), .ZN(n337) );
  XOR2_X1 U328 ( .A(G176GAT), .B(G64GAT), .Z(n385) );
  XNOR2_X1 U329 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U330 ( .A(n367), .B(n322), .ZN(n323) );
  XOR2_X1 U331 ( .A(n385), .B(n384), .Z(n293) );
  OR2_X1 U332 ( .A1(n577), .A2(n440), .ZN(n294) );
  AND2_X1 U333 ( .A1(n533), .A2(n521), .ZN(n462) );
  INV_X1 U334 ( .A(n475), .ZN(n440) );
  XNOR2_X1 U335 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U336 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U337 ( .A(n302), .B(n301), .ZN(n303) );
  OR2_X1 U338 ( .A1(n576), .A2(n294), .ZN(n441) );
  XNOR2_X1 U339 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U340 ( .A(n324), .B(n323), .ZN(n326) );
  XNOR2_X1 U341 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U342 ( .A(n310), .B(n325), .Z(n585) );
  NOR2_X1 U343 ( .A1(n551), .A2(n550), .ZN(n563) );
  XNOR2_X1 U344 ( .A(n457), .B(n456), .ZN(n533) );
  XNOR2_X1 U345 ( .A(n459), .B(G176GAT), .ZN(n460) );
  XNOR2_X1 U346 ( .A(n461), .B(n460), .ZN(G1349GAT) );
  INV_X1 U347 ( .A(KEYINPUT41), .ZN(n311) );
  XOR2_X1 U348 ( .A(KEYINPUT77), .B(KEYINPUT31), .Z(n296) );
  XNOR2_X1 U349 ( .A(KEYINPUT32), .B(KEYINPUT75), .ZN(n295) );
  XNOR2_X1 U350 ( .A(n296), .B(n295), .ZN(n306) );
  XOR2_X1 U351 ( .A(KEYINPUT76), .B(n385), .Z(n298) );
  XOR2_X1 U352 ( .A(G57GAT), .B(KEYINPUT13), .Z(n334) );
  XNOR2_X1 U353 ( .A(G204GAT), .B(n334), .ZN(n297) );
  XNOR2_X1 U354 ( .A(n298), .B(n297), .ZN(n304) );
  XOR2_X1 U355 ( .A(KEYINPUT33), .B(KEYINPUT73), .Z(n300) );
  NAND2_X1 U356 ( .A1(G230GAT), .A2(G233GAT), .ZN(n299) );
  XOR2_X1 U357 ( .A(n300), .B(n299), .Z(n302) );
  XOR2_X1 U358 ( .A(G120GAT), .B(G71GAT), .Z(n454) );
  XOR2_X1 U359 ( .A(G148GAT), .B(G78GAT), .Z(n429) );
  XNOR2_X1 U360 ( .A(n454), .B(n429), .ZN(n301) );
  XNOR2_X1 U361 ( .A(n306), .B(n305), .ZN(n310) );
  XOR2_X1 U362 ( .A(KEYINPUT74), .B(G92GAT), .Z(n308) );
  XNOR2_X1 U363 ( .A(G99GAT), .B(G85GAT), .ZN(n307) );
  XNOR2_X1 U364 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U365 ( .A(G106GAT), .B(n309), .ZN(n325) );
  XNOR2_X1 U366 ( .A(n311), .B(n585), .ZN(n536) );
  XNOR2_X1 U367 ( .A(G36GAT), .B(G190GAT), .ZN(n312) );
  XNOR2_X1 U368 ( .A(n312), .B(G218GAT), .ZN(n392) );
  XOR2_X1 U369 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n314) );
  XNOR2_X1 U370 ( .A(G134GAT), .B(KEYINPUT78), .ZN(n313) );
  XNOR2_X1 U371 ( .A(n314), .B(n313), .ZN(n317) );
  XOR2_X1 U372 ( .A(G50GAT), .B(G162GAT), .Z(n436) );
  AND2_X1 U373 ( .A1(G232GAT), .A2(G233GAT), .ZN(n315) );
  XOR2_X1 U374 ( .A(n392), .B(n318), .Z(n324) );
  XOR2_X1 U375 ( .A(KEYINPUT7), .B(KEYINPUT70), .Z(n320) );
  XNOR2_X1 U376 ( .A(G43GAT), .B(G29GAT), .ZN(n319) );
  XNOR2_X1 U377 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U378 ( .A(KEYINPUT8), .B(n321), .Z(n367) );
  XNOR2_X1 U379 ( .A(KEYINPUT10), .B(KEYINPUT66), .ZN(n322) );
  XNOR2_X1 U380 ( .A(n326), .B(n325), .ZN(n374) );
  XNOR2_X1 U381 ( .A(n374), .B(KEYINPUT79), .ZN(n569) );
  XNOR2_X1 U382 ( .A(n569), .B(KEYINPUT104), .ZN(n327) );
  NAND2_X1 U383 ( .A1(n327), .A2(KEYINPUT36), .ZN(n331) );
  INV_X1 U384 ( .A(n327), .ZN(n329) );
  INV_X1 U385 ( .A(KEYINPUT36), .ZN(n328) );
  NAND2_X1 U386 ( .A1(n329), .A2(n328), .ZN(n330) );
  NAND2_X1 U387 ( .A1(n331), .A2(n330), .ZN(n490) );
  XOR2_X1 U388 ( .A(KEYINPUT15), .B(KEYINPUT81), .Z(n333) );
  XNOR2_X1 U389 ( .A(G71GAT), .B(G64GAT), .ZN(n332) );
  XNOR2_X1 U390 ( .A(n333), .B(n332), .ZN(n348) );
  XOR2_X1 U391 ( .A(n334), .B(G78GAT), .Z(n336) );
  XOR2_X1 U392 ( .A(G15GAT), .B(G127GAT), .Z(n455) );
  XNOR2_X1 U393 ( .A(n455), .B(G211GAT), .ZN(n335) );
  XNOR2_X1 U394 ( .A(n336), .B(n335), .ZN(n341) );
  XNOR2_X1 U395 ( .A(n337), .B(KEYINPUT80), .ZN(n384) );
  XOR2_X1 U396 ( .A(G22GAT), .B(G155GAT), .Z(n428) );
  XOR2_X1 U397 ( .A(n384), .B(n428), .Z(n339) );
  NAND2_X1 U398 ( .A1(G231GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U399 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U400 ( .A(n341), .B(n340), .Z(n346) );
  XOR2_X1 U401 ( .A(KEYINPUT71), .B(G1GAT), .Z(n353) );
  XOR2_X1 U402 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n343) );
  XNOR2_X1 U403 ( .A(KEYINPUT82), .B(KEYINPUT83), .ZN(n342) );
  XNOR2_X1 U404 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U405 ( .A(n353), .B(n344), .ZN(n345) );
  XNOR2_X1 U406 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U407 ( .A(n348), .B(n347), .Z(n560) );
  NAND2_X1 U408 ( .A1(n490), .A2(n560), .ZN(n350) );
  XOR2_X1 U409 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n349) );
  XNOR2_X1 U410 ( .A(n350), .B(n349), .ZN(n371) );
  XOR2_X1 U411 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n352) );
  XNOR2_X1 U412 ( .A(KEYINPUT29), .B(KEYINPUT67), .ZN(n351) );
  XNOR2_X1 U413 ( .A(n352), .B(n351), .ZN(n357) );
  XOR2_X1 U414 ( .A(G50GAT), .B(G36GAT), .Z(n355) );
  XNOR2_X1 U415 ( .A(n353), .B(KEYINPUT72), .ZN(n354) );
  XNOR2_X1 U416 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U417 ( .A(n357), .B(n356), .Z(n359) );
  NAND2_X1 U418 ( .A1(G229GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U419 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U420 ( .A(G113GAT), .B(G141GAT), .Z(n361) );
  XNOR2_X1 U421 ( .A(G197GAT), .B(G22GAT), .ZN(n360) );
  XNOR2_X1 U422 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U423 ( .A(n363), .B(n362), .Z(n369) );
  XOR2_X1 U424 ( .A(KEYINPUT69), .B(G8GAT), .Z(n365) );
  XNOR2_X1 U425 ( .A(G169GAT), .B(G15GAT), .ZN(n364) );
  XNOR2_X1 U426 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U427 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U428 ( .A(n369), .B(n368), .ZN(n580) );
  NAND2_X1 U429 ( .A1(n580), .A2(n585), .ZN(n370) );
  NOR2_X1 U430 ( .A1(n580), .A2(n536), .ZN(n372) );
  XNOR2_X1 U431 ( .A(n372), .B(KEYINPUT46), .ZN(n373) );
  NOR2_X1 U432 ( .A1(n560), .A2(n373), .ZN(n375) );
  NAND2_X1 U433 ( .A1(n375), .A2(n374), .ZN(n377) );
  XOR2_X1 U434 ( .A(KEYINPUT47), .B(KEYINPUT114), .Z(n376) );
  NAND2_X1 U435 ( .A1(n379), .A2(n378), .ZN(n381) );
  XOR2_X1 U436 ( .A(KEYINPUT48), .B(KEYINPUT64), .Z(n380) );
  XNOR2_X1 U437 ( .A(n381), .B(n380), .ZN(n530) );
  XOR2_X1 U438 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n383) );
  XNOR2_X1 U439 ( .A(G92GAT), .B(KEYINPUT95), .ZN(n382) );
  XNOR2_X1 U440 ( .A(n383), .B(n382), .ZN(n398) );
  NAND2_X1 U441 ( .A1(G226GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U442 ( .A(n293), .B(n386), .ZN(n387) );
  XOR2_X1 U443 ( .A(n387), .B(KEYINPUT94), .Z(n396) );
  XOR2_X1 U444 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n389) );
  XNOR2_X1 U445 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n388) );
  XNOR2_X1 U446 ( .A(n389), .B(n388), .ZN(n446) );
  XOR2_X1 U447 ( .A(G204GAT), .B(G211GAT), .Z(n391) );
  XNOR2_X1 U448 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n390) );
  XNOR2_X1 U449 ( .A(n391), .B(n390), .ZN(n425) );
  XNOR2_X1 U450 ( .A(n446), .B(n425), .ZN(n394) );
  XNOR2_X1 U451 ( .A(n392), .B(KEYINPUT93), .ZN(n393) );
  XNOR2_X1 U452 ( .A(n398), .B(n397), .ZN(n468) );
  NOR2_X1 U453 ( .A1(n530), .A2(n468), .ZN(n399) );
  XOR2_X1 U454 ( .A(KEYINPUT54), .B(n399), .Z(n576) );
  XOR2_X1 U455 ( .A(KEYINPUT6), .B(KEYINPUT90), .Z(n401) );
  XNOR2_X1 U456 ( .A(KEYINPUT4), .B(KEYINPUT92), .ZN(n400) );
  XNOR2_X1 U457 ( .A(n401), .B(n400), .ZN(n420) );
  XOR2_X1 U458 ( .A(G155GAT), .B(G148GAT), .Z(n403) );
  XNOR2_X1 U459 ( .A(G29GAT), .B(G127GAT), .ZN(n402) );
  XNOR2_X1 U460 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U461 ( .A(KEYINPUT5), .B(G57GAT), .Z(n405) );
  XNOR2_X1 U462 ( .A(G1GAT), .B(G120GAT), .ZN(n404) );
  XNOR2_X1 U463 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U464 ( .A(n407), .B(n406), .Z(n413) );
  XNOR2_X1 U465 ( .A(G113GAT), .B(G134GAT), .ZN(n408) );
  XNOR2_X1 U466 ( .A(n408), .B(KEYINPUT0), .ZN(n447) );
  XOR2_X1 U467 ( .A(G85GAT), .B(G162GAT), .Z(n410) );
  NAND2_X1 U468 ( .A1(G225GAT), .A2(G233GAT), .ZN(n409) );
  XNOR2_X1 U469 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U470 ( .A(n447), .B(n411), .ZN(n412) );
  XNOR2_X1 U471 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U472 ( .A(n414), .B(KEYINPUT1), .Z(n418) );
  XOR2_X1 U473 ( .A(KEYINPUT2), .B(KEYINPUT86), .Z(n416) );
  XNOR2_X1 U474 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n415) );
  XNOR2_X1 U475 ( .A(n416), .B(n415), .ZN(n424) );
  XNOR2_X1 U476 ( .A(n424), .B(KEYINPUT91), .ZN(n417) );
  XNOR2_X1 U477 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U478 ( .A(n420), .B(n419), .ZN(n577) );
  XOR2_X1 U479 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n422) );
  NAND2_X1 U480 ( .A1(G228GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U481 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U482 ( .A(n423), .B(KEYINPUT22), .Z(n427) );
  XNOR2_X1 U483 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U484 ( .A(n427), .B(n426), .ZN(n433) );
  XOR2_X1 U485 ( .A(G106GAT), .B(G218GAT), .Z(n431) );
  XNOR2_X1 U486 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U487 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U488 ( .A(n433), .B(n432), .Z(n439) );
  XOR2_X1 U489 ( .A(KEYINPUT23), .B(KEYINPUT89), .Z(n435) );
  XNOR2_X1 U490 ( .A(KEYINPUT24), .B(KEYINPUT85), .ZN(n434) );
  XNOR2_X1 U491 ( .A(n435), .B(n434), .ZN(n437) );
  XNOR2_X1 U492 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U493 ( .A(n439), .B(n438), .ZN(n475) );
  XNOR2_X1 U494 ( .A(n441), .B(KEYINPUT55), .ZN(n442) );
  XNOR2_X1 U495 ( .A(n442), .B(KEYINPUT122), .ZN(n458) );
  XOR2_X1 U496 ( .A(G176GAT), .B(G183GAT), .Z(n444) );
  NAND2_X1 U497 ( .A1(G227GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U498 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U499 ( .A(n445), .B(KEYINPUT20), .Z(n449) );
  XNOR2_X1 U500 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U501 ( .A(n449), .B(n448), .ZN(n453) );
  XOR2_X1 U502 ( .A(KEYINPUT84), .B(G190GAT), .Z(n451) );
  XNOR2_X1 U503 ( .A(G43GAT), .B(G99GAT), .ZN(n450) );
  XNOR2_X1 U504 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U505 ( .A(n453), .B(n452), .Z(n457) );
  XNOR2_X1 U506 ( .A(n455), .B(n454), .ZN(n456) );
  NAND2_X1 U507 ( .A1(n458), .A2(n533), .ZN(n568) );
  NOR2_X1 U508 ( .A1(n536), .A2(n568), .ZN(n461) );
  XNOR2_X1 U509 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n459) );
  XOR2_X1 U510 ( .A(KEYINPUT34), .B(KEYINPUT103), .Z(n482) );
  INV_X1 U511 ( .A(n468), .ZN(n521) );
  XOR2_X1 U512 ( .A(KEYINPUT100), .B(n462), .Z(n463) );
  NAND2_X1 U513 ( .A1(n463), .A2(n475), .ZN(n464) );
  XNOR2_X1 U514 ( .A(n464), .B(KEYINPUT25), .ZN(n470) );
  XNOR2_X1 U515 ( .A(KEYINPUT99), .B(KEYINPUT26), .ZN(n466) );
  NOR2_X1 U516 ( .A1(n533), .A2(n475), .ZN(n465) );
  XNOR2_X1 U517 ( .A(n466), .B(n465), .ZN(n467) );
  XOR2_X1 U518 ( .A(KEYINPUT98), .B(n467), .Z(n578) );
  INV_X1 U519 ( .A(n578), .ZN(n551) );
  XNOR2_X1 U520 ( .A(KEYINPUT27), .B(n468), .ZN(n473) );
  NOR2_X1 U521 ( .A1(n551), .A2(n473), .ZN(n469) );
  NOR2_X1 U522 ( .A1(n470), .A2(n469), .ZN(n471) );
  NOR2_X1 U523 ( .A1(n471), .A2(n577), .ZN(n472) );
  XOR2_X1 U524 ( .A(KEYINPUT101), .B(n472), .Z(n477) );
  INV_X1 U525 ( .A(n577), .ZN(n474) );
  NOR2_X1 U526 ( .A1(n474), .A2(n473), .ZN(n549) );
  XNOR2_X1 U527 ( .A(n475), .B(KEYINPUT28), .ZN(n487) );
  NAND2_X1 U528 ( .A1(n549), .A2(n487), .ZN(n531) );
  NOR2_X1 U529 ( .A1(n533), .A2(n531), .ZN(n476) );
  NOR2_X1 U530 ( .A1(n477), .A2(n476), .ZN(n491) );
  INV_X1 U531 ( .A(n560), .ZN(n589) );
  NOR2_X1 U532 ( .A1(n569), .A2(n589), .ZN(n478) );
  XOR2_X1 U533 ( .A(KEYINPUT16), .B(n478), .Z(n479) );
  NOR2_X1 U534 ( .A1(n491), .A2(n479), .ZN(n480) );
  XOR2_X1 U535 ( .A(KEYINPUT102), .B(n480), .Z(n506) );
  INV_X1 U536 ( .A(n580), .ZN(n552) );
  NAND2_X1 U537 ( .A1(n585), .A2(n552), .ZN(n495) );
  NOR2_X1 U538 ( .A1(n506), .A2(n495), .ZN(n488) );
  NAND2_X1 U539 ( .A1(n488), .A2(n577), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U541 ( .A(G1GAT), .B(n483), .ZN(G1324GAT) );
  NAND2_X1 U542 ( .A1(n488), .A2(n521), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n484), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U544 ( .A(G15GAT), .B(KEYINPUT35), .Z(n486) );
  NAND2_X1 U545 ( .A1(n488), .A2(n533), .ZN(n485) );
  XNOR2_X1 U546 ( .A(n486), .B(n485), .ZN(G1326GAT) );
  INV_X1 U547 ( .A(n487), .ZN(n525) );
  NAND2_X1 U548 ( .A1(n488), .A2(n525), .ZN(n489) );
  XNOR2_X1 U549 ( .A(n489), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U550 ( .A1(n560), .A2(n491), .ZN(n492) );
  NAND2_X1 U551 ( .A1(n490), .A2(n492), .ZN(n493) );
  XNOR2_X1 U552 ( .A(n493), .B(KEYINPUT37), .ZN(n494) );
  XNOR2_X1 U553 ( .A(KEYINPUT105), .B(n494), .ZN(n519) );
  NOR2_X1 U554 ( .A1(n519), .A2(n495), .ZN(n496) );
  XNOR2_X1 U555 ( .A(n496), .B(KEYINPUT38), .ZN(n501) );
  NAND2_X1 U556 ( .A1(n577), .A2(n501), .ZN(n498) );
  XOR2_X1 U557 ( .A(KEYINPUT106), .B(KEYINPUT39), .Z(n497) );
  XNOR2_X1 U558 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U559 ( .A(G29GAT), .B(n499), .ZN(G1328GAT) );
  NAND2_X1 U560 ( .A1(n521), .A2(n501), .ZN(n500) );
  XNOR2_X1 U561 ( .A(G36GAT), .B(n500), .ZN(G1329GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n503) );
  NAND2_X1 U563 ( .A1(n501), .A2(n533), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U565 ( .A(G43GAT), .B(n504), .ZN(G1330GAT) );
  NAND2_X1 U566 ( .A1(n525), .A2(n501), .ZN(n505) );
  XNOR2_X1 U567 ( .A(G50GAT), .B(n505), .ZN(G1331GAT) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n510) );
  XOR2_X1 U569 ( .A(KEYINPUT110), .B(KEYINPUT109), .Z(n508) );
  INV_X1 U570 ( .A(n536), .ZN(n557) );
  NAND2_X1 U571 ( .A1(n580), .A2(n557), .ZN(n518) );
  NOR2_X1 U572 ( .A1(n506), .A2(n518), .ZN(n514) );
  NAND2_X1 U573 ( .A1(n514), .A2(n577), .ZN(n507) );
  XNOR2_X1 U574 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U576 ( .A(KEYINPUT108), .B(n511), .ZN(G1332GAT) );
  NAND2_X1 U577 ( .A1(n514), .A2(n521), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n512), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U579 ( .A1(n514), .A2(n533), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n513), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT111), .B(KEYINPUT43), .Z(n516) );
  NAND2_X1 U582 ( .A1(n514), .A2(n525), .ZN(n515) );
  XNOR2_X1 U583 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U584 ( .A(G78GAT), .B(n517), .Z(G1335GAT) );
  NOR2_X1 U585 ( .A1(n519), .A2(n518), .ZN(n526) );
  NAND2_X1 U586 ( .A1(n526), .A2(n577), .ZN(n520) );
  XNOR2_X1 U587 ( .A(G85GAT), .B(n520), .ZN(G1336GAT) );
  NAND2_X1 U588 ( .A1(n526), .A2(n521), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n522), .B(KEYINPUT112), .ZN(n523) );
  XNOR2_X1 U590 ( .A(G92GAT), .B(n523), .ZN(G1337GAT) );
  NAND2_X1 U591 ( .A1(n526), .A2(n533), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n524), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT44), .B(KEYINPUT113), .Z(n528) );
  NAND2_X1 U594 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  NOR2_X1 U597 ( .A1(n530), .A2(n531), .ZN(n532) );
  NAND2_X1 U598 ( .A1(n533), .A2(n532), .ZN(n543) );
  NOR2_X1 U599 ( .A1(n580), .A2(n543), .ZN(n535) );
  XNOR2_X1 U600 ( .A(G113GAT), .B(KEYINPUT115), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n535), .B(n534), .ZN(G1340GAT) );
  NOR2_X1 U602 ( .A1(n536), .A2(n543), .ZN(n538) );
  XNOR2_X1 U603 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(G1341GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n540) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(KEYINPUT117), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(n542) );
  NOR2_X1 U608 ( .A1(n589), .A2(n543), .ZN(n541) );
  XOR2_X1 U609 ( .A(n542), .B(n541), .Z(G1342GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT51), .B(KEYINPUT118), .Z(n546) );
  INV_X1 U611 ( .A(n543), .ZN(n544) );
  NAND2_X1 U612 ( .A1(n544), .A2(n569), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U614 ( .A(G134GAT), .B(n547), .ZN(G1343GAT) );
  INV_X1 U615 ( .A(n530), .ZN(n548) );
  NAND2_X1 U616 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U617 ( .A1(n552), .A2(n563), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n553), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n555) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U622 ( .A(KEYINPUT119), .B(n556), .Z(n559) );
  NAND2_X1 U623 ( .A1(n563), .A2(n557), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(G1345GAT) );
  XOR2_X1 U625 ( .A(G155GAT), .B(KEYINPUT121), .Z(n562) );
  NAND2_X1 U626 ( .A1(n563), .A2(n560), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(G1346GAT) );
  INV_X1 U628 ( .A(n563), .ZN(n564) );
  NOR2_X1 U629 ( .A1(n374), .A2(n564), .ZN(n565) );
  XOR2_X1 U630 ( .A(G162GAT), .B(n565), .Z(G1347GAT) );
  NOR2_X1 U631 ( .A1(n580), .A2(n568), .ZN(n566) );
  XOR2_X1 U632 ( .A(G169GAT), .B(n566), .Z(G1348GAT) );
  NOR2_X1 U633 ( .A1(n589), .A2(n568), .ZN(n567) );
  XOR2_X1 U634 ( .A(G183GAT), .B(n567), .Z(G1350GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n572) );
  INV_X1 U636 ( .A(n568), .ZN(n570) );
  NAND2_X1 U637 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(G190GAT), .B(n573), .ZN(G1351GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT126), .B(KEYINPUT60), .Z(n575) );
  XNOR2_X1 U641 ( .A(KEYINPUT124), .B(KEYINPUT125), .ZN(n574) );
  XNOR2_X1 U642 ( .A(n575), .B(n574), .ZN(n584) );
  NOR2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n591) );
  NOR2_X1 U645 ( .A1(n580), .A2(n591), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(G1352GAT) );
  NOR2_X1 U649 ( .A1(n585), .A2(n591), .ZN(n587) );
  XNOR2_X1 U650 ( .A(KEYINPUT61), .B(KEYINPUT127), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(n588) );
  XOR2_X1 U652 ( .A(G204GAT), .B(n588), .Z(G1353GAT) );
  NOR2_X1 U653 ( .A1(n589), .A2(n591), .ZN(n590) );
  XOR2_X1 U654 ( .A(G211GAT), .B(n590), .Z(G1354GAT) );
  INV_X1 U655 ( .A(n591), .ZN(n592) );
  NAND2_X1 U656 ( .A1(n592), .A2(n490), .ZN(n593) );
  XNOR2_X1 U657 ( .A(n593), .B(KEYINPUT62), .ZN(n594) );
  XNOR2_X1 U658 ( .A(G218GAT), .B(n594), .ZN(G1355GAT) );
endmodule

