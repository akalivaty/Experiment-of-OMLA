

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U554 ( .A(n734), .B(KEYINPUT91), .ZN(n736) );
  XNOR2_X1 U555 ( .A(KEYINPUT1), .B(n545), .ZN(n674) );
  XNOR2_X1 U556 ( .A(n538), .B(n723), .ZN(n724) );
  AND2_X1 U557 ( .A1(n793), .A2(n791), .ZN(n734) );
  INV_X1 U558 ( .A(KEYINPUT28), .ZN(n729) );
  XNOR2_X1 U559 ( .A(n532), .B(KEYINPUT96), .ZN(n758) );
  NAND2_X1 U560 ( .A1(n535), .A2(n533), .ZN(n532) );
  XNOR2_X1 U561 ( .A(n534), .B(KEYINPUT31), .ZN(n533) );
  NAND2_X1 U562 ( .A1(n536), .A2(n519), .ZN(n535) );
  INV_X1 U563 ( .A(n736), .ZN(n722) );
  NAND2_X1 U564 ( .A1(n736), .A2(G1956), .ZN(n538) );
  XNOR2_X1 U565 ( .A(n733), .B(n537), .ZN(n536) );
  INV_X1 U566 ( .A(KEYINPUT29), .ZN(n537) );
  NAND2_X1 U567 ( .A1(n745), .A2(n744), .ZN(n534) );
  XNOR2_X1 U568 ( .A(n762), .B(n525), .ZN(n779) );
  INV_X1 U569 ( .A(KEYINPUT97), .ZN(n525) );
  NAND2_X1 U570 ( .A1(n746), .A2(G8), .ZN(n780) );
  XNOR2_X1 U571 ( .A(KEYINPUT87), .B(n707), .ZN(n791) );
  NAND2_X1 U572 ( .A1(G2105), .A2(KEYINPUT17), .ZN(n527) );
  NAND2_X1 U573 ( .A1(G2104), .A2(KEYINPUT17), .ZN(n528) );
  AND2_X1 U574 ( .A1(n784), .A2(n783), .ZN(n790) );
  NAND2_X1 U575 ( .A1(n529), .A2(n526), .ZN(n905) );
  NAND2_X1 U576 ( .A1(n531), .A2(n530), .ZN(n529) );
  AND2_X1 U577 ( .A1(n528), .A2(n527), .ZN(n526) );
  NOR2_X1 U578 ( .A1(G2104), .A2(KEYINPUT17), .ZN(n531) );
  NAND2_X1 U579 ( .A1(n905), .A2(G137), .ZN(n559) );
  OR2_X1 U580 ( .A1(G301), .A2(n743), .ZN(n519) );
  INV_X1 U581 ( .A(G2105), .ZN(n530) );
  AND2_X1 U582 ( .A1(n773), .A2(n772), .ZN(n520) );
  XNOR2_X1 U583 ( .A(n521), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U584 ( .A1(n522), .A2(n836), .ZN(n521) );
  NAND2_X1 U585 ( .A1(n523), .A2(n822), .ZN(n522) );
  NAND2_X1 U586 ( .A1(n790), .A2(n789), .ZN(n523) );
  AND2_X1 U587 ( .A1(n524), .A2(n520), .ZN(n776) );
  NAND2_X1 U588 ( .A1(n779), .A2(n768), .ZN(n524) );
  NOR2_X1 U589 ( .A1(n984), .A2(n728), .ZN(n730) );
  INV_X1 U590 ( .A(KEYINPUT94), .ZN(n723) );
  INV_X1 U591 ( .A(G651), .ZN(n543) );
  NOR2_X1 U592 ( .A1(n645), .A2(n543), .ZN(n667) );
  INV_X1 U593 ( .A(G2104), .ZN(n557) );
  XNOR2_X1 U594 ( .A(n607), .B(KEYINPUT72), .ZN(n993) );
  AND2_X1 U595 ( .A1(n530), .A2(G2104), .ZN(n904) );
  INV_X1 U596 ( .A(n993), .ZN(n846) );
  NOR2_X1 U597 ( .A1(G651), .A2(n645), .ZN(n670) );
  NOR2_X1 U598 ( .A1(n561), .A2(n560), .ZN(G160) );
  NOR2_X1 U599 ( .A1(G651), .A2(G543), .ZN(n666) );
  NAND2_X1 U600 ( .A1(n666), .A2(G89), .ZN(n539) );
  XNOR2_X1 U601 ( .A(n539), .B(KEYINPUT4), .ZN(n541) );
  XOR2_X1 U602 ( .A(KEYINPUT0), .B(G543), .Z(n645) );
  NAND2_X1 U603 ( .A1(G76), .A2(n667), .ZN(n540) );
  NAND2_X1 U604 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U605 ( .A(KEYINPUT5), .B(n542), .ZN(n551) );
  NOR2_X1 U606 ( .A1(G543), .A2(n543), .ZN(n544) );
  XOR2_X1 U607 ( .A(KEYINPUT64), .B(n544), .Z(n545) );
  NAND2_X1 U608 ( .A1(G63), .A2(n674), .ZN(n546) );
  XOR2_X1 U609 ( .A(KEYINPUT73), .B(n546), .Z(n548) );
  NAND2_X1 U610 ( .A1(n670), .A2(G51), .ZN(n547) );
  NAND2_X1 U611 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U612 ( .A(KEYINPUT6), .B(n549), .Z(n550) );
  NAND2_X1 U613 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U614 ( .A(KEYINPUT7), .B(n552), .ZN(G168) );
  XOR2_X1 U615 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  AND2_X1 U616 ( .A1(G2104), .A2(G2105), .ZN(n901) );
  NAND2_X1 U617 ( .A1(n901), .A2(G113), .ZN(n556) );
  NAND2_X1 U618 ( .A1(G2104), .A2(G101), .ZN(n553) );
  OR2_X1 U619 ( .A1(G2105), .A2(n553), .ZN(n554) );
  XOR2_X1 U620 ( .A(n554), .B(KEYINPUT23), .Z(n555) );
  NAND2_X1 U621 ( .A1(n556), .A2(n555), .ZN(n561) );
  AND2_X1 U622 ( .A1(n557), .A2(G2105), .ZN(n900) );
  NAND2_X1 U623 ( .A1(G125), .A2(n900), .ZN(n558) );
  NAND2_X1 U624 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U625 ( .A(G2443), .B(G2446), .Z(n563) );
  XNOR2_X1 U626 ( .A(G2427), .B(G2451), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n563), .B(n562), .ZN(n569) );
  XOR2_X1 U628 ( .A(G2430), .B(G2454), .Z(n565) );
  XNOR2_X1 U629 ( .A(G1341), .B(G1348), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(n567) );
  XOR2_X1 U631 ( .A(G2435), .B(G2438), .Z(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n568) );
  XOR2_X1 U633 ( .A(n569), .B(n568), .Z(n570) );
  AND2_X1 U634 ( .A1(G14), .A2(n570), .ZN(G401) );
  INV_X1 U635 ( .A(G69), .ZN(G235) );
  NAND2_X1 U636 ( .A1(n670), .A2(G52), .ZN(n572) );
  NAND2_X1 U637 ( .A1(G64), .A2(n674), .ZN(n571) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n577) );
  NAND2_X1 U639 ( .A1(G90), .A2(n666), .ZN(n574) );
  NAND2_X1 U640 ( .A1(G77), .A2(n667), .ZN(n573) );
  NAND2_X1 U641 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U642 ( .A(KEYINPUT9), .B(n575), .Z(n576) );
  NOR2_X1 U643 ( .A1(n577), .A2(n576), .ZN(G171) );
  INV_X1 U644 ( .A(G171), .ZN(G301) );
  NAND2_X1 U645 ( .A1(G102), .A2(n904), .ZN(n579) );
  NAND2_X1 U646 ( .A1(G138), .A2(n905), .ZN(n578) );
  NAND2_X1 U647 ( .A1(n579), .A2(n578), .ZN(n583) );
  NAND2_X1 U648 ( .A1(G126), .A2(n900), .ZN(n581) );
  NAND2_X1 U649 ( .A1(G114), .A2(n901), .ZN(n580) );
  NAND2_X1 U650 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U651 ( .A1(n583), .A2(n582), .ZN(G164) );
  NAND2_X1 U652 ( .A1(G94), .A2(G452), .ZN(n584) );
  XOR2_X1 U653 ( .A(KEYINPUT66), .B(n584), .Z(G173) );
  NAND2_X1 U654 ( .A1(G7), .A2(G661), .ZN(n585) );
  XOR2_X1 U655 ( .A(n585), .B(KEYINPUT10), .Z(n924) );
  NAND2_X1 U656 ( .A1(n924), .A2(G567), .ZN(n586) );
  XOR2_X1 U657 ( .A(KEYINPUT11), .B(n586), .Z(G234) );
  XOR2_X1 U658 ( .A(KEYINPUT68), .B(KEYINPUT14), .Z(n588) );
  NAND2_X1 U659 ( .A1(G56), .A2(n674), .ZN(n587) );
  XNOR2_X1 U660 ( .A(n588), .B(n587), .ZN(n595) );
  NAND2_X1 U661 ( .A1(G81), .A2(n666), .ZN(n589) );
  XOR2_X1 U662 ( .A(KEYINPUT12), .B(n589), .Z(n590) );
  XNOR2_X1 U663 ( .A(n590), .B(KEYINPUT69), .ZN(n592) );
  NAND2_X1 U664 ( .A1(G68), .A2(n667), .ZN(n591) );
  NAND2_X1 U665 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U666 ( .A(KEYINPUT13), .B(n593), .Z(n594) );
  NOR2_X1 U667 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U668 ( .A1(n670), .A2(G43), .ZN(n596) );
  NAND2_X1 U669 ( .A1(n597), .A2(n596), .ZN(n992) );
  INV_X1 U670 ( .A(G860), .ZN(n636) );
  OR2_X1 U671 ( .A1(n992), .A2(n636), .ZN(G153) );
  NAND2_X1 U672 ( .A1(G301), .A2(G868), .ZN(n598) );
  XNOR2_X1 U673 ( .A(n598), .B(KEYINPUT70), .ZN(n609) );
  INV_X1 U674 ( .A(G868), .ZN(n688) );
  NAND2_X1 U675 ( .A1(G54), .A2(n670), .ZN(n605) );
  NAND2_X1 U676 ( .A1(G79), .A2(n667), .ZN(n599) );
  XNOR2_X1 U677 ( .A(KEYINPUT71), .B(n599), .ZN(n603) );
  NAND2_X1 U678 ( .A1(G66), .A2(n674), .ZN(n601) );
  NAND2_X1 U679 ( .A1(n666), .A2(G92), .ZN(n600) );
  NAND2_X1 U680 ( .A1(n601), .A2(n600), .ZN(n602) );
  NOR2_X1 U681 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U682 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U683 ( .A(n606), .B(KEYINPUT15), .ZN(n607) );
  NAND2_X1 U684 ( .A1(n688), .A2(n846), .ZN(n608) );
  NAND2_X1 U685 ( .A1(n609), .A2(n608), .ZN(G284) );
  NAND2_X1 U686 ( .A1(n670), .A2(G53), .ZN(n611) );
  NAND2_X1 U687 ( .A1(G65), .A2(n674), .ZN(n610) );
  NAND2_X1 U688 ( .A1(n611), .A2(n610), .ZN(n615) );
  NAND2_X1 U689 ( .A1(G91), .A2(n666), .ZN(n613) );
  NAND2_X1 U690 ( .A1(G78), .A2(n667), .ZN(n612) );
  NAND2_X1 U691 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n984) );
  XNOR2_X1 U693 ( .A(n984), .B(KEYINPUT67), .ZN(G299) );
  XOR2_X1 U694 ( .A(KEYINPUT74), .B(G868), .Z(n616) );
  NOR2_X1 U695 ( .A1(G286), .A2(n616), .ZN(n619) );
  NOR2_X1 U696 ( .A1(G868), .A2(G299), .ZN(n617) );
  XOR2_X1 U697 ( .A(KEYINPUT75), .B(n617), .Z(n618) );
  NOR2_X1 U698 ( .A1(n619), .A2(n618), .ZN(G297) );
  NAND2_X1 U699 ( .A1(n636), .A2(G559), .ZN(n620) );
  NAND2_X1 U700 ( .A1(n620), .A2(n993), .ZN(n621) );
  XNOR2_X1 U701 ( .A(n621), .B(KEYINPUT76), .ZN(n622) );
  XNOR2_X1 U702 ( .A(KEYINPUT16), .B(n622), .ZN(G148) );
  NOR2_X1 U703 ( .A1(G868), .A2(n992), .ZN(n625) );
  NAND2_X1 U704 ( .A1(n993), .A2(G868), .ZN(n623) );
  NOR2_X1 U705 ( .A1(G559), .A2(n623), .ZN(n624) );
  NOR2_X1 U706 ( .A1(n625), .A2(n624), .ZN(G282) );
  NAND2_X1 U707 ( .A1(G123), .A2(n900), .ZN(n626) );
  XNOR2_X1 U708 ( .A(n626), .B(KEYINPUT18), .ZN(n629) );
  NAND2_X1 U709 ( .A1(G111), .A2(n901), .ZN(n627) );
  XOR2_X1 U710 ( .A(KEYINPUT77), .B(n627), .Z(n628) );
  NAND2_X1 U711 ( .A1(n629), .A2(n628), .ZN(n633) );
  NAND2_X1 U712 ( .A1(G99), .A2(n904), .ZN(n631) );
  NAND2_X1 U713 ( .A1(G135), .A2(n905), .ZN(n630) );
  NAND2_X1 U714 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U715 ( .A1(n633), .A2(n632), .ZN(n930) );
  XNOR2_X1 U716 ( .A(n930), .B(G2096), .ZN(n634) );
  INV_X1 U717 ( .A(G2100), .ZN(n863) );
  NAND2_X1 U718 ( .A1(n634), .A2(n863), .ZN(G156) );
  NAND2_X1 U719 ( .A1(n993), .A2(G559), .ZN(n635) );
  XOR2_X1 U720 ( .A(n992), .B(n635), .Z(n685) );
  NAND2_X1 U721 ( .A1(n636), .A2(n685), .ZN(n644) );
  NAND2_X1 U722 ( .A1(G67), .A2(n674), .ZN(n637) );
  XNOR2_X1 U723 ( .A(n637), .B(KEYINPUT78), .ZN(n639) );
  NAND2_X1 U724 ( .A1(G80), .A2(n667), .ZN(n638) );
  NAND2_X1 U725 ( .A1(n639), .A2(n638), .ZN(n643) );
  NAND2_X1 U726 ( .A1(G93), .A2(n666), .ZN(n641) );
  NAND2_X1 U727 ( .A1(G55), .A2(n670), .ZN(n640) );
  NAND2_X1 U728 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U729 ( .A1(n643), .A2(n642), .ZN(n687) );
  XOR2_X1 U730 ( .A(n644), .B(n687), .Z(G145) );
  NAND2_X1 U731 ( .A1(G87), .A2(n645), .ZN(n647) );
  NAND2_X1 U732 ( .A1(G74), .A2(G651), .ZN(n646) );
  NAND2_X1 U733 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U734 ( .A1(n674), .A2(n648), .ZN(n650) );
  NAND2_X1 U735 ( .A1(n670), .A2(G49), .ZN(n649) );
  NAND2_X1 U736 ( .A1(n650), .A2(n649), .ZN(G288) );
  NAND2_X1 U737 ( .A1(G85), .A2(n666), .ZN(n652) );
  NAND2_X1 U738 ( .A1(G72), .A2(n667), .ZN(n651) );
  NAND2_X1 U739 ( .A1(n652), .A2(n651), .ZN(n655) );
  NAND2_X1 U740 ( .A1(G60), .A2(n674), .ZN(n653) );
  XNOR2_X1 U741 ( .A(KEYINPUT65), .B(n653), .ZN(n654) );
  NOR2_X1 U742 ( .A1(n655), .A2(n654), .ZN(n657) );
  NAND2_X1 U743 ( .A1(n670), .A2(G47), .ZN(n656) );
  NAND2_X1 U744 ( .A1(n657), .A2(n656), .ZN(G290) );
  NAND2_X1 U745 ( .A1(n666), .A2(G86), .ZN(n659) );
  NAND2_X1 U746 ( .A1(G61), .A2(n674), .ZN(n658) );
  NAND2_X1 U747 ( .A1(n659), .A2(n658), .ZN(n663) );
  NAND2_X1 U748 ( .A1(G73), .A2(n667), .ZN(n660) );
  XNOR2_X1 U749 ( .A(n660), .B(KEYINPUT79), .ZN(n661) );
  XNOR2_X1 U750 ( .A(n661), .B(KEYINPUT2), .ZN(n662) );
  NOR2_X1 U751 ( .A1(n663), .A2(n662), .ZN(n665) );
  NAND2_X1 U752 ( .A1(n670), .A2(G48), .ZN(n664) );
  NAND2_X1 U753 ( .A1(n665), .A2(n664), .ZN(G305) );
  NAND2_X1 U754 ( .A1(G88), .A2(n666), .ZN(n669) );
  NAND2_X1 U755 ( .A1(G75), .A2(n667), .ZN(n668) );
  NAND2_X1 U756 ( .A1(n669), .A2(n668), .ZN(n673) );
  NAND2_X1 U757 ( .A1(n670), .A2(G50), .ZN(n671) );
  XOR2_X1 U758 ( .A(KEYINPUT80), .B(n671), .Z(n672) );
  NOR2_X1 U759 ( .A1(n673), .A2(n672), .ZN(n676) );
  NAND2_X1 U760 ( .A1(G62), .A2(n674), .ZN(n675) );
  NAND2_X1 U761 ( .A1(n676), .A2(n675), .ZN(G303) );
  XNOR2_X1 U762 ( .A(KEYINPUT82), .B(KEYINPUT19), .ZN(n678) );
  XNOR2_X1 U763 ( .A(G288), .B(KEYINPUT81), .ZN(n677) );
  XNOR2_X1 U764 ( .A(n678), .B(n677), .ZN(n681) );
  XNOR2_X1 U765 ( .A(n687), .B(G290), .ZN(n679) );
  XNOR2_X1 U766 ( .A(n679), .B(G299), .ZN(n680) );
  XNOR2_X1 U767 ( .A(n681), .B(n680), .ZN(n683) );
  XOR2_X1 U768 ( .A(G305), .B(G303), .Z(n682) );
  XNOR2_X1 U769 ( .A(n683), .B(n682), .ZN(n845) );
  XNOR2_X1 U770 ( .A(KEYINPUT83), .B(n845), .ZN(n684) );
  XNOR2_X1 U771 ( .A(n685), .B(n684), .ZN(n686) );
  NOR2_X1 U772 ( .A1(n688), .A2(n686), .ZN(n690) );
  AND2_X1 U773 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U774 ( .A1(n690), .A2(n689), .ZN(G295) );
  NAND2_X1 U775 ( .A1(G2078), .A2(G2084), .ZN(n692) );
  XOR2_X1 U776 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n691) );
  XNOR2_X1 U777 ( .A(n692), .B(n691), .ZN(n693) );
  NAND2_X1 U778 ( .A1(G2090), .A2(n693), .ZN(n694) );
  XNOR2_X1 U779 ( .A(KEYINPUT21), .B(n694), .ZN(n695) );
  NAND2_X1 U780 ( .A1(n695), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U781 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U782 ( .A1(G120), .A2(G57), .ZN(n696) );
  NOR2_X1 U783 ( .A1(G235), .A2(n696), .ZN(n697) );
  XNOR2_X1 U784 ( .A(KEYINPUT86), .B(n697), .ZN(n698) );
  NAND2_X1 U785 ( .A1(n698), .A2(G108), .ZN(n843) );
  NAND2_X1 U786 ( .A1(n843), .A2(G567), .ZN(n704) );
  XOR2_X1 U787 ( .A(KEYINPUT22), .B(KEYINPUT85), .Z(n700) );
  NAND2_X1 U788 ( .A1(G132), .A2(G82), .ZN(n699) );
  XNOR2_X1 U789 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X1 U790 ( .A1(n701), .A2(G218), .ZN(n702) );
  NAND2_X1 U791 ( .A1(G96), .A2(n702), .ZN(n842) );
  NAND2_X1 U792 ( .A1(n842), .A2(G2106), .ZN(n703) );
  NAND2_X1 U793 ( .A1(n704), .A2(n703), .ZN(n923) );
  NAND2_X1 U794 ( .A1(G661), .A2(G483), .ZN(n705) );
  NOR2_X1 U795 ( .A1(n923), .A2(n705), .ZN(n839) );
  NAND2_X1 U796 ( .A1(n839), .A2(G36), .ZN(G176) );
  NOR2_X1 U797 ( .A1(G1981), .A2(G305), .ZN(n706) );
  XNOR2_X1 U798 ( .A(n706), .B(KEYINPUT24), .ZN(n708) );
  NOR2_X1 U799 ( .A1(G164), .A2(G1384), .ZN(n793) );
  NAND2_X1 U800 ( .A1(G40), .A2(G160), .ZN(n707) );
  NAND2_X1 U801 ( .A1(n793), .A2(n791), .ZN(n746) );
  INV_X1 U802 ( .A(n780), .ZN(n770) );
  NAND2_X1 U803 ( .A1(n708), .A2(n770), .ZN(n784) );
  INV_X1 U804 ( .A(G1996), .ZN(n854) );
  NOR2_X1 U805 ( .A1(n746), .A2(n854), .ZN(n709) );
  XOR2_X1 U806 ( .A(n709), .B(KEYINPUT26), .Z(n711) );
  NAND2_X1 U807 ( .A1(n746), .A2(G1341), .ZN(n710) );
  NAND2_X1 U808 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U809 ( .A1(n992), .A2(n712), .ZN(n715) );
  OR2_X1 U810 ( .A1(n993), .A2(n715), .ZN(n719) );
  NAND2_X1 U811 ( .A1(n722), .A2(G2067), .ZN(n714) );
  NAND2_X1 U812 ( .A1(G1348), .A2(n746), .ZN(n713) );
  NAND2_X1 U813 ( .A1(n714), .A2(n713), .ZN(n717) );
  NAND2_X1 U814 ( .A1(n715), .A2(n993), .ZN(n716) );
  NAND2_X1 U815 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U816 ( .A1(n719), .A2(n718), .ZN(n727) );
  XOR2_X1 U817 ( .A(KEYINPUT93), .B(KEYINPUT27), .Z(n721) );
  NAND2_X1 U818 ( .A1(G2072), .A2(n722), .ZN(n720) );
  XNOR2_X1 U819 ( .A(n721), .B(n720), .ZN(n725) );
  NOR2_X1 U820 ( .A1(n725), .A2(n724), .ZN(n728) );
  NAND2_X1 U821 ( .A1(n984), .A2(n728), .ZN(n726) );
  NAND2_X1 U822 ( .A1(n727), .A2(n726), .ZN(n732) );
  XNOR2_X1 U823 ( .A(n730), .B(n729), .ZN(n731) );
  NAND2_X1 U824 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U825 ( .A1(n734), .A2(G1961), .ZN(n738) );
  XOR2_X1 U826 ( .A(G2078), .B(KEYINPUT25), .Z(n735) );
  XNOR2_X1 U827 ( .A(KEYINPUT92), .B(n735), .ZN(n955) );
  NOR2_X1 U828 ( .A1(n736), .A2(n955), .ZN(n737) );
  NOR2_X1 U829 ( .A1(n738), .A2(n737), .ZN(n743) );
  NOR2_X1 U830 ( .A1(G1966), .A2(n780), .ZN(n757) );
  NOR2_X1 U831 ( .A1(G2084), .A2(n746), .ZN(n754) );
  NOR2_X1 U832 ( .A1(n757), .A2(n754), .ZN(n739) );
  NAND2_X1 U833 ( .A1(G8), .A2(n739), .ZN(n740) );
  XNOR2_X1 U834 ( .A(KEYINPUT30), .B(n740), .ZN(n741) );
  NOR2_X1 U835 ( .A1(G168), .A2(n741), .ZN(n742) );
  XNOR2_X1 U836 ( .A(n742), .B(KEYINPUT95), .ZN(n745) );
  NAND2_X1 U837 ( .A1(n743), .A2(G301), .ZN(n744) );
  NAND2_X1 U838 ( .A1(n758), .A2(G286), .ZN(n751) );
  NOR2_X1 U839 ( .A1(G1971), .A2(n780), .ZN(n748) );
  NOR2_X1 U840 ( .A1(G2090), .A2(n746), .ZN(n747) );
  NOR2_X1 U841 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U842 ( .A1(n749), .A2(G303), .ZN(n750) );
  NAND2_X1 U843 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U844 ( .A1(n752), .A2(G8), .ZN(n753) );
  XNOR2_X1 U845 ( .A(n753), .B(KEYINPUT32), .ZN(n761) );
  NAND2_X1 U846 ( .A1(G8), .A2(n754), .ZN(n755) );
  XOR2_X1 U847 ( .A(KEYINPUT90), .B(n755), .Z(n756) );
  NOR2_X1 U848 ( .A1(n757), .A2(n756), .ZN(n759) );
  NAND2_X1 U849 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U850 ( .A1(n761), .A2(n760), .ZN(n762) );
  NOR2_X1 U851 ( .A1(G288), .A2(G1976), .ZN(n763) );
  XOR2_X1 U852 ( .A(n763), .B(KEYINPUT98), .Z(n989) );
  NOR2_X1 U853 ( .A1(G1971), .A2(G303), .ZN(n764) );
  XNOR2_X1 U854 ( .A(n764), .B(KEYINPUT99), .ZN(n765) );
  AND2_X1 U855 ( .A1(n989), .A2(n765), .ZN(n767) );
  INV_X1 U856 ( .A(KEYINPUT33), .ZN(n766) );
  AND2_X1 U857 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U858 ( .A1(G288), .A2(G1976), .ZN(n769) );
  XNOR2_X1 U859 ( .A(n769), .B(KEYINPUT100), .ZN(n982) );
  AND2_X1 U860 ( .A1(n770), .A2(n982), .ZN(n771) );
  OR2_X1 U861 ( .A1(KEYINPUT33), .A2(n771), .ZN(n773) );
  XNOR2_X1 U862 ( .A(G1981), .B(G305), .ZN(n980) );
  INV_X1 U863 ( .A(n980), .ZN(n772) );
  NOR2_X1 U864 ( .A1(n780), .A2(n989), .ZN(n774) );
  NAND2_X1 U865 ( .A1(KEYINPUT33), .A2(n774), .ZN(n775) );
  NAND2_X1 U866 ( .A1(n776), .A2(n775), .ZN(n786) );
  NOR2_X1 U867 ( .A1(G2090), .A2(G303), .ZN(n777) );
  NAND2_X1 U868 ( .A1(G8), .A2(n777), .ZN(n778) );
  NAND2_X1 U869 ( .A1(n779), .A2(n778), .ZN(n781) );
  NAND2_X1 U870 ( .A1(n781), .A2(n780), .ZN(n785) );
  AND2_X1 U871 ( .A1(n785), .A2(KEYINPUT101), .ZN(n782) );
  NAND2_X1 U872 ( .A1(n786), .A2(n782), .ZN(n783) );
  NAND2_X1 U873 ( .A1(n785), .A2(n786), .ZN(n788) );
  INV_X1 U874 ( .A(KEYINPUT101), .ZN(n787) );
  NAND2_X1 U875 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U876 ( .A(G1986), .B(G290), .ZN(n991) );
  INV_X1 U877 ( .A(n791), .ZN(n792) );
  NOR2_X1 U878 ( .A1(n793), .A2(n792), .ZN(n834) );
  NAND2_X1 U879 ( .A1(n991), .A2(n834), .ZN(n821) );
  XNOR2_X1 U880 ( .A(KEYINPUT37), .B(G2067), .ZN(n832) );
  NAND2_X1 U881 ( .A1(n904), .A2(G104), .ZN(n794) );
  XNOR2_X1 U882 ( .A(n794), .B(KEYINPUT88), .ZN(n796) );
  NAND2_X1 U883 ( .A1(G140), .A2(n905), .ZN(n795) );
  NAND2_X1 U884 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U885 ( .A(KEYINPUT34), .B(n797), .ZN(n802) );
  NAND2_X1 U886 ( .A1(G128), .A2(n900), .ZN(n799) );
  NAND2_X1 U887 ( .A1(G116), .A2(n901), .ZN(n798) );
  NAND2_X1 U888 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U889 ( .A(KEYINPUT35), .B(n800), .Z(n801) );
  NOR2_X1 U890 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U891 ( .A(KEYINPUT36), .B(n803), .ZN(n885) );
  NOR2_X1 U892 ( .A1(n832), .A2(n885), .ZN(n925) );
  NAND2_X1 U893 ( .A1(n925), .A2(n834), .ZN(n804) );
  XNOR2_X1 U894 ( .A(KEYINPUT89), .B(n804), .ZN(n829) );
  NAND2_X1 U895 ( .A1(G119), .A2(n900), .ZN(n806) );
  NAND2_X1 U896 ( .A1(G107), .A2(n901), .ZN(n805) );
  NAND2_X1 U897 ( .A1(n806), .A2(n805), .ZN(n810) );
  NAND2_X1 U898 ( .A1(G95), .A2(n904), .ZN(n808) );
  NAND2_X1 U899 ( .A1(G131), .A2(n905), .ZN(n807) );
  NAND2_X1 U900 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U901 ( .A1(n810), .A2(n809), .ZN(n897) );
  INV_X1 U902 ( .A(G1991), .ZN(n823) );
  NOR2_X1 U903 ( .A1(n897), .A2(n823), .ZN(n819) );
  NAND2_X1 U904 ( .A1(G129), .A2(n900), .ZN(n812) );
  NAND2_X1 U905 ( .A1(G117), .A2(n901), .ZN(n811) );
  NAND2_X1 U906 ( .A1(n812), .A2(n811), .ZN(n815) );
  NAND2_X1 U907 ( .A1(n904), .A2(G105), .ZN(n813) );
  XOR2_X1 U908 ( .A(KEYINPUT38), .B(n813), .Z(n814) );
  NOR2_X1 U909 ( .A1(n815), .A2(n814), .ZN(n817) );
  NAND2_X1 U910 ( .A1(n905), .A2(G141), .ZN(n816) );
  NAND2_X1 U911 ( .A1(n817), .A2(n816), .ZN(n911) );
  AND2_X1 U912 ( .A1(G1996), .A2(n911), .ZN(n818) );
  OR2_X1 U913 ( .A1(n819), .A2(n818), .ZN(n926) );
  AND2_X1 U914 ( .A1(n926), .A2(n834), .ZN(n826) );
  NOR2_X1 U915 ( .A1(n829), .A2(n826), .ZN(n820) );
  AND2_X1 U916 ( .A1(n821), .A2(n820), .ZN(n822) );
  NOR2_X1 U917 ( .A1(G1996), .A2(n911), .ZN(n928) );
  AND2_X1 U918 ( .A1(n823), .A2(n897), .ZN(n931) );
  NOR2_X1 U919 ( .A1(G1986), .A2(G290), .ZN(n824) );
  NOR2_X1 U920 ( .A1(n931), .A2(n824), .ZN(n825) );
  NOR2_X1 U921 ( .A1(n826), .A2(n825), .ZN(n827) );
  NOR2_X1 U922 ( .A1(n928), .A2(n827), .ZN(n828) );
  XNOR2_X1 U923 ( .A(n828), .B(KEYINPUT39), .ZN(n831) );
  INV_X1 U924 ( .A(n829), .ZN(n830) );
  NAND2_X1 U925 ( .A1(n831), .A2(n830), .ZN(n833) );
  NAND2_X1 U926 ( .A1(n832), .A2(n885), .ZN(n938) );
  NAND2_X1 U927 ( .A1(n833), .A2(n938), .ZN(n835) );
  NAND2_X1 U928 ( .A1(n835), .A2(n834), .ZN(n836) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n924), .ZN(G217) );
  NAND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n837) );
  XOR2_X1 U931 ( .A(KEYINPUT102), .B(n837), .Z(n838) );
  NAND2_X1 U932 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U933 ( .A1(G3), .A2(G1), .ZN(n840) );
  NAND2_X1 U934 ( .A1(n840), .A2(n839), .ZN(n841) );
  XOR2_X1 U935 ( .A(KEYINPUT103), .B(n841), .Z(G188) );
  XOR2_X1 U936 ( .A(G120), .B(KEYINPUT104), .Z(G236) );
  XNOR2_X1 U937 ( .A(G108), .B(KEYINPUT115), .ZN(G238) );
  INV_X1 U939 ( .A(G132), .ZN(G219) );
  INV_X1 U940 ( .A(G96), .ZN(G221) );
  INV_X1 U941 ( .A(G82), .ZN(G220) );
  INV_X1 U942 ( .A(G57), .ZN(G237) );
  NOR2_X1 U943 ( .A1(n843), .A2(n842), .ZN(n844) );
  XOR2_X1 U944 ( .A(n844), .B(KEYINPUT105), .Z(G325) );
  INV_X1 U945 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U946 ( .A(n992), .B(n845), .ZN(n848) );
  XOR2_X1 U947 ( .A(G301), .B(n846), .Z(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n849), .B(G286), .ZN(n850) );
  NOR2_X1 U950 ( .A1(G37), .A2(n850), .ZN(G397) );
  XOR2_X1 U951 ( .A(KEYINPUT41), .B(G1971), .Z(n852) );
  XNOR2_X1 U952 ( .A(G1961), .B(G1956), .ZN(n851) );
  XNOR2_X1 U953 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U954 ( .A(n853), .B(KEYINPUT109), .Z(n856) );
  XOR2_X1 U955 ( .A(n854), .B(G1991), .Z(n855) );
  XNOR2_X1 U956 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U957 ( .A(G1966), .B(G1976), .Z(n858) );
  XNOR2_X1 U958 ( .A(G1986), .B(G1981), .ZN(n857) );
  XNOR2_X1 U959 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U960 ( .A(n860), .B(n859), .Z(n862) );
  XNOR2_X1 U961 ( .A(KEYINPUT108), .B(G2474), .ZN(n861) );
  XNOR2_X1 U962 ( .A(n862), .B(n861), .ZN(G229) );
  XNOR2_X1 U963 ( .A(n863), .B(KEYINPUT43), .ZN(n865) );
  XNOR2_X1 U964 ( .A(KEYINPUT42), .B(G2678), .ZN(n864) );
  XNOR2_X1 U965 ( .A(n865), .B(n864), .ZN(n869) );
  XOR2_X1 U966 ( .A(KEYINPUT106), .B(G2090), .Z(n867) );
  XNOR2_X1 U967 ( .A(G2067), .B(G2072), .ZN(n866) );
  XNOR2_X1 U968 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U969 ( .A(n869), .B(n868), .Z(n871) );
  XNOR2_X1 U970 ( .A(KEYINPUT107), .B(G2096), .ZN(n870) );
  XNOR2_X1 U971 ( .A(n871), .B(n870), .ZN(n873) );
  XOR2_X1 U972 ( .A(G2078), .B(G2084), .Z(n872) );
  XNOR2_X1 U973 ( .A(n873), .B(n872), .ZN(G227) );
  NAND2_X1 U974 ( .A1(n905), .A2(G136), .ZN(n880) );
  NAND2_X1 U975 ( .A1(G100), .A2(n904), .ZN(n875) );
  NAND2_X1 U976 ( .A1(G112), .A2(n901), .ZN(n874) );
  NAND2_X1 U977 ( .A1(n875), .A2(n874), .ZN(n878) );
  NAND2_X1 U978 ( .A1(n900), .A2(G124), .ZN(n876) );
  XOR2_X1 U979 ( .A(KEYINPUT44), .B(n876), .Z(n877) );
  NOR2_X1 U980 ( .A1(n878), .A2(n877), .ZN(n879) );
  NAND2_X1 U981 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U982 ( .A(KEYINPUT110), .B(n881), .Z(G162) );
  XOR2_X1 U983 ( .A(KEYINPUT46), .B(KEYINPUT112), .Z(n883) );
  XNOR2_X1 U984 ( .A(KEYINPUT113), .B(KEYINPUT48), .ZN(n882) );
  XNOR2_X1 U985 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U986 ( .A(n885), .B(n884), .ZN(n887) );
  XNOR2_X1 U987 ( .A(G164), .B(G160), .ZN(n886) );
  XNOR2_X1 U988 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U989 ( .A(G162), .B(n888), .ZN(n899) );
  NAND2_X1 U990 ( .A1(G103), .A2(n904), .ZN(n890) );
  NAND2_X1 U991 ( .A1(G139), .A2(n905), .ZN(n889) );
  NAND2_X1 U992 ( .A1(n890), .A2(n889), .ZN(n896) );
  NAND2_X1 U993 ( .A1(G127), .A2(n900), .ZN(n892) );
  NAND2_X1 U994 ( .A1(G115), .A2(n901), .ZN(n891) );
  NAND2_X1 U995 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U996 ( .A(KEYINPUT111), .B(n893), .ZN(n894) );
  XNOR2_X1 U997 ( .A(KEYINPUT47), .B(n894), .ZN(n895) );
  NOR2_X1 U998 ( .A1(n896), .A2(n895), .ZN(n943) );
  XNOR2_X1 U999 ( .A(n897), .B(n943), .ZN(n898) );
  XNOR2_X1 U1000 ( .A(n899), .B(n898), .ZN(n915) );
  NAND2_X1 U1001 ( .A1(G130), .A2(n900), .ZN(n903) );
  NAND2_X1 U1002 ( .A1(G118), .A2(n901), .ZN(n902) );
  NAND2_X1 U1003 ( .A1(n903), .A2(n902), .ZN(n910) );
  NAND2_X1 U1004 ( .A1(G106), .A2(n904), .ZN(n907) );
  NAND2_X1 U1005 ( .A1(G142), .A2(n905), .ZN(n906) );
  NAND2_X1 U1006 ( .A1(n907), .A2(n906), .ZN(n908) );
  XOR2_X1 U1007 ( .A(n908), .B(KEYINPUT45), .Z(n909) );
  NOR2_X1 U1008 ( .A1(n910), .A2(n909), .ZN(n912) );
  XNOR2_X1 U1009 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1010 ( .A(n930), .B(n913), .Z(n914) );
  XNOR2_X1 U1011 ( .A(n915), .B(n914), .ZN(n916) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n916), .ZN(G395) );
  NOR2_X1 U1013 ( .A1(G401), .A2(n923), .ZN(n920) );
  NOR2_X1 U1014 ( .A1(G229), .A2(G227), .ZN(n917) );
  XNOR2_X1 U1015 ( .A(KEYINPUT49), .B(n917), .ZN(n918) );
  NOR2_X1 U1016 ( .A1(G397), .A2(n918), .ZN(n919) );
  NAND2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(n921) );
  NOR2_X1 U1018 ( .A1(n921), .A2(G395), .ZN(n922) );
  XOR2_X1 U1019 ( .A(n922), .B(KEYINPUT114), .Z(G225) );
  INV_X1 U1020 ( .A(G225), .ZN(G308) );
  INV_X1 U1021 ( .A(n923), .ZN(G319) );
  INV_X1 U1022 ( .A(n924), .ZN(G223) );
  XNOR2_X1 U1023 ( .A(KEYINPUT119), .B(KEYINPUT52), .ZN(n950) );
  OR2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n941) );
  XOR2_X1 U1025 ( .A(G2090), .B(G162), .Z(n927) );
  NOR2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1027 ( .A(KEYINPUT51), .B(n929), .ZN(n937) );
  NOR2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1029 ( .A(KEYINPUT116), .B(n932), .Z(n934) );
  XOR2_X1 U1030 ( .A(G160), .B(G2084), .Z(n933) );
  NOR2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1032 ( .A(KEYINPUT117), .B(n935), .ZN(n936) );
  NOR2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n939) );
  NAND2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1036 ( .A(KEYINPUT118), .B(n942), .ZN(n948) );
  XOR2_X1 U1037 ( .A(G2072), .B(n943), .Z(n945) );
  XOR2_X1 U1038 ( .A(G164), .B(G2078), .Z(n944) );
  NOR2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1040 ( .A(KEYINPUT50), .B(n946), .ZN(n947) );
  NAND2_X1 U1041 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1042 ( .A(n950), .B(n949), .ZN(n952) );
  INV_X1 U1043 ( .A(KEYINPUT55), .ZN(n951) );
  NAND2_X1 U1044 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1045 ( .A1(n953), .A2(G29), .ZN(n1033) );
  XOR2_X1 U1046 ( .A(G2084), .B(G34), .Z(n954) );
  XNOR2_X1 U1047 ( .A(KEYINPUT54), .B(n954), .ZN(n973) );
  XNOR2_X1 U1048 ( .A(G2090), .B(G35), .ZN(n971) );
  XOR2_X1 U1049 ( .A(G32), .B(G1996), .Z(n959) );
  XNOR2_X1 U1050 ( .A(n955), .B(G27), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(G26), .B(G2067), .ZN(n956) );
  NOR2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n961) );
  XNOR2_X1 U1054 ( .A(G33), .B(G2072), .ZN(n960) );
  NOR2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1056 ( .A(KEYINPUT122), .B(n962), .ZN(n967) );
  XNOR2_X1 U1057 ( .A(KEYINPUT120), .B(G25), .ZN(n963) );
  XOR2_X1 U1058 ( .A(n963), .B(G1991), .Z(n964) );
  NAND2_X1 U1059 ( .A1(G28), .A2(n964), .ZN(n965) );
  XNOR2_X1 U1060 ( .A(KEYINPUT121), .B(n965), .ZN(n966) );
  NAND2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1062 ( .A(n968), .B(KEYINPUT123), .ZN(n969) );
  XNOR2_X1 U1063 ( .A(n969), .B(KEYINPUT53), .ZN(n970) );
  NOR2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1066 ( .A(n974), .B(KEYINPUT124), .ZN(n975) );
  XOR2_X1 U1067 ( .A(n975), .B(KEYINPUT55), .Z(n977) );
  INV_X1 U1068 ( .A(G29), .ZN(n976) );
  NAND2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1070 ( .A1(G11), .A2(n978), .ZN(n1031) );
  INV_X1 U1071 ( .A(G16), .ZN(n1027) );
  XOR2_X1 U1072 ( .A(n1027), .B(KEYINPUT56), .Z(n1003) );
  XOR2_X1 U1073 ( .A(G1966), .B(G168), .Z(n979) );
  NOR2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1075 ( .A(KEYINPUT57), .B(n981), .Z(n1001) );
  XOR2_X1 U1076 ( .A(G303), .B(G1971), .Z(n983) );
  NAND2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n987) );
  XNOR2_X1 U1078 ( .A(G1956), .B(n984), .ZN(n985) );
  XNOR2_X1 U1079 ( .A(KEYINPUT125), .B(n985), .ZN(n986) );
  NOR2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n999) );
  XOR2_X1 U1082 ( .A(G1961), .B(G171), .Z(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n997) );
  XNOR2_X1 U1084 ( .A(n992), .B(G1341), .ZN(n995) );
  XOR2_X1 U1085 ( .A(n993), .B(G1348), .Z(n994) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n998) );
  NOR2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1090 ( .A1(n1003), .A2(n1002), .ZN(n1029) );
  XOR2_X1 U1091 ( .A(G1348), .B(KEYINPUT59), .Z(n1004) );
  XNOR2_X1 U1092 ( .A(G4), .B(n1004), .ZN(n1006) );
  XNOR2_X1 U1093 ( .A(G6), .B(G1981), .ZN(n1005) );
  NOR2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1010) );
  XNOR2_X1 U1095 ( .A(G1341), .B(G19), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(G1956), .B(G20), .ZN(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(n1011), .B(KEYINPUT60), .ZN(n1012) );
  XNOR2_X1 U1100 ( .A(KEYINPUT127), .B(n1012), .ZN(n1022) );
  XNOR2_X1 U1101 ( .A(G1961), .B(KEYINPUT126), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(n1013), .B(G5), .ZN(n1020) );
  XNOR2_X1 U1103 ( .A(G1976), .B(G23), .ZN(n1015) );
  XNOR2_X1 U1104 ( .A(G1971), .B(G22), .ZN(n1014) );
  NOR2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1017) );
  XOR2_X1 U1106 ( .A(G1986), .B(G24), .Z(n1016) );
  NAND2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1108 ( .A(KEYINPUT58), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1109 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1024) );
  XNOR2_X1 U1111 ( .A(G21), .B(G1966), .ZN(n1023) );
  NOR2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1113 ( .A(KEYINPUT61), .B(n1025), .ZN(n1026) );
  NAND2_X1 U1114 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1115 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NOR2_X1 U1116 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NAND2_X1 U1117 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XNOR2_X1 U1118 ( .A(KEYINPUT62), .B(n1034), .ZN(G150) );
  INV_X1 U1119 ( .A(G150), .ZN(G311) );
  INV_X1 U1120 ( .A(G303), .ZN(G166) );
endmodule

