//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 0 1 1 1 1 0 1 0 0 1 0 0 1 0 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n811, new_n812, new_n813,
    new_n814, new_n816, new_n817, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT67), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT67), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n204), .A2(G183gat), .A3(G190gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT24), .ZN(new_n206));
  AND3_X1   g005(.A1(new_n203), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  NAND3_X1  g006(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT68), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND4_X1  g009(.A1(KEYINPUT68), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n210), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n207), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216));
  OR2_X1    g015(.A1(new_n216), .A2(KEYINPUT66), .ZN(new_n217));
  NOR2_X1   g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT23), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n216), .A2(KEYINPUT66), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(G169gat), .B2(G176gat), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n217), .A2(new_n219), .A3(new_n220), .A4(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT25), .B1(new_n215), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n202), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT71), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT71), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n228), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n216), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT26), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n231), .B1(new_n232), .B2(new_n218), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n225), .B1(new_n230), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(G183gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT27), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT27), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(G183gat), .ZN(new_n238));
  INV_X1    g037(.A(G190gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n236), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT69), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AND2_X1   g041(.A1(KEYINPUT70), .A2(KEYINPUT28), .ZN(new_n243));
  NOR2_X1   g042(.A1(KEYINPUT70), .A2(KEYINPUT28), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n242), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n240), .A2(new_n241), .A3(new_n245), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n234), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT25), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n222), .A2(new_n250), .A3(new_n216), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n202), .B1(new_n212), .B2(new_n206), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n251), .B1(new_n208), .B2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT64), .B(G169gat), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n221), .A2(G176gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT65), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT65), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n254), .A2(new_n258), .A3(new_n255), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n253), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n224), .A2(new_n249), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT73), .ZN(new_n262));
  INV_X1    g061(.A(G226gat), .ZN(new_n263));
  INV_X1    g062(.A(G233gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT73), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n224), .A2(new_n249), .A3(new_n266), .A4(new_n260), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n262), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n265), .A2(KEYINPUT29), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n261), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  AND2_X1   g070(.A1(G211gat), .A2(G218gat), .ZN(new_n272));
  NOR2_X1   g071(.A1(G211gat), .A2(G218gat), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT72), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G211gat), .ZN(new_n275));
  INV_X1    g074(.A(G218gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT72), .ZN(new_n278));
  NAND2_X1  g077(.A1(G211gat), .A2(G218gat), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n274), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(G197gat), .ZN(new_n282));
  INV_X1    g081(.A(G204gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(G197gat), .A2(G204gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT22), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n279), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n281), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n274), .A2(new_n280), .A3(new_n288), .A4(new_n286), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n271), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n262), .A2(new_n267), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(new_n269), .ZN(new_n295));
  INV_X1    g094(.A(new_n292), .ZN(new_n296));
  INV_X1    g095(.A(new_n265), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n261), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n295), .A2(new_n296), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n293), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G8gat), .B(G36gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(G64gat), .B(G92gat), .ZN(new_n303));
  XOR2_X1   g102(.A(new_n302), .B(new_n303), .Z(new_n304));
  NAND2_X1  g103(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n304), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n293), .A2(new_n300), .A3(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n305), .A2(KEYINPUT30), .A3(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT30), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n301), .A2(new_n309), .A3(new_n304), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  AND2_X1   g110(.A1(G155gat), .A2(G162gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(G155gat), .A2(G162gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G141gat), .B(G148gat), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n314), .B1(new_n315), .B2(KEYINPUT2), .ZN(new_n316));
  INV_X1    g115(.A(G141gat), .ZN(new_n317));
  AND2_X1   g116(.A1(new_n317), .A2(G148gat), .ZN(new_n318));
  AND2_X1   g117(.A1(KEYINPUT74), .A2(G148gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(KEYINPUT74), .A2(G148gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n318), .B1(new_n321), .B2(G141gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT2), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n312), .B1(new_n323), .B2(new_n313), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n316), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT75), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  XOR2_X1   g126(.A(G127gat), .B(G134gat), .Z(new_n328));
  XNOR2_X1  g127(.A(G113gat), .B(G120gat), .ZN(new_n329));
  OR3_X1    g128(.A1(new_n328), .A2(KEYINPUT1), .A3(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n328), .B1(KEYINPUT1), .B2(new_n329), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NOR3_X1   g131(.A1(new_n319), .A2(new_n320), .A3(new_n317), .ZN(new_n333));
  NOR3_X1   g132(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n334));
  OAI22_X1  g133(.A1(new_n333), .A2(new_n318), .B1(new_n312), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n335), .A2(KEYINPUT75), .A3(new_n316), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n327), .A2(new_n332), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n325), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n329), .A2(KEYINPUT1), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(new_n328), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(G225gat), .A2(G233gat), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n345), .A2(KEYINPUT77), .A3(KEYINPUT5), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT77), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n343), .B1(new_n337), .B2(new_n341), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT5), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT3), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n351), .B(new_n316), .C1(new_n322), .C2(new_n324), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT76), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n335), .A2(KEYINPUT76), .A3(new_n351), .A4(new_n316), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n327), .A2(new_n336), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n356), .B(new_n332), .C1(new_n357), .C2(new_n351), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT4), .B1(new_n338), .B2(new_n340), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT4), .ZN(new_n360));
  NOR3_X1   g159(.A1(new_n332), .A2(new_n325), .A3(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n358), .A2(new_n362), .A3(new_n343), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n346), .A2(new_n350), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT78), .ZN(new_n365));
  XNOR2_X1  g164(.A(G1gat), .B(G29gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n366), .B(KEYINPUT0), .ZN(new_n367));
  XNOR2_X1  g166(.A(G57gat), .B(G85gat), .ZN(new_n368));
  XOR2_X1   g167(.A(new_n367), .B(new_n368), .Z(new_n369));
  OR2_X1    g168(.A1(new_n363), .A2(KEYINPUT5), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT78), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n346), .A2(new_n350), .A3(new_n363), .A4(new_n371), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n365), .A2(new_n369), .A3(new_n370), .A4(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT6), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AND2_X1   g174(.A1(new_n372), .A2(new_n370), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n369), .B1(new_n376), .B2(new_n365), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n365), .A2(new_n370), .A3(new_n372), .ZN(new_n379));
  INV_X1    g178(.A(new_n369), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n379), .A2(KEYINPUT6), .A3(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n311), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(G228gat), .A2(G233gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n383), .B(KEYINPUT80), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT29), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n290), .A2(new_n386), .A3(new_n291), .ZN(new_n387));
  AND2_X1   g186(.A1(new_n387), .A2(new_n351), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n388), .A2(new_n338), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n356), .A2(new_n386), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n292), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n389), .B1(new_n391), .B2(KEYINPUT81), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT81), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n390), .A2(new_n393), .A3(new_n292), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n385), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n296), .B1(new_n356), .B2(new_n386), .ZN(new_n396));
  INV_X1    g195(.A(new_n383), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n397), .B1(new_n388), .B2(new_n357), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(G22gat), .B1(new_n395), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n389), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT29), .B1(new_n354), .B2(new_n355), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT81), .B1(new_n402), .B2(new_n296), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n394), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n384), .ZN(new_n405));
  INV_X1    g204(.A(G22gat), .ZN(new_n406));
  INV_X1    g205(.A(new_n399), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(G78gat), .B(G106gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(KEYINPUT31), .B(G50gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n400), .A2(new_n408), .A3(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(KEYINPUT79), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n406), .B1(new_n405), .B2(new_n407), .ZN(new_n414));
  AOI211_X1 g213(.A(G22gat), .B(new_n399), .C1(new_n404), .C2(new_n384), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n412), .A2(new_n416), .A3(KEYINPUT82), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT82), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n418), .B(new_n413), .C1(new_n414), .C2(new_n415), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n382), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n261), .A2(new_n332), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n340), .A2(new_n224), .A3(new_n249), .A4(new_n260), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(G227gat), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n425), .A2(new_n264), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT33), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(G15gat), .B(G43gat), .ZN(new_n428));
  XNOR2_X1  g227(.A(G71gat), .B(G99gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n428), .B(new_n429), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT34), .B1(new_n424), .B2(new_n426), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT34), .ZN(new_n433));
  INV_X1    g232(.A(new_n426), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n422), .A2(new_n433), .A3(new_n434), .A4(new_n423), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n431), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT32), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n438), .B1(new_n424), .B2(new_n426), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n432), .B(new_n435), .C1(new_n427), .C2(new_n430), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n437), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n439), .B1(new_n437), .B2(new_n440), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n443), .B(KEYINPUT36), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n271), .A2(new_n292), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT37), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n269), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n448), .B1(new_n262), .B2(new_n267), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n292), .B1(new_n449), .B2(new_n298), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT38), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n304), .A2(new_n446), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n307), .A2(new_n453), .ZN(new_n454));
  AOI22_X1  g253(.A1(new_n451), .A2(new_n454), .B1(new_n301), .B2(new_n304), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT38), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n293), .A2(new_n300), .A3(KEYINPUT37), .ZN(new_n457));
  AOI211_X1 g256(.A(KEYINPUT85), .B(new_n456), .C1(new_n454), .C2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT85), .ZN(new_n459));
  NOR3_X1   g258(.A1(new_n449), .A2(new_n292), .A3(new_n298), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n296), .B1(new_n268), .B2(new_n270), .ZN(new_n461));
  NOR3_X1   g260(.A1(new_n460), .A2(new_n461), .A3(new_n304), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n457), .B1(new_n462), .B2(new_n452), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n459), .B1(new_n463), .B2(KEYINPUT38), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n455), .B1(new_n458), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n379), .A2(new_n380), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n466), .A2(new_n374), .A3(new_n373), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n375), .A2(new_n377), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n358), .A2(new_n362), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n344), .B1(new_n471), .B2(KEYINPUT39), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n342), .A2(KEYINPUT39), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n344), .B1(KEYINPUT83), .B2(KEYINPUT39), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n474), .B1(KEYINPUT83), .B2(KEYINPUT39), .ZN(new_n475));
  AOI22_X1  g274(.A1(new_n472), .A2(new_n473), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(KEYINPUT84), .B1(new_n476), .B2(new_n380), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT40), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT40), .ZN(new_n479));
  OAI211_X1 g278(.A(KEYINPUT84), .B(new_n479), .C1(new_n476), .C2(new_n380), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n310), .A3(new_n308), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n417), .B(new_n419), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n421), .B(new_n444), .C1(new_n470), .C2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n417), .A2(new_n419), .A3(new_n443), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT86), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT86), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n417), .A2(new_n487), .A3(new_n443), .A4(new_n419), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT35), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n382), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n490), .B1(new_n382), .B2(new_n485), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n484), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(G29gat), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n495), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n496));
  XOR2_X1   g295(.A(KEYINPUT14), .B(G29gat), .Z(new_n497));
  OAI21_X1  g296(.A(new_n496), .B1(new_n497), .B2(G36gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(G43gat), .B(G50gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT15), .ZN(new_n500));
  OR2_X1    g299(.A1(new_n499), .A2(KEYINPUT15), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n498), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT87), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n498), .A2(new_n501), .A3(KEYINPUT87), .A4(new_n500), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n504), .B(new_n505), .C1(new_n498), .C2(new_n500), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT17), .ZN(new_n507));
  OR2_X1    g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(G15gat), .B(G22gat), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT16), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n509), .B1(new_n510), .B2(G1gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(KEYINPUT88), .A2(G8gat), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n511), .B(new_n512), .C1(G1gat), .C2(new_n509), .ZN(new_n513));
  NOR2_X1   g312(.A1(KEYINPUT88), .A2(G8gat), .ZN(new_n514));
  XOR2_X1   g313(.A(new_n513), .B(new_n514), .Z(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n506), .A2(new_n507), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n508), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(G229gat), .A2(G233gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n515), .A2(new_n506), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT89), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT18), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n515), .B(new_n506), .ZN(new_n525));
  XOR2_X1   g324(.A(new_n519), .B(KEYINPUT13), .Z(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n522), .A2(new_n523), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n518), .A2(new_n519), .A3(new_n520), .A4(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n524), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G113gat), .B(G141gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(G197gat), .ZN(new_n532));
  XOR2_X1   g331(.A(KEYINPUT11), .B(G169gat), .Z(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  XOR2_X1   g333(.A(new_n534), .B(KEYINPUT12), .Z(new_n535));
  NAND2_X1  g334(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n535), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n524), .A2(new_n537), .A3(new_n527), .A4(new_n529), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n494), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(G64gat), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n541), .A2(G57gat), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(G57gat), .ZN(new_n543));
  AND2_X1   g342(.A1(G71gat), .A2(G78gat), .ZN(new_n544));
  OAI22_X1  g343(.A1(new_n542), .A2(new_n543), .B1(KEYINPUT9), .B2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G71gat), .B(G78gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT21), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(G231gat), .A2(G233gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(G127gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n516), .B1(new_n549), .B2(new_n548), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G183gat), .B(G211gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT90), .ZN(new_n558));
  XNOR2_X1  g357(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n559));
  INV_X1    g358(.A(G155gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n558), .B(new_n561), .ZN(new_n562));
  OR2_X1    g361(.A1(new_n556), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n556), .A2(new_n562), .ZN(new_n564));
  AND2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(KEYINPUT91), .B(KEYINPUT7), .ZN(new_n566));
  NAND2_X1  g365(.A1(G85gat), .A2(G92gat), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n567), .ZN(new_n569));
  NAND2_X1  g368(.A1(G99gat), .A2(G106gat), .ZN(new_n570));
  INV_X1    g369(.A(G85gat), .ZN(new_n571));
  INV_X1    g370(.A(G92gat), .ZN(new_n572));
  AOI22_X1  g371(.A1(KEYINPUT8), .A2(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n568), .A2(new_n569), .A3(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G99gat), .B(G106gat), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n568), .A2(new_n575), .A3(new_n569), .A4(new_n573), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n508), .A2(new_n517), .A3(new_n579), .ZN(new_n580));
  AND3_X1   g379(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n581));
  AND2_X1   g380(.A1(new_n577), .A2(new_n578), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n581), .B1(new_n506), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT92), .ZN(new_n584));
  AND2_X1   g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n583), .A2(new_n584), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n580), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G190gat), .B(G218gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT93), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT94), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n589), .B(new_n580), .C1(new_n585), .C2(new_n586), .ZN(new_n594));
  XNOR2_X1  g393(.A(G134gat), .B(G162gat), .ZN(new_n595));
  AOI21_X1  g394(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n595), .B(new_n596), .Z(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n587), .A2(KEYINPUT94), .A3(new_n590), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n593), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT95), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n593), .A2(new_n599), .A3(KEYINPUT95), .A4(new_n600), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n591), .A2(new_n594), .ZN(new_n605));
  AOI22_X1  g404(.A1(new_n603), .A2(new_n604), .B1(new_n605), .B2(new_n597), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n565), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(G230gat), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n608), .A2(new_n264), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT96), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n578), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n579), .A2(new_n547), .A3(new_n612), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n578), .B(new_n577), .C1(new_n548), .C2(new_n611), .ZN(new_n614));
  AOI21_X1  g413(.A(KEYINPUT10), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AND3_X1   g414(.A1(new_n582), .A2(KEYINPUT10), .A3(new_n547), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n610), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n613), .A2(new_n614), .A3(new_n609), .ZN(new_n618));
  XNOR2_X1  g417(.A(G120gat), .B(G148gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(G176gat), .B(G204gat), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n619), .B(new_n620), .Z(new_n621));
  NAND3_X1  g420(.A1(new_n617), .A2(new_n618), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT97), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n617), .A2(new_n618), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n621), .B(KEYINPUT98), .Z(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  OR3_X1    g426(.A1(new_n607), .A2(KEYINPUT99), .A3(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(KEYINPUT99), .B1(new_n607), .B2(new_n627), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n540), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n469), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g432(.A(KEYINPUT100), .B(G1gat), .Z(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(G1324gat));
  INV_X1    g434(.A(new_n311), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n631), .A2(new_n636), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n637), .A2(G8gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(KEYINPUT16), .B(G8gat), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(KEYINPUT42), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n641), .B1(KEYINPUT42), .B2(new_n640), .ZN(G1325gat));
  INV_X1    g441(.A(new_n631), .ZN(new_n643));
  OAI21_X1  g442(.A(G15gat), .B1(new_n643), .B2(new_n444), .ZN(new_n644));
  INV_X1    g443(.A(new_n443), .ZN(new_n645));
  OR2_X1    g444(.A1(new_n645), .A2(G15gat), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n644), .B1(new_n643), .B2(new_n646), .ZN(G1326gat));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n420), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT101), .ZN(new_n649));
  XNOR2_X1  g448(.A(KEYINPUT43), .B(G22gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(G1327gat));
  INV_X1    g450(.A(new_n565), .ZN(new_n652));
  INV_X1    g451(.A(new_n627), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n603), .A2(new_n604), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n605), .A2(new_n597), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT102), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(new_n540), .ZN(new_n661));
  NOR3_X1   g460(.A1(new_n661), .A2(G29gat), .A3(new_n469), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n662), .B(KEYINPUT45), .Z(new_n663));
  NAND2_X1  g462(.A1(new_n494), .A2(KEYINPUT103), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT103), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n484), .A2(new_n492), .A3(new_n665), .A4(new_n493), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n606), .A2(KEYINPUT44), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n664), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n494), .A2(new_n658), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(KEYINPUT44), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n671), .A2(new_n539), .A3(new_n655), .ZN(new_n672));
  OAI21_X1  g471(.A(G29gat), .B1(new_n672), .B2(new_n469), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n663), .A2(new_n673), .ZN(G1328gat));
  NOR3_X1   g473(.A1(new_n661), .A2(G36gat), .A3(new_n311), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(KEYINPUT46), .ZN(new_n676));
  OAI21_X1  g475(.A(G36gat), .B1(new_n672), .B2(new_n311), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(G1329gat));
  NOR3_X1   g477(.A1(new_n661), .A2(G43gat), .A3(new_n645), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n672), .A2(new_n444), .ZN(new_n681));
  OAI21_X1  g480(.A(G43gat), .B1(new_n681), .B2(KEYINPUT104), .ZN(new_n682));
  INV_X1    g481(.A(new_n539), .ZN(new_n683));
  AOI211_X1 g482(.A(new_n683), .B(new_n654), .C1(new_n668), .C2(new_n670), .ZN(new_n684));
  INV_X1    g483(.A(new_n444), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n684), .A2(KEYINPUT104), .A3(new_n685), .ZN(new_n686));
  OAI211_X1 g485(.A(KEYINPUT47), .B(new_n680), .C1(new_n682), .C2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(G43gat), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n680), .B1(new_n681), .B2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT47), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n687), .A2(new_n691), .ZN(G1330gat));
  INV_X1    g491(.A(G50gat), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n420), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g493(.A(new_n694), .B(KEYINPUT105), .Z(new_n695));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n696));
  OAI22_X1  g495(.A1(new_n661), .A2(new_n695), .B1(new_n696), .B2(KEYINPUT48), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n684), .A2(new_n420), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n697), .B1(new_n698), .B2(G50gat), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n696), .A2(KEYINPUT48), .ZN(new_n700));
  XOR2_X1   g499(.A(new_n700), .B(KEYINPUT107), .Z(new_n701));
  XNOR2_X1  g500(.A(new_n699), .B(new_n701), .ZN(G1331gat));
  AND2_X1   g501(.A1(new_n664), .A2(new_n666), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n607), .A2(new_n539), .A3(new_n653), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(new_n632), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g507(.A(new_n311), .B(KEYINPUT108), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT49), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n709), .B1(new_n710), .B2(new_n541), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT109), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n706), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n710), .A2(new_n541), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(G1333gat));
  OAI21_X1  g514(.A(G71gat), .B1(new_n705), .B2(new_n444), .ZN(new_n716));
  OR2_X1    g515(.A1(new_n645), .A2(G71gat), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n716), .B1(new_n705), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1334gat));
  NAND2_X1  g519(.A1(new_n706), .A2(new_n420), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g521(.A1(new_n652), .A2(new_n683), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n723), .A2(new_n653), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n725), .B1(new_n668), .B2(new_n670), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(G85gat), .B1(new_n727), .B2(new_n469), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT112), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT51), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n723), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n494), .A2(KEYINPUT111), .A3(new_n658), .ZN(new_n732));
  AOI21_X1  g531(.A(KEYINPUT111), .B1(new_n494), .B2(new_n658), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n731), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n729), .A2(new_n730), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OAI221_X1 g535(.A(new_n731), .B1(new_n729), .B2(new_n730), .C1(new_n732), .C2(new_n733), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n632), .A2(new_n571), .A3(new_n627), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT113), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n736), .A2(new_n737), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n728), .A2(new_n740), .ZN(G1336gat));
  INV_X1    g540(.A(new_n709), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n742), .A2(G92gat), .A3(new_n653), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n736), .A2(new_n737), .A3(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n671), .A2(new_n709), .A3(new_n724), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G92gat), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT52), .ZN(new_n747));
  AND3_X1   g546(.A1(new_n744), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n671), .A2(new_n636), .A3(new_n724), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G92gat), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n747), .B1(new_n744), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(KEYINPUT114), .B1(new_n748), .B2(new_n751), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n736), .A2(new_n737), .A3(new_n743), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n572), .B1(new_n726), .B2(new_n636), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT52), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT114), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n744), .A2(new_n746), .A3(new_n747), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n755), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n752), .A2(new_n758), .ZN(G1337gat));
  OAI21_X1  g558(.A(G99gat), .B1(new_n727), .B2(new_n444), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n653), .A2(new_n645), .A3(G99gat), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n736), .A2(new_n737), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n762), .ZN(G1338gat));
  NAND2_X1  g562(.A1(new_n726), .A2(new_n420), .ZN(new_n764));
  AOI22_X1  g563(.A1(new_n764), .A2(G106gat), .B1(KEYINPUT115), .B2(KEYINPUT53), .ZN(new_n765));
  INV_X1    g564(.A(new_n420), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n766), .A2(G106gat), .A3(new_n653), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n736), .A2(new_n737), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  OR2_X1    g568(.A1(KEYINPUT115), .A2(KEYINPUT53), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n769), .B(new_n770), .ZN(G1339gat));
  NAND4_X1  g570(.A1(new_n565), .A2(new_n606), .A3(new_n683), .A4(new_n653), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT116), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n519), .B1(new_n518), .B2(new_n520), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n525), .A2(new_n526), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n534), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n538), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n627), .ZN(new_n779));
  OR3_X1    g578(.A1(new_n615), .A2(new_n610), .A3(new_n616), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n780), .A2(KEYINPUT54), .A3(new_n617), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT54), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n782), .B(new_n610), .C1(new_n615), .C2(new_n616), .ZN(new_n783));
  INV_X1    g582(.A(new_n621), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n783), .A2(KEYINPUT117), .A3(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT117), .B1(new_n783), .B2(new_n784), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n781), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n781), .B(KEYINPUT55), .C1(new_n786), .C2(new_n787), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n790), .A2(new_n623), .A3(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n539), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n658), .B1(new_n779), .B2(new_n794), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n606), .A2(new_n777), .A3(new_n792), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n652), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n773), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n798), .A2(new_n469), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n489), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n800), .A2(new_n709), .ZN(new_n801));
  INV_X1    g600(.A(G113gat), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n801), .A2(new_n802), .A3(new_n539), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n798), .A2(new_n420), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n709), .A2(new_n469), .A3(new_n645), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n804), .A2(new_n539), .A3(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n806), .A2(KEYINPUT118), .A3(G113gat), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(KEYINPUT118), .B1(new_n806), .B2(G113gat), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n803), .B1(new_n808), .B2(new_n809), .ZN(G1340gat));
  NAND2_X1  g609(.A1(new_n804), .A2(new_n805), .ZN(new_n811));
  INV_X1    g610(.A(G120gat), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n811), .A2(new_n812), .A3(new_n653), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n801), .A2(new_n627), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n813), .B1(new_n814), .B2(new_n812), .ZN(G1341gat));
  NAND3_X1  g614(.A1(new_n801), .A2(new_n553), .A3(new_n565), .ZN(new_n816));
  OAI21_X1  g615(.A(G127gat), .B1(new_n811), .B2(new_n652), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(G1342gat));
  NOR4_X1   g617(.A1(new_n800), .A2(G134gat), .A3(new_n636), .A4(new_n606), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT56), .ZN(new_n820));
  OR2_X1    g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n820), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n804), .A2(new_n658), .A3(new_n805), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT119), .B1(new_n823), .B2(G134gat), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n823), .A2(KEYINPUT119), .A3(G134gat), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n821), .B(new_n822), .C1(new_n824), .C2(new_n826), .ZN(G1343gat));
  NOR3_X1   g626(.A1(new_n685), .A2(new_n709), .A3(new_n469), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT57), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n830), .B1(new_n798), .B2(new_n766), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT120), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n791), .A2(new_n623), .ZN(new_n833));
  INV_X1    g632(.A(new_n787), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n785), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT55), .B1(new_n835), .B2(new_n781), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n832), .B1(new_n833), .B2(new_n836), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n790), .A2(KEYINPUT120), .A3(new_n623), .A4(new_n791), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n837), .A2(new_n539), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n658), .B1(new_n839), .B2(new_n779), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n652), .B1(new_n840), .B2(new_n796), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n773), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n766), .A2(new_n830), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n829), .B1(new_n831), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n317), .B1(new_n845), .B2(new_n539), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n685), .A2(new_n766), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n799), .A2(new_n847), .ZN(new_n848));
  NOR4_X1   g647(.A1(new_n848), .A2(G141gat), .A3(new_n683), .A4(new_n709), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT58), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(KEYINPUT58), .B1(new_n846), .B2(new_n849), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(G1344gat));
  NOR2_X1   g653(.A1(new_n848), .A2(new_n709), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n321), .A3(new_n627), .ZN(new_n856));
  AOI211_X1 g655(.A(KEYINPUT59), .B(new_n321), .C1(new_n845), .C2(new_n627), .ZN(new_n857));
  XNOR2_X1  g656(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n858));
  INV_X1    g657(.A(new_n796), .ZN(new_n859));
  INV_X1    g658(.A(new_n779), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n683), .B1(new_n792), .B2(new_n832), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n860), .B1(new_n861), .B2(new_n838), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n859), .B(KEYINPUT122), .C1(new_n862), .C2(new_n658), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT122), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n864), .B1(new_n840), .B2(new_n796), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n863), .A2(new_n865), .A3(new_n652), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n628), .A2(new_n683), .A3(new_n629), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(KEYINPUT57), .B1(new_n868), .B2(new_n420), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n773), .A2(new_n797), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n843), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n627), .B(new_n828), .C1(new_n869), .C2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n858), .B1(new_n873), .B2(G148gat), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n856), .B1(new_n857), .B2(new_n874), .ZN(G1345gat));
  INV_X1    g674(.A(new_n845), .ZN(new_n876));
  OAI21_X1  g675(.A(G155gat), .B1(new_n876), .B2(new_n652), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n855), .A2(new_n560), .A3(new_n565), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(G1346gat));
  OAI21_X1  g678(.A(G162gat), .B1(new_n876), .B2(new_n606), .ZN(new_n880));
  INV_X1    g679(.A(G162gat), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n658), .A2(new_n881), .A3(new_n311), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n880), .B1(new_n848), .B2(new_n882), .ZN(G1347gat));
  NOR2_X1   g682(.A1(new_n632), .A2(new_n311), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(new_n645), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n804), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(G169gat), .B1(new_n887), .B2(new_n683), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n798), .A2(new_n632), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n742), .B1(new_n486), .B2(new_n488), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n539), .A2(new_n254), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n888), .B1(new_n891), .B2(new_n892), .ZN(G1348gat));
  INV_X1    g692(.A(G176gat), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n887), .A2(new_n894), .A3(new_n653), .ZN(new_n895));
  INV_X1    g694(.A(new_n891), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n627), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n895), .B1(new_n894), .B2(new_n897), .ZN(G1349gat));
  NAND4_X1  g697(.A1(new_n896), .A2(new_n236), .A3(new_n238), .A4(new_n565), .ZN(new_n899));
  OAI21_X1  g698(.A(G183gat), .B1(new_n887), .B2(new_n652), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n899), .A2(KEYINPUT123), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(KEYINPUT60), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT60), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n899), .A2(new_n900), .A3(KEYINPUT123), .A4(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(G1350gat));
  NAND3_X1  g704(.A1(new_n896), .A2(new_n239), .A3(new_n658), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n804), .A2(new_n658), .A3(new_n886), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT61), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n907), .A2(new_n908), .A3(G190gat), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n908), .B1(new_n907), .B2(G190gat), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n906), .B1(new_n910), .B2(new_n911), .ZN(G1351gat));
  NAND4_X1  g711(.A1(new_n870), .A2(new_n469), .A3(new_n709), .A4(new_n847), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(G197gat), .B1(new_n914), .B2(new_n539), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n869), .A2(new_n872), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n885), .A2(new_n685), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n683), .A2(new_n282), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n915), .B1(new_n919), .B2(new_n920), .ZN(G1352gat));
  OAI211_X1 g720(.A(new_n627), .B(new_n917), .C1(new_n869), .C2(new_n872), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(G204gat), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n870), .A2(new_n469), .A3(new_n847), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n709), .A2(new_n283), .A3(new_n627), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n926), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n927));
  XNOR2_X1  g726(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n923), .A2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT125), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n923), .A2(new_n929), .A3(KEYINPUT125), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1353gat));
  NAND3_X1  g733(.A1(new_n914), .A2(new_n275), .A3(new_n565), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n565), .B(new_n917), .C1(new_n869), .C2(new_n872), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n936), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n937));
  AOI21_X1  g736(.A(KEYINPUT63), .B1(new_n936), .B2(G211gat), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n935), .B1(new_n937), .B2(new_n938), .ZN(G1354gat));
  OAI21_X1  g738(.A(new_n276), .B1(new_n913), .B2(new_n606), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT126), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n658), .A2(G218gat), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT127), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n942), .B1(new_n919), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g743(.A(KEYINPUT127), .B1(new_n916), .B2(new_n918), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n941), .B1(new_n944), .B2(new_n945), .ZN(G1355gat));
endmodule


