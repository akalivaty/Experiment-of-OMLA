//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 0 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 1 1 1 0 1 1 0 0 1 1 1 0 1 0 1 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n736, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  AND2_X1   g003(.A1(KEYINPUT72), .A2(G953), .ZN(new_n190));
  NOR2_X1   g004(.A1(KEYINPUT72), .A2(G953), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(G221), .A3(G234), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT22), .B(G137), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n193), .B(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT77), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(new_n193), .B(new_n194), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT77), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT76), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT16), .ZN(new_n204));
  AND2_X1   g018(.A1(KEYINPUT75), .A2(G125), .ZN(new_n205));
  NOR2_X1   g019(.A1(KEYINPUT75), .A2(G125), .ZN(new_n206));
  OAI21_X1  g020(.A(G140), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(G125), .A2(G140), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n204), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n205), .A2(new_n206), .ZN(new_n211));
  NOR3_X1   g025(.A1(new_n211), .A2(KEYINPUT16), .A3(G140), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n203), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT75), .B(G125), .ZN(new_n214));
  INV_X1    g028(.A(G140), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(new_n204), .A3(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n208), .B1(new_n214), .B2(G140), .ZN(new_n217));
  OAI211_X1 g031(.A(G146), .B(new_n216), .C1(new_n217), .C2(new_n204), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n213), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT69), .B(G128), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G119), .ZN(new_n221));
  INV_X1    g035(.A(G119), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G128), .ZN(new_n223));
  XOR2_X1   g037(.A(KEYINPUT24), .B(G110), .Z(new_n224));
  NAND3_X1  g038(.A1(new_n221), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT23), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n226), .B1(new_n222), .B2(G128), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(new_n223), .ZN(new_n228));
  INV_X1    g042(.A(G128), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT69), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G128), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n230), .A2(new_n232), .A3(KEYINPUT23), .A4(G119), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT74), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n220), .A2(KEYINPUT74), .A3(KEYINPUT23), .A4(G119), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n228), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G110), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n225), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n202), .B1(new_n219), .B2(new_n239), .ZN(new_n240));
  OR2_X1    g054(.A1(new_n237), .A2(new_n238), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n213), .A2(new_n218), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n241), .A2(KEYINPUT76), .A3(new_n242), .A4(new_n225), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n224), .B1(new_n221), .B2(new_n223), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n245), .B1(new_n237), .B2(new_n238), .ZN(new_n246));
  XNOR2_X1  g060(.A(G125), .B(G140), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(new_n203), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n218), .A2(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n201), .B1(new_n244), .B2(new_n251), .ZN(new_n252));
  AOI211_X1 g066(.A(new_n250), .B(new_n196), .C1(new_n240), .C2(new_n243), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(KEYINPUT25), .B1(new_n254), .B2(new_n188), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT25), .ZN(new_n256));
  NOR4_X1   g070(.A1(new_n252), .A2(new_n253), .A3(new_n256), .A4(G902), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n189), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n254), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n189), .A2(G902), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n258), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G237), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n192), .A2(G210), .A3(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n264), .B(KEYINPUT27), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT26), .B(G101), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n265), .B(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT28), .ZN(new_n269));
  XOR2_X1   g083(.A(KEYINPUT2), .B(G113), .Z(new_n270));
  XNOR2_X1  g084(.A(G116), .B(G119), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT71), .ZN(new_n273));
  INV_X1    g087(.A(new_n271), .ZN(new_n274));
  XNOR2_X1  g088(.A(KEYINPUT2), .B(G113), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n273), .B(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(G134), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT66), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT66), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G134), .ZN(new_n281));
  AOI21_X1  g095(.A(G137), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G137), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(G134), .ZN(new_n284));
  OAI21_X1  g098(.A(G131), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n279), .A2(new_n281), .A3(G137), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n283), .A2(KEYINPUT11), .A3(G134), .ZN(new_n287));
  XNOR2_X1  g101(.A(KEYINPUT65), .B(KEYINPUT11), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n286), .B(new_n287), .C1(new_n282), .C2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n285), .B1(new_n289), .B2(G131), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n203), .A2(G143), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT64), .ZN(new_n293));
  INV_X1    g107(.A(G143), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n293), .B1(new_n294), .B2(G146), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n203), .A2(KEYINPUT64), .A3(G143), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n291), .B(new_n292), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT68), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT64), .B1(new_n203), .B2(G143), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n293), .A2(new_n294), .A3(G146), .ZN(new_n301));
  AOI22_X1  g115(.A1(new_n300), .A2(new_n301), .B1(G143), .B2(new_n203), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n302), .A2(KEYINPUT68), .A3(new_n292), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n294), .A2(G146), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n291), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT1), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n307), .B1(G143), .B2(new_n203), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n306), .B1(new_n220), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT70), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n306), .B(KEYINPUT70), .C1(new_n220), .C2(new_n308), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n290), .B1(new_n304), .B2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n302), .A2(KEYINPUT0), .A3(G128), .ZN(new_n315));
  NAND2_X1  g129(.A1(KEYINPUT0), .A2(G128), .ZN(new_n316));
  OR2_X1    g130(.A1(KEYINPUT0), .A2(G128), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n306), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT67), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G131), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n289), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n286), .A2(new_n287), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  XOR2_X1   g139(.A(KEYINPUT65), .B(KEYINPUT11), .Z(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT66), .B(G134), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n326), .B1(new_n327), .B2(G137), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n325), .A2(new_n321), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n319), .B1(new_n323), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n277), .B1(new_n314), .B2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(KEYINPUT68), .B1(new_n302), .B2(new_n292), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n300), .A2(new_n301), .ZN(new_n333));
  AND4_X1   g147(.A1(KEYINPUT68), .A2(new_n333), .A3(new_n291), .A4(new_n292), .ZN(new_n334));
  INV_X1    g148(.A(new_n312), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT1), .B1(new_n294), .B2(G146), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n231), .A2(G128), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n229), .A2(KEYINPUT69), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(KEYINPUT70), .B1(new_n339), .B2(new_n306), .ZN(new_n340));
  OAI22_X1  g154(.A1(new_n332), .A2(new_n334), .B1(new_n335), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G131), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n279), .A2(new_n281), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n283), .ZN(new_n344));
  INV_X1    g158(.A(new_n284), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n342), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n288), .B1(new_n283), .B2(new_n343), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n347), .A2(new_n324), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n346), .B1(new_n348), .B2(new_n342), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n341), .A2(new_n349), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n315), .A2(new_n318), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n321), .B1(new_n325), .B2(new_n328), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n289), .A2(new_n322), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n276), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(new_n273), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n350), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n269), .B1(new_n331), .B2(new_n357), .ZN(new_n358));
  NOR3_X1   g172(.A1(new_n314), .A2(new_n330), .A3(new_n277), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n359), .A2(KEYINPUT28), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n268), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  NOR3_X1   g175(.A1(new_n314), .A2(new_n330), .A3(KEYINPUT30), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT30), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n363), .B1(new_n350), .B2(new_n354), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n277), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(new_n267), .A3(new_n357), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT31), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n361), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G472), .ZN(new_n369));
  OAI21_X1  g183(.A(KEYINPUT30), .B1(new_n314), .B2(new_n330), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n350), .A2(new_n363), .A3(new_n354), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n356), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n372), .A2(new_n359), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(KEYINPUT31), .A3(new_n267), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n368), .A2(new_n369), .A3(new_n188), .A4(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT73), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT32), .ZN(new_n378));
  NOR3_X1   g192(.A1(new_n372), .A2(new_n268), .A3(new_n359), .ZN(new_n379));
  AOI21_X1  g193(.A(G902), .B1(new_n379), .B2(KEYINPUT31), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n380), .A2(new_n368), .A3(KEYINPUT73), .A4(new_n369), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n377), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n268), .B1(new_n372), .B2(new_n359), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n356), .B1(new_n350), .B2(new_n354), .ZN(new_n384));
  OAI21_X1  g198(.A(KEYINPUT28), .B1(new_n359), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n357), .A2(new_n269), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n267), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT29), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n383), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n188), .B1(new_n387), .B2(new_n388), .ZN(new_n390));
  OAI21_X1  g204(.A(G472), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n380), .A2(new_n368), .A3(KEYINPUT32), .A4(new_n369), .ZN(new_n392));
  AND2_X1   g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n262), .B1(new_n382), .B2(new_n393), .ZN(new_n394));
  XOR2_X1   g208(.A(G110), .B(G122), .Z(new_n395));
  INV_X1    g209(.A(KEYINPUT4), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT3), .ZN(new_n397));
  INV_X1    g211(.A(G104), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n397), .B1(new_n398), .B2(KEYINPUT79), .ZN(new_n399));
  INV_X1    g213(.A(G107), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(KEYINPUT80), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT80), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G107), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT79), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT3), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n399), .A2(new_n401), .A3(new_n403), .A4(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT3), .B1(new_n398), .B2(G107), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n398), .A2(G107), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G101), .ZN(new_n410));
  AOI21_X1  g224(.A(G101), .B1(new_n398), .B2(G107), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n406), .A2(new_n407), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n396), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(KEYINPUT4), .B1(new_n409), .B2(G101), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n277), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n272), .ZN(new_n416));
  XNOR2_X1  g230(.A(KEYINPUT88), .B(KEYINPUT5), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(G116), .A3(new_n222), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n418), .A2(G113), .ZN(new_n419));
  OR2_X1    g233(.A1(new_n274), .A2(new_n417), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n416), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(G104), .B1(new_n401), .B2(new_n403), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n398), .A2(G107), .ZN(new_n423));
  OAI21_X1  g237(.A(G101), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n412), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT81), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT89), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT81), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n412), .A2(new_n424), .A3(new_n428), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n421), .A2(new_n426), .A3(new_n427), .A4(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n415), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n421), .A2(new_n426), .A3(new_n429), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT89), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n395), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n395), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n433), .A2(new_n415), .A3(new_n436), .A4(new_n430), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n435), .A2(KEYINPUT6), .A3(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G953), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n214), .B1(new_n304), .B2(new_n313), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n319), .A2(new_n211), .ZN(new_n441));
  OAI211_X1 g255(.A(G224), .B(new_n439), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n341), .A2(new_n211), .ZN(new_n443));
  INV_X1    g257(.A(new_n441), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n439), .A2(G224), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT6), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n448), .B(new_n395), .C1(new_n431), .C2(new_n434), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n438), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT7), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n445), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n442), .A2(new_n446), .A3(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT90), .B(KEYINPUT8), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n395), .B(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n455), .B1(new_n421), .B2(new_n425), .ZN(new_n456));
  INV_X1    g270(.A(new_n419), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT91), .ZN(new_n458));
  AOI22_X1  g272(.A1(new_n457), .A2(new_n458), .B1(KEYINPUT5), .B2(new_n271), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n419), .A2(KEYINPUT91), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n416), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n456), .B1(new_n461), .B2(new_n425), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n443), .A2(new_n444), .A3(new_n451), .A4(new_n445), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n453), .A2(new_n462), .A3(new_n437), .A4(new_n463), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n464), .A2(new_n188), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n450), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(G210), .B1(G237), .B2(G902), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT92), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n450), .A2(new_n465), .A3(new_n467), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(G214), .B1(G237), .B2(G902), .ZN(new_n473));
  OR2_X1    g287(.A1(new_n471), .A2(new_n470), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT18), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT93), .B(G143), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n192), .A2(new_n477), .A3(G214), .A4(new_n263), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT72), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n439), .ZN(new_n480));
  NAND2_X1  g294(.A1(KEYINPUT72), .A2(G953), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n480), .A2(G214), .A3(new_n263), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(KEYINPUT93), .A2(G143), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI211_X1 g298(.A(new_n476), .B(new_n342), .C1(new_n478), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(KEYINPUT18), .A2(G131), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n478), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n207), .A2(G146), .A3(new_n209), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n248), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(KEYINPUT94), .B1(new_n485), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n478), .A2(new_n484), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(KEYINPUT18), .A3(G131), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT94), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n493), .A2(new_n494), .A3(new_n487), .A4(new_n489), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(G113), .B(G122), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(new_n398), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n492), .A2(G131), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT17), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n478), .A2(new_n484), .A3(new_n342), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n492), .A2(KEYINPUT17), .A3(G131), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n219), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n496), .A2(new_n498), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n498), .B1(new_n496), .B2(new_n504), .ZN(new_n506));
  NOR3_X1   g320(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT96), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(KEYINPUT96), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n188), .ZN(new_n509));
  OAI21_X1  g323(.A(G475), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT97), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT95), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n217), .A2(KEYINPUT19), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT19), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n247), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n513), .A2(new_n203), .A3(new_n515), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n516), .A2(new_n218), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n499), .A2(new_n501), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n498), .B1(new_n496), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n512), .B1(new_n505), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT20), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n496), .A2(new_n498), .A3(new_n504), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n491), .A2(new_n495), .B1(new_n517), .B2(new_n518), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n523), .B1(new_n498), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(G475), .A2(G902), .ZN(new_n526));
  AOI22_X1  g340(.A1(new_n521), .A2(new_n522), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AND4_X1   g341(.A1(KEYINPUT95), .A2(new_n525), .A3(new_n522), .A4(new_n526), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n510), .B(new_n511), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n510), .B1(new_n527), .B2(new_n528), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT97), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n220), .A2(G143), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n294), .A2(G128), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n532), .A2(new_n327), .A3(new_n533), .ZN(new_n534));
  OR2_X1    g348(.A1(new_n534), .A2(KEYINPUT98), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(KEYINPUT98), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n401), .A2(new_n403), .ZN(new_n537));
  XNOR2_X1  g351(.A(G116), .B(G122), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n537), .B(new_n538), .ZN(new_n539));
  XOR2_X1   g353(.A(new_n533), .B(KEYINPUT13), .Z(new_n540));
  INV_X1    g354(.A(new_n532), .ZN(new_n541));
  OAI21_X1  g355(.A(G134), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n535), .A2(new_n536), .A3(new_n539), .A4(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT14), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n538), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(G122), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n546), .A2(G116), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n400), .B1(new_n547), .B2(KEYINPUT14), .ZN(new_n548));
  AOI22_X1  g362(.A1(new_n545), .A2(new_n548), .B1(new_n537), .B2(new_n538), .ZN(new_n549));
  INV_X1    g363(.A(new_n534), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n327), .B1(new_n532), .B2(new_n533), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(KEYINPUT9), .B(G234), .ZN(new_n553));
  NOR3_X1   g367(.A1(new_n553), .A2(new_n187), .A3(G953), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n543), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n554), .B1(new_n543), .B2(new_n552), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n188), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT99), .ZN(new_n558));
  INV_X1    g372(.A(G478), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n559), .A2(KEYINPUT15), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT99), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n561), .B(new_n188), .C1(new_n555), .C2(new_n556), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n558), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  OR2_X1    g377(.A1(new_n557), .A2(new_n560), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(KEYINPUT100), .B(G952), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(G953), .ZN(new_n568));
  NAND2_X1  g382(.A1(G234), .A2(G237), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n192), .ZN(new_n572));
  AND3_X1   g386(.A1(new_n572), .A2(G902), .A3(new_n569), .ZN(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT21), .B(G898), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n571), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  AND4_X1   g390(.A1(new_n529), .A2(new_n531), .A3(new_n566), .A4(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(G221), .B1(new_n553), .B2(G902), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(KEYINPUT78), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n329), .A2(new_n323), .ZN(new_n580));
  XNOR2_X1  g394(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n304), .A2(new_n313), .A3(new_n425), .ZN(new_n582));
  INV_X1    g396(.A(new_n302), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n336), .A2(G128), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n425), .B1(new_n304), .B2(new_n585), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n580), .B(new_n581), .C1(new_n582), .C2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT83), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n304), .A2(new_n313), .A3(new_n425), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n299), .A2(new_n303), .B1(new_n583), .B2(new_n584), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n589), .B1(new_n425), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT83), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n591), .A2(new_n592), .A3(new_n580), .A4(new_n581), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n580), .B1(new_n582), .B2(new_n586), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT12), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n588), .A2(new_n593), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n351), .B1(new_n413), .B2(new_n414), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n341), .A2(KEYINPUT10), .A3(new_n426), .A4(new_n429), .ZN(new_n599));
  INV_X1    g413(.A(new_n580), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT10), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n601), .B1(new_n590), .B2(new_n425), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n598), .A2(new_n599), .A3(new_n600), .A4(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n192), .A2(G227), .ZN(new_n604));
  XOR2_X1   g418(.A(G110), .B(G140), .Z(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n603), .A2(KEYINPUT86), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(KEYINPUT86), .B1(new_n603), .B2(new_n607), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n597), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT87), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI211_X1 g426(.A(KEYINPUT87), .B(new_n597), .C1(new_n608), .C2(new_n609), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n598), .A2(new_n599), .A3(new_n602), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n614), .A2(KEYINPUT85), .A3(new_n580), .ZN(new_n615));
  AOI21_X1  g429(.A(KEYINPUT85), .B1(new_n614), .B2(new_n580), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n603), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n606), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n612), .A2(new_n613), .A3(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(G469), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n619), .A2(new_n620), .A3(new_n188), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n607), .B1(new_n597), .B2(new_n603), .ZN(new_n622));
  AND3_X1   g436(.A1(new_n603), .A2(KEYINPUT84), .A3(new_n607), .ZN(new_n623));
  INV_X1    g437(.A(new_n616), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n614), .A2(KEYINPUT85), .A3(new_n580), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n603), .A2(new_n607), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT84), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n622), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(G469), .B1(new_n630), .B2(G902), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n579), .B1(new_n621), .B2(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n394), .A2(new_n475), .A3(new_n577), .A4(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G101), .ZN(G3));
  AND3_X1   g448(.A1(new_n361), .A2(new_n367), .A3(new_n366), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n188), .B1(new_n366), .B2(new_n367), .ZN(new_n636));
  OAI21_X1  g450(.A(G472), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n377), .A2(new_n381), .A3(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n638), .A2(new_n262), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n632), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n531), .A2(new_n529), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n555), .A2(new_n556), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT33), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n555), .A2(new_n556), .A3(KEYINPUT33), .ZN(new_n645));
  OAI211_X1 g459(.A(G478), .B(new_n188), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n558), .A2(new_n559), .A3(new_n562), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n641), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n473), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n650), .B1(new_n469), .B2(new_n471), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n576), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n640), .A2(new_n649), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT34), .B(G104), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G6));
  INV_X1    g469(.A(new_n640), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n525), .A2(new_n526), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(new_n522), .ZN(new_n658));
  INV_X1    g472(.A(new_n510), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AND4_X1   g474(.A1(new_n565), .A2(new_n651), .A3(new_n576), .A4(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT35), .B(G107), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G9));
  AOI21_X1  g478(.A(new_n250), .B1(new_n240), .B2(new_n243), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT101), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT36), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n667), .B1(new_n201), .B2(new_n668), .ZN(new_n669));
  AOI211_X1 g483(.A(KEYINPUT101), .B(KEYINPUT36), .C1(new_n198), .C2(new_n200), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n666), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n669), .A2(new_n670), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n665), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n674), .A2(new_n261), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n665), .A2(new_n199), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n676), .B(new_n188), .C1(new_n665), .C2(new_n201), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n256), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n254), .A2(KEYINPUT25), .A3(new_n188), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n675), .B1(new_n680), .B2(new_n189), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n638), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n475), .A2(new_n577), .A3(new_n682), .A4(new_n632), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT37), .B(G110), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G12));
  AOI21_X1  g499(.A(new_n681), .B1(new_n382), .B2(new_n393), .ZN(new_n686));
  INV_X1    g500(.A(G900), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n571), .B1(new_n573), .B2(new_n687), .ZN(new_n688));
  NOR4_X1   g502(.A1(new_n658), .A2(new_n566), .A3(new_n659), .A4(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n686), .A2(new_n632), .A3(new_n651), .A4(new_n689), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT102), .B(G128), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G30));
  XOR2_X1   g506(.A(new_n688), .B(KEYINPUT39), .Z(new_n693));
  NAND2_X1  g507(.A1(new_n632), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(KEYINPUT104), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT40), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT104), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n694), .B(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT40), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n472), .A2(new_n474), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n701), .A2(KEYINPUT38), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT38), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n703), .B1(new_n472), .B2(new_n474), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n675), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n258), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n707), .A2(new_n650), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(new_n641), .A3(new_n565), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n380), .A2(new_n369), .A3(new_n368), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n267), .B1(new_n331), .B2(new_n357), .ZN(new_n711));
  OAI21_X1  g525(.A(KEYINPUT103), .B1(new_n379), .B2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT103), .ZN(new_n713));
  INV_X1    g527(.A(new_n711), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n366), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n712), .A2(new_n188), .A3(new_n715), .ZN(new_n716));
  AOI22_X1  g530(.A1(new_n710), .A2(KEYINPUT32), .B1(new_n716), .B2(G472), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n709), .B1(new_n382), .B2(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n697), .A2(new_n700), .A3(new_n705), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G143), .ZN(G45));
  INV_X1    g534(.A(new_n648), .ZN(new_n721));
  AOI211_X1 g535(.A(new_n721), .B(new_n688), .C1(new_n531), .C2(new_n529), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n686), .A2(new_n722), .A3(new_n632), .A4(new_n651), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G146), .ZN(G48));
  INV_X1    g538(.A(new_n652), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n619), .A2(new_n620), .A3(new_n188), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n620), .B1(new_n619), .B2(new_n188), .ZN(new_n727));
  INV_X1    g541(.A(new_n578), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n721), .B1(new_n531), .B2(new_n529), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n725), .A2(new_n729), .A3(new_n394), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(KEYINPUT41), .B(G113), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n731), .B(new_n732), .ZN(G15));
  NAND3_X1  g547(.A1(new_n661), .A2(new_n394), .A3(new_n729), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G116), .ZN(G18));
  NAND4_X1  g549(.A1(new_n729), .A2(new_n686), .A3(new_n577), .A4(new_n651), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G119), .ZN(G21));
  AND3_X1   g551(.A1(new_n641), .A2(new_n651), .A3(new_n565), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n637), .A2(new_n375), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n262), .A2(new_n739), .A3(new_n575), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n738), .A2(new_n729), .A3(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G122), .ZN(G24));
  INV_X1    g556(.A(KEYINPUT105), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n743), .B1(new_n739), .B2(new_n681), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n707), .A2(KEYINPUT105), .A3(new_n375), .A4(new_n637), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n746), .A2(new_n729), .A3(new_n651), .A4(new_n722), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G125), .ZN(G27));
  NAND2_X1  g562(.A1(new_n391), .A2(new_n392), .ZN(new_n749));
  AOI21_X1  g563(.A(KEYINPUT107), .B1(new_n375), .B2(new_n378), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n375), .A2(KEYINPUT107), .A3(new_n378), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n262), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n650), .B1(new_n472), .B2(new_n474), .ZN(new_n754));
  AOI21_X1  g568(.A(KEYINPUT106), .B1(new_n630), .B2(G469), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n597), .A2(new_n603), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n606), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n603), .A2(KEYINPUT84), .A3(new_n607), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n629), .B(new_n758), .C1(new_n616), .C2(new_n615), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n757), .A2(new_n759), .A3(KEYINPUT106), .A4(G469), .ZN(new_n760));
  NAND2_X1  g574(.A1(G469), .A2(G902), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n755), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n728), .B1(new_n763), .B2(new_n621), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n753), .A2(new_n722), .A3(new_n754), .A4(new_n764), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n764), .A2(new_n394), .A3(new_n754), .ZN(new_n766));
  INV_X1    g580(.A(new_n722), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(KEYINPUT42), .ZN(new_n768));
  AOI22_X1  g582(.A1(KEYINPUT42), .A2(new_n765), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G131), .ZN(G33));
  AND2_X1   g584(.A1(new_n394), .A2(new_n754), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n771), .A2(KEYINPUT108), .A3(new_n689), .A4(new_n764), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n764), .A2(new_n394), .A3(new_n689), .A4(new_n754), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT108), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G134), .ZN(G36));
  NAND2_X1  g591(.A1(new_n757), .A2(new_n759), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT45), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n620), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT109), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n630), .A2(KEYINPUT45), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n784), .B1(new_n780), .B2(new_n781), .ZN(new_n785));
  OAI211_X1 g599(.A(KEYINPUT46), .B(new_n761), .C1(new_n783), .C2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n621), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n780), .A2(new_n781), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n788), .A2(new_n782), .A3(new_n784), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT46), .B1(new_n789), .B2(new_n761), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT110), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n791), .A2(new_n792), .A3(new_n578), .A4(new_n693), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n578), .B1(new_n787), .B2(new_n790), .ZN(new_n794));
  INV_X1    g608(.A(new_n693), .ZN(new_n795));
  OAI21_X1  g609(.A(KEYINPUT110), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n531), .A2(new_n529), .A3(new_n648), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT43), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT43), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n531), .A2(new_n799), .A3(new_n529), .A4(new_n648), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n638), .A2(new_n707), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT44), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AND4_X1   g618(.A1(KEYINPUT44), .A2(new_n803), .A3(new_n798), .A4(new_n800), .ZN(new_n805));
  INV_X1    g619(.A(new_n754), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n793), .A2(new_n796), .A3(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G137), .ZN(G39));
  XNOR2_X1  g623(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n791), .A2(new_n578), .A3(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n810), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n794), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n382), .A2(new_n393), .A3(new_n262), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n767), .A2(new_n806), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n811), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G140), .ZN(G42));
  NAND3_X1  g631(.A1(new_n729), .A2(new_n571), .A3(new_n754), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n818), .A2(new_n801), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT118), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT48), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n819), .A2(new_n753), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n822), .B1(new_n819), .B2(new_n753), .ZN(new_n824));
  OAI22_X1  g638(.A1(new_n823), .A2(new_n824), .B1(new_n820), .B2(new_n821), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n262), .A2(new_n739), .A3(new_n570), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n802), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n729), .A2(new_n651), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n568), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n262), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n830), .A2(new_n382), .A3(new_n717), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n818), .A2(new_n649), .A3(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n825), .A2(new_n833), .ZN(new_n834));
  OR2_X1    g648(.A1(new_n702), .A2(new_n704), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n835), .A2(KEYINPUT115), .A3(new_n650), .A4(new_n729), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT115), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n729), .A2(new_n650), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n837), .B1(new_n705), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n827), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n840), .A2(KEYINPUT50), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT50), .ZN(new_n842));
  AOI211_X1 g656(.A(new_n842), .B(new_n827), .C1(new_n836), .C2(new_n839), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n819), .A2(new_n746), .ZN(new_n845));
  NOR4_X1   g659(.A1(new_n818), .A2(new_n641), .A3(new_n648), .A4(new_n831), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n845), .A2(new_n846), .A3(KEYINPUT117), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n845), .A2(new_n846), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT117), .ZN(new_n849));
  OAI21_X1  g663(.A(KEYINPUT51), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n844), .A2(new_n847), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n827), .A2(new_n806), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n794), .B(new_n810), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n726), .A2(new_n727), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n854), .A2(new_n579), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n852), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n834), .B1(new_n851), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n848), .B1(new_n841), .B2(new_n843), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT116), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT114), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n856), .A2(new_n861), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n848), .B(KEYINPUT116), .C1(new_n841), .C2(new_n843), .ZN(new_n863));
  OAI211_X1 g677(.A(KEYINPUT114), .B(new_n852), .C1(new_n853), .C2(new_n855), .ZN(new_n864));
  AND4_X1   g678(.A1(new_n860), .A2(new_n862), .A3(new_n863), .A4(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n857), .B1(new_n865), .B2(KEYINPUT51), .ZN(new_n866));
  INV_X1    g680(.A(new_n688), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n258), .A2(new_n706), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n868), .B1(new_n382), .B2(new_n717), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n738), .A2(new_n764), .A3(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n747), .A2(new_n870), .A3(new_n723), .A4(new_n690), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT52), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT112), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OR2_X1    g689(.A1(new_n871), .A2(new_n872), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n871), .A2(KEYINPUT112), .A3(new_n872), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n746), .A2(new_n764), .A3(new_n722), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n565), .A2(new_n688), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n686), .A2(new_n632), .A3(new_n660), .A4(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n754), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n769), .A2(new_n776), .A3(new_n885), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n731), .A2(new_n633), .A3(new_n741), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n734), .A2(new_n736), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n531), .A2(new_n529), .A3(new_n565), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n575), .B1(new_n649), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n656), .A2(new_n475), .A3(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n887), .A2(new_n888), .A3(new_n891), .A4(new_n683), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n886), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT53), .B1(new_n880), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n890), .A2(new_n475), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n734), .B(new_n736), .C1(new_n895), .C2(new_n640), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n731), .A2(new_n633), .A3(new_n741), .A4(new_n683), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n898), .A2(new_n769), .A3(new_n776), .A4(new_n885), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n871), .B(KEYINPUT52), .ZN(new_n900));
  XOR2_X1   g714(.A(KEYINPUT113), .B(KEYINPUT53), .Z(new_n901));
  NOR3_X1   g715(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(KEYINPUT54), .B1(new_n894), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT112), .B1(new_n871), .B2(new_n872), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n871), .A2(new_n872), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n893), .B(KEYINPUT53), .C1(new_n906), .C2(new_n878), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT54), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n901), .B1(new_n899), .B2(new_n900), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n903), .A2(new_n910), .ZN(new_n911));
  OAI22_X1  g725(.A1(new_n866), .A2(new_n911), .B1(G952), .B2(G953), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n854), .B(KEYINPUT49), .ZN(new_n913));
  NOR4_X1   g727(.A1(new_n831), .A2(new_n579), .A3(new_n650), .A4(new_n797), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n835), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n912), .A2(new_n915), .ZN(G75));
  NAND2_X1  g730(.A1(new_n907), .A2(new_n909), .ZN(new_n917));
  NAND2_X1  g731(.A1(G210), .A2(G902), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT56), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n438), .A2(new_n449), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(new_n447), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT55), .Z(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n920), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n192), .A2(G952), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n918), .B1(new_n907), .B2(new_n909), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n923), .B1(new_n928), .B2(KEYINPUT56), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n925), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT119), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n925), .A2(KEYINPUT119), .A3(new_n927), .A4(new_n929), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(G51));
  NAND2_X1  g748(.A1(new_n917), .A2(KEYINPUT54), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n910), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n761), .B(KEYINPUT57), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n619), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n188), .B1(new_n907), .B2(new_n909), .ZN(new_n940));
  INV_X1    g754(.A(new_n789), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n926), .B1(new_n939), .B2(new_n942), .ZN(G54));
  AND2_X1   g757(.A1(KEYINPUT58), .A2(G475), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n940), .A2(new_n525), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n525), .B1(new_n940), .B2(new_n944), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n945), .A2(new_n946), .A3(new_n926), .ZN(G60));
  NAND2_X1  g761(.A1(G478), .A2(G902), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT59), .Z(new_n949));
  AOI21_X1  g763(.A(new_n949), .B1(new_n903), .B2(new_n910), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n644), .A2(new_n645), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(KEYINPUT120), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n949), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT53), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n906), .A2(new_n878), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n955), .B1(new_n956), .B2(new_n899), .ZN(new_n957));
  OR3_X1    g771(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n908), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n954), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT120), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n961), .A2(new_n962), .A3(new_n951), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n951), .A2(new_n949), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n926), .B1(new_n936), .B2(new_n964), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n953), .A2(new_n963), .A3(new_n965), .ZN(G63));
  NAND2_X1  g780(.A1(G217), .A2(G902), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT60), .Z(new_n968));
  NAND2_X1  g782(.A1(new_n917), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n259), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n917), .A2(new_n673), .A3(new_n671), .A4(new_n968), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n970), .A2(new_n927), .A3(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT61), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n970), .A2(KEYINPUT61), .A3(new_n927), .A4(new_n971), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(G66));
  INV_X1    g790(.A(G224), .ZN(new_n977));
  OAI21_X1  g791(.A(G953), .B1(new_n574), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n978), .B1(new_n898), .B2(new_n572), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT121), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n921), .B1(G898), .B2(new_n192), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n980), .B(new_n981), .ZN(G69));
  AND3_X1   g796(.A1(new_n747), .A2(new_n690), .A3(new_n723), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n719), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(KEYINPUT62), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n649), .A2(new_n889), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n695), .A2(new_n771), .A3(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT62), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n719), .A2(new_n988), .A3(new_n983), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n985), .A2(new_n987), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n808), .A2(new_n816), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n192), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n362), .A2(new_n364), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n513), .A2(new_n515), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n993), .B(new_n994), .Z(new_n995));
  AOI21_X1  g809(.A(new_n192), .B1(G227), .B2(G900), .ZN(new_n996));
  AOI22_X1  g810(.A1(new_n992), .A2(new_n995), .B1(KEYINPUT124), .B2(new_n996), .ZN(new_n997));
  AND2_X1   g811(.A1(new_n808), .A2(new_n816), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT122), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n773), .B(KEYINPUT108), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n765), .A2(KEYINPUT42), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n766), .A2(new_n768), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n999), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n769), .A2(new_n776), .A3(KEYINPUT122), .ZN(new_n1005));
  AND3_X1   g819(.A1(new_n1004), .A2(new_n1005), .A3(new_n983), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT123), .ZN(new_n1007));
  AND2_X1   g821(.A1(new_n753), .A2(new_n738), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n793), .A2(new_n796), .A3(new_n1008), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n998), .A2(new_n1006), .A3(new_n1007), .A4(new_n1009), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n1009), .A2(new_n1005), .A3(new_n983), .A4(new_n1004), .ZN(new_n1011));
  OAI21_X1  g825(.A(KEYINPUT123), .B1(new_n1011), .B2(new_n991), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1010), .A2(new_n1012), .A3(new_n192), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n995), .B1(G900), .B2(new_n572), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  OR2_X1    g829(.A1(new_n996), .A2(KEYINPUT124), .ZN(new_n1016));
  AND3_X1   g830(.A1(new_n997), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1016), .B1(new_n997), .B2(new_n1015), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1017), .A2(new_n1018), .ZN(G72));
  NAND3_X1  g833(.A1(new_n1010), .A2(new_n1012), .A3(new_n898), .ZN(new_n1020));
  XNOR2_X1  g834(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n369), .A2(new_n188), .ZN(new_n1022));
  XNOR2_X1  g836(.A(new_n1021), .B(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g837(.A(new_n1023), .B(KEYINPUT126), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n1025), .A2(new_n268), .A3(new_n373), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n373), .A2(new_n268), .ZN(new_n1027));
  NOR3_X1   g841(.A1(new_n990), .A2(new_n892), .A3(new_n991), .ZN(new_n1028));
  INV_X1    g842(.A(new_n1024), .ZN(new_n1029));
  OAI211_X1 g843(.A(KEYINPUT127), .B(new_n1027), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1030));
  INV_X1    g844(.A(KEYINPUT127), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n989), .A2(new_n987), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n988), .B1(new_n719), .B2(new_n983), .ZN(new_n1033));
  NOR3_X1   g847(.A1(new_n1032), .A2(new_n991), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n1029), .B1(new_n1034), .B2(new_n898), .ZN(new_n1035));
  INV_X1    g849(.A(new_n1027), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1031), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n957), .A2(new_n958), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n1023), .B1(new_n383), .B2(new_n366), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n926), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  AND4_X1   g854(.A1(new_n1026), .A2(new_n1030), .A3(new_n1037), .A4(new_n1040), .ZN(G57));
endmodule


