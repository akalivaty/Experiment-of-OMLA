//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 1 1 1 0 0 0 1 1 0 0 0 1 1 0 1 0 0 1 1 0 0 0 1 0 1 0 1 0 1 0 1 0 1 0 1 1 1 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1238, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  INV_X1    g0010(.A(new_n201), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  INV_X1    g0020(.A(G107), .ZN(new_n221));
  INV_X1    g0021(.A(G264), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n207), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n210), .B(new_n217), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XOR2_X1   g0038(.A(G107), .B(G116), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT66), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT65), .ZN(new_n243));
  XOR2_X1   g0043(.A(G58), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(KEYINPUT3), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G33), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n250));
  AND3_X1   g0050(.A1(new_n248), .A2(new_n250), .A3(KEYINPUT68), .ZN(new_n251));
  AOI21_X1  g0051(.A(KEYINPUT68), .B1(new_n248), .B2(new_n250), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G1698), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n253), .A2(G222), .A3(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n253), .A2(G223), .A3(G1698), .ZN(new_n256));
  OAI211_X1 g0056(.A(new_n255), .B(new_n256), .C1(new_n219), .C2(new_n253), .ZN(new_n257));
  AND2_X1   g0057(.A1(G1), .A2(G13), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT69), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  AND3_X1   g0060(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n259), .B1(new_n258), .B2(new_n260), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G274), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n265), .B1(new_n258), .B2(new_n260), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(G41), .B2(G45), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G226), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n258), .A2(new_n260), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n268), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n270), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  XOR2_X1   g0074(.A(new_n274), .B(KEYINPUT67), .Z(new_n275));
  AND2_X1   g0075(.A1(new_n264), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G190), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n264), .A2(new_n275), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G200), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n214), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT8), .B(G58), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n249), .A2(G20), .ZN(new_n285));
  NOR2_X1   g0085(.A1(G20), .A2(G33), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n284), .A2(new_n285), .B1(G150), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n203), .A2(G20), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n282), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G13), .ZN(new_n290));
  NOR3_X1   g0090(.A1(new_n290), .A2(new_n215), .A3(G1), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n291), .A2(new_n281), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n267), .A2(G20), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n292), .A2(G50), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n291), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n294), .B1(G50), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n289), .A2(new_n296), .ZN(new_n297));
  XOR2_X1   g0097(.A(new_n297), .B(KEYINPUT9), .Z(new_n298));
  NAND3_X1  g0098(.A1(new_n277), .A2(new_n279), .A3(new_n298), .ZN(new_n299));
  XOR2_X1   g0099(.A(new_n299), .B(KEYINPUT10), .Z(new_n300));
  INV_X1    g0100(.A(KEYINPUT70), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT68), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n247), .A2(G33), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n248), .A2(new_n250), .A3(KEYINPUT68), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n305), .A2(G226), .A3(new_n254), .A4(new_n306), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n305), .A2(G232), .A3(G1698), .A4(new_n306), .ZN(new_n308));
  NAND2_X1  g0108(.A1(G33), .A2(G97), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n263), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT13), .ZN(new_n312));
  INV_X1    g0112(.A(new_n270), .ZN(new_n313));
  INV_X1    g0113(.A(new_n273), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n313), .B1(G238), .B2(new_n314), .ZN(new_n315));
  AND3_X1   g0115(.A1(new_n311), .A2(new_n312), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n312), .B1(new_n311), .B2(new_n315), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G200), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n301), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n317), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n311), .A2(new_n312), .A3(new_n315), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n323), .A2(KEYINPUT70), .A3(G200), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n320), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n286), .A2(G50), .ZN(new_n326));
  XNOR2_X1  g0126(.A(new_n326), .B(KEYINPUT71), .ZN(new_n327));
  INV_X1    g0127(.A(G68), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n285), .A2(G77), .B1(G20), .B2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n282), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  OR2_X1    g0130(.A1(new_n330), .A2(KEYINPUT11), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(KEYINPUT11), .ZN(new_n332));
  OR3_X1    g0132(.A1(new_n295), .A2(KEYINPUT12), .A3(G68), .ZN(new_n333));
  OAI21_X1  g0133(.A(KEYINPUT12), .B1(new_n295), .B2(G68), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n328), .B1(new_n267), .B2(G20), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n333), .A2(new_n334), .B1(new_n292), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n331), .A2(new_n332), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n337), .B1(new_n318), .B2(G190), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n325), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G179), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n276), .A2(new_n341), .ZN(new_n342));
  OAI221_X1 g0142(.A(new_n342), .B1(G169), .B2(new_n276), .C1(new_n289), .C2(new_n296), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n270), .B1(new_n220), .B2(new_n273), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n253), .A2(G232), .A3(new_n254), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n253), .A2(G238), .A3(G1698), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n345), .B(new_n346), .C1(new_n221), .C2(new_n253), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n344), .B1(new_n347), .B2(new_n263), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G200), .ZN(new_n350));
  INV_X1    g0150(.A(new_n292), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n293), .A2(G77), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n353), .B1(new_n219), .B2(new_n291), .ZN(new_n354));
  XNOR2_X1  g0154(.A(KEYINPUT15), .B(G87), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n285), .ZN(new_n357));
  INV_X1    g0157(.A(new_n286), .ZN(new_n358));
  OAI221_X1 g0158(.A(new_n357), .B1(new_n215), .B2(new_n219), .C1(new_n358), .C2(new_n283), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n281), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n354), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n361), .B1(new_n348), .B2(G190), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n350), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G169), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n349), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n348), .A2(new_n341), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n365), .A2(new_n366), .A3(new_n361), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n343), .A2(new_n363), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT14), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n369), .B(G169), .C1(new_n316), .C2(new_n317), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(new_n323), .B2(new_n341), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n369), .B1(new_n323), .B2(G169), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n337), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  NOR4_X1   g0174(.A1(new_n300), .A2(new_n340), .A3(new_n368), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(G58), .A2(G68), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n211), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT73), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(new_n378), .A3(G20), .ZN(new_n379));
  INV_X1    g0179(.A(G159), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n379), .B1(new_n380), .B2(new_n358), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n378), .B1(new_n377), .B2(G20), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT7), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n384), .A2(KEYINPUT72), .ZN(new_n385));
  XNOR2_X1  g0185(.A(KEYINPUT3), .B(G33), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n385), .B1(new_n386), .B2(G20), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n248), .A2(new_n250), .ZN(new_n388));
  XNOR2_X1  g0188(.A(KEYINPUT72), .B(KEYINPUT7), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(new_n389), .A3(new_n215), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n387), .A2(new_n390), .A3(G68), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n383), .A2(KEYINPUT16), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n281), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n215), .B1(new_n251), .B2(new_n252), .ZN(new_n394));
  OR3_X1    g0194(.A1(new_n249), .A2(KEYINPUT74), .A3(KEYINPUT3), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n248), .A2(KEYINPUT74), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n395), .A2(new_n396), .A3(new_n250), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n384), .A2(G20), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n394), .A2(new_n384), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(KEYINPUT75), .B1(new_n399), .B2(new_n328), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n397), .A2(new_n398), .ZN(new_n401));
  AOI21_X1  g0201(.A(G20), .B1(new_n305), .B2(new_n306), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n401), .B1(new_n402), .B2(KEYINPUT7), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT75), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n403), .A2(new_n404), .A3(G68), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n400), .A2(new_n383), .A3(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT16), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n393), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n284), .A2(new_n293), .ZN(new_n409));
  OAI22_X1  g0209(.A1(new_n351), .A2(new_n409), .B1(new_n295), .B2(new_n284), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n271), .A2(G1698), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n386), .B(new_n412), .C1(G223), .C2(G1698), .ZN(new_n413));
  INV_X1    g0213(.A(G87), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n413), .B1(new_n249), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n263), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n313), .B1(G232), .B2(new_n314), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(G190), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n319), .B1(new_n416), .B2(new_n417), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n411), .A2(KEYINPUT17), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n410), .ZN(new_n424));
  OR2_X1    g0224(.A1(new_n381), .A2(new_n382), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n403), .A2(G68), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n425), .B1(new_n426), .B2(KEYINPUT75), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT16), .B1(new_n427), .B2(new_n405), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n422), .B(new_n424), .C1(new_n428), .C2(new_n393), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT17), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n423), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT18), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n424), .B1(new_n428), .B2(new_n393), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n418), .A2(G169), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(new_n341), .B2(new_n418), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n433), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n433), .B(new_n436), .C1(new_n408), .C2(new_n410), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT76), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n436), .B1(new_n408), .B2(new_n410), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT18), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT76), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(new_n443), .A3(new_n438), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n432), .B1(new_n440), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n375), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NOR3_X1   g0247(.A1(new_n414), .A2(KEYINPUT22), .A3(G20), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n253), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n386), .A2(new_n215), .A3(G87), .ZN(new_n450));
  AND3_X1   g0250(.A1(new_n450), .A2(KEYINPUT86), .A3(KEYINPUT22), .ZN(new_n451));
  AOI21_X1  g0251(.A(KEYINPUT86), .B1(new_n450), .B2(KEYINPUT22), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n449), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT24), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT23), .B1(new_n221), .B2(G20), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n221), .A2(KEYINPUT23), .A3(G20), .ZN(new_n457));
  INV_X1    g0257(.A(G116), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n249), .A2(new_n458), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n456), .A2(new_n457), .B1(new_n459), .B2(new_n215), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n453), .A2(new_n454), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n454), .B1(new_n453), .B2(new_n460), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n281), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(G45), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(G1), .ZN(new_n465));
  XNOR2_X1  g0265(.A(KEYINPUT5), .B(G41), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n266), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n465), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n272), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n272), .A2(KEYINPUT69), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(G250), .A2(G1698), .ZN(new_n473));
  INV_X1    g0273(.A(G257), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n473), .B1(new_n474), .B2(G1698), .ZN(new_n475));
  AOI22_X1  g0275(.A1(new_n475), .A2(new_n386), .B1(G33), .B2(G294), .ZN(new_n476));
  OAI221_X1 g0276(.A(new_n467), .B1(new_n469), .B2(new_n222), .C1(new_n472), .C2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n477), .A2(new_n419), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n478), .B1(G200), .B2(new_n477), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n292), .B1(G1), .B2(new_n249), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT25), .B1(new_n291), .B2(new_n221), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n291), .A2(KEYINPUT25), .A3(new_n221), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n481), .A2(G107), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AND3_X1   g0285(.A1(new_n463), .A2(new_n479), .A3(new_n485), .ZN(new_n486));
  OR2_X1    g0286(.A1(new_n477), .A2(G179), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n477), .A2(new_n364), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n489), .B1(new_n463), .B2(new_n485), .ZN(new_n490));
  OAI21_X1  g0290(.A(KEYINPUT87), .B1(new_n486), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT87), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n463), .A2(new_n479), .A3(new_n485), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n453), .A2(new_n460), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT24), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n453), .A2(new_n454), .A3(new_n460), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n282), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n485), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n492), .B(new_n493), .C1(new_n499), .C2(new_n489), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n491), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(G303), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n253), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT84), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G264), .A2(G1698), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n504), .B1(new_n388), .B2(new_n505), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n386), .A2(KEYINPUT84), .A3(G264), .A4(G1698), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n386), .A2(G257), .A3(new_n254), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n263), .B1(new_n503), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n467), .ZN(new_n511));
  INV_X1    g0311(.A(new_n469), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n511), .B1(new_n512), .B2(G270), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G33), .A2(G283), .ZN(new_n516));
  INV_X1    g0316(.A(G97), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n516), .B(new_n215), .C1(G33), .C2(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n518), .B(new_n281), .C1(new_n215), .C2(G116), .ZN(new_n519));
  XNOR2_X1  g0319(.A(new_n519), .B(KEYINPUT20), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n291), .A2(new_n458), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(new_n480), .B2(new_n458), .ZN(new_n522));
  OAI21_X1  g0322(.A(G169), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(KEYINPUT85), .B1(new_n515), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT21), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT21), .ZN(new_n526));
  OAI211_X1 g0326(.A(KEYINPUT85), .B(new_n526), .C1(new_n515), .C2(new_n523), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n510), .A2(G179), .A3(new_n513), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n520), .A2(new_n522), .ZN(new_n529));
  OR2_X1    g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n514), .A2(G200), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n531), .B(new_n529), .C1(new_n419), .C2(new_n514), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n525), .A2(new_n527), .A3(new_n530), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n403), .A2(G107), .ZN(new_n534));
  OR3_X1    g0334(.A1(new_n517), .A2(KEYINPUT78), .A3(G107), .ZN(new_n535));
  OAI21_X1  g0335(.A(KEYINPUT78), .B1(new_n517), .B2(G107), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT6), .ZN(new_n538));
  AOI22_X1  g0338(.A1(KEYINPUT77), .A2(new_n538), .B1(new_n517), .B2(G107), .ZN(new_n539));
  OR2_X1    g0339(.A1(new_n538), .A2(KEYINPUT77), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n535), .A2(new_n539), .A3(new_n536), .A4(new_n540), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n544), .A2(G20), .B1(G77), .B2(new_n286), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n282), .B1(new_n534), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n295), .A2(G97), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n547), .B1(new_n481), .B2(G97), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n467), .B1(new_n469), .B2(new_n474), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n305), .A2(G250), .A3(G1698), .A4(new_n306), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT4), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n553), .A2(new_n220), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n305), .A2(new_n254), .A3(new_n306), .A4(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n386), .A2(G244), .A3(new_n254), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n553), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n552), .A2(new_n555), .A3(new_n557), .A4(new_n516), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n551), .B1(new_n558), .B2(new_n263), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(G190), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n550), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n551), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT79), .ZN(new_n563));
  AND3_X1   g0363(.A1(new_n558), .A2(new_n563), .A3(new_n263), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n563), .B1(new_n558), .B2(new_n263), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n562), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G200), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n534), .A2(new_n545), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n281), .ZN(new_n569));
  INV_X1    g0369(.A(new_n559), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n569), .A2(new_n548), .B1(new_n364), .B2(new_n570), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n341), .B(new_n562), .C1(new_n564), .C2(new_n565), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n561), .A2(new_n567), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT80), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n533), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n567), .A2(new_n550), .A3(new_n560), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n571), .A2(new_n572), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT83), .ZN(new_n579));
  INV_X1    g0379(.A(G250), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n580), .B1(new_n267), .B2(G45), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n266), .A2(new_n465), .B1(new_n272), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(G238), .A2(G1698), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n583), .B1(new_n220), .B2(G1698), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n459), .B1(new_n584), .B2(new_n386), .ZN(new_n585));
  OAI211_X1 g0385(.A(G190), .B(new_n582), .C1(new_n585), .C2(new_n472), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n220), .A2(G1698), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(G238), .B2(G1698), .ZN(new_n589));
  OAI22_X1  g0389(.A1(new_n589), .A2(new_n388), .B1(new_n249), .B2(new_n458), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n263), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n319), .B1(new_n591), .B2(new_n582), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n587), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n481), .A2(G87), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT82), .ZN(new_n595));
  NOR3_X1   g0395(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n596));
  AOI21_X1  g0396(.A(G20), .B1(G33), .B2(G97), .ZN(new_n597));
  OAI21_X1  g0397(.A(KEYINPUT19), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT19), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n285), .A2(new_n599), .A3(G97), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n386), .A2(KEYINPUT81), .A3(new_n215), .A4(G68), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n248), .A2(new_n250), .A3(new_n215), .A4(G68), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT81), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n601), .A2(new_n602), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n281), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n356), .A2(new_n295), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n595), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  AOI211_X1 g0410(.A(KEYINPUT82), .B(new_n608), .C1(new_n606), .C2(new_n281), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n593), .B(new_n594), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n266), .A2(new_n465), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n272), .A2(new_n581), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(new_n263), .B2(new_n590), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n341), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n591), .A2(new_n582), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n364), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n598), .A2(new_n600), .B1(new_n603), .B2(new_n604), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n282), .B1(new_n622), .B2(new_n602), .ZN(new_n623));
  OAI21_X1  g0423(.A(KEYINPUT82), .B1(new_n623), .B2(new_n608), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n607), .A2(new_n595), .A3(new_n609), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n481), .A2(new_n356), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n621), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n579), .B1(new_n613), .B2(new_n628), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n624), .A2(new_n625), .B1(new_n356), .B2(new_n481), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n612), .B(KEYINPUT83), .C1(new_n630), .C2(new_n621), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n578), .A2(KEYINPUT80), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  AND4_X1   g0432(.A1(new_n447), .A2(new_n501), .A3(new_n575), .A4(new_n632), .ZN(G372));
  INV_X1    g0433(.A(new_n343), .ZN(new_n634));
  XNOR2_X1  g0434(.A(new_n300), .B(KEYINPUT91), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n437), .A2(new_n439), .ZN(new_n636));
  INV_X1    g0436(.A(new_n366), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n361), .B1(new_n348), .B2(G169), .ZN(new_n638));
  OAI21_X1  g0438(.A(KEYINPUT90), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT90), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n365), .A2(new_n640), .A3(new_n366), .A4(new_n361), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n374), .B1(new_n339), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n636), .B1(new_n643), .B2(new_n432), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n634), .B1(new_n635), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n627), .B1(new_n610), .B2(new_n611), .ZN(new_n646));
  INV_X1    g0446(.A(new_n621), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT88), .ZN(new_n649));
  INV_X1    g0449(.A(new_n572), .ZN(new_n650));
  OAI22_X1  g0450(.A1(new_n546), .A2(new_n549), .B1(G169), .B2(new_n559), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n613), .A2(new_n628), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT26), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n569), .A2(new_n548), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n570), .A2(new_n364), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n655), .A2(new_n572), .A3(KEYINPUT88), .A4(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n652), .A2(new_n653), .A3(new_n654), .A4(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n577), .B1(new_n629), .B2(new_n631), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n648), .B(new_n658), .C1(new_n659), .C2(new_n654), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(KEYINPUT89), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n650), .A2(new_n651), .ZN(new_n662));
  INV_X1    g0462(.A(new_n631), .ZN(new_n663));
  AOI21_X1  g0463(.A(KEYINPUT83), .B1(new_n648), .B2(new_n612), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(KEYINPUT26), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT89), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n666), .A2(new_n667), .A3(new_n648), .A4(new_n658), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n648), .A2(new_n612), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n486), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n525), .A2(new_n527), .A3(new_n530), .ZN(new_n671));
  OAI211_X1 g0471(.A(new_n670), .B(new_n573), .C1(new_n490), .C2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n661), .A2(new_n668), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n645), .B1(new_n446), .B2(new_n674), .ZN(G369));
  NAND3_X1  g0475(.A1(new_n267), .A2(new_n215), .A3(G13), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT92), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT27), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(new_n680), .A3(G213), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  XNOR2_X1  g0482(.A(KEYINPUT93), .B(G343), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n682), .A2(KEYINPUT94), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT94), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n681), .B2(new_n683), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(new_n497), .B2(new_n498), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT95), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n501), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n688), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n671), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  AOI22_X1  g0494(.A1(new_n691), .A2(new_n694), .B1(new_n490), .B2(new_n692), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n691), .B1(new_n490), .B2(new_n688), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n692), .A2(new_n529), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n671), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n533), .B2(new_n697), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(G330), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n695), .B1(new_n696), .B2(new_n700), .ZN(G399));
  INV_X1    g0501(.A(new_n208), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(G41), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n596), .A2(new_n458), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n704), .A2(G1), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(new_n212), .B2(new_n704), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT28), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n628), .B(KEYINPUT99), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n672), .B(new_n710), .C1(KEYINPUT26), .C2(new_n665), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n669), .B1(new_n577), .B2(new_n649), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n654), .B1(new_n712), .B2(new_n657), .ZN(new_n713));
  OAI211_X1 g0513(.A(KEYINPUT29), .B(new_n692), .C1(new_n711), .C2(new_n713), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n673), .A2(new_n692), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n714), .B1(new_n715), .B2(KEYINPUT29), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n632), .A2(new_n575), .A3(new_n501), .A4(new_n692), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n476), .A2(new_n472), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n718), .B1(G264), .B2(new_n512), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n559), .A2(new_n719), .A3(new_n617), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT30), .ZN(new_n721));
  OR3_X1    g0521(.A1(new_n720), .A2(new_n528), .A3(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n617), .A2(G179), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n566), .A2(new_n477), .A3(new_n514), .A4(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n721), .B1(new_n720), .B2(new_n528), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n722), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g0526(.A(KEYINPUT96), .B(KEYINPUT31), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n726), .A2(new_n688), .A3(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT97), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n725), .A2(new_n730), .ZN(new_n731));
  OAI211_X1 g0531(.A(KEYINPUT97), .B(new_n721), .C1(new_n720), .C2(new_n528), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n731), .A2(new_n722), .A3(new_n732), .A4(new_n724), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(new_n688), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT31), .ZN(new_n735));
  AOI21_X1  g0535(.A(KEYINPUT98), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n734), .A2(new_n735), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT98), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  OAI211_X1 g0539(.A(new_n717), .B(new_n729), .C1(new_n736), .C2(new_n739), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n740), .A2(G330), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AND2_X1   g0542(.A1(new_n716), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n709), .B1(new_n743), .B2(G1), .ZN(G364));
  NOR2_X1   g0544(.A1(new_n699), .A2(G330), .ZN(new_n745));
  XOR2_X1   g0545(.A(new_n745), .B(KEYINPUT100), .Z(new_n746));
  NOR2_X1   g0546(.A1(new_n290), .A2(G20), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n267), .B1(new_n747), .B2(G45), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n703), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n746), .A2(new_n700), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n253), .A2(new_n208), .ZN(new_n753));
  INV_X1    g0553(.A(G355), .ZN(new_n754));
  OAI22_X1  g0554(.A1(new_n753), .A2(new_n754), .B1(G116), .B2(new_n208), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n245), .A2(G45), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n702), .A2(new_n386), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n758), .B1(new_n464), .B2(new_n213), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n755), .B1(new_n756), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G13), .A2(G33), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G20), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n214), .B1(G20), .B2(new_n364), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n750), .B1(new_n760), .B2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n764), .ZN(new_n768));
  NAND2_X1  g0568(.A1(G20), .A2(G179), .ZN(new_n769));
  XOR2_X1   g0569(.A(new_n769), .B(KEYINPUT101), .Z(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G190), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n319), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(G200), .ZN(new_n773));
  AOI22_X1  g0573(.A1(G50), .A2(new_n772), .B1(new_n773), .B2(G58), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n770), .A2(new_n419), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n319), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(G200), .ZN(new_n777));
  AOI22_X1  g0577(.A1(G68), .A2(new_n776), .B1(new_n777), .B2(G77), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n215), .A2(G179), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n779), .A2(new_n419), .A3(new_n319), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n380), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT32), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n419), .A2(G179), .A3(G200), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n215), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n779), .A2(G190), .A3(G200), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n785), .A2(G97), .B1(new_n787), .B2(G87), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n779), .A2(new_n419), .A3(G200), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G107), .ZN(new_n791));
  AND3_X1   g0591(.A1(new_n788), .A2(new_n253), .A3(new_n791), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n774), .A2(new_n778), .A3(new_n782), .A4(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(KEYINPUT33), .B(G317), .ZN(new_n794));
  AOI22_X1  g0594(.A1(G322), .A2(new_n773), .B1(new_n776), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n777), .A2(G311), .ZN(new_n796));
  INV_X1    g0596(.A(G294), .ZN(new_n797));
  INV_X1    g0597(.A(G283), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n784), .A2(new_n797), .B1(new_n789), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n780), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n253), .B(new_n799), .C1(G329), .C2(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n786), .B(KEYINPUT102), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n772), .A2(G326), .B1(G303), .B2(new_n802), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n795), .A2(new_n796), .A3(new_n801), .A4(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n768), .B1(new_n793), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n767), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n763), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n806), .B1(new_n699), .B2(new_n807), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n752), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(G396));
  AND2_X1   g0610(.A1(new_n688), .A2(new_n361), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n639), .A2(new_n641), .A3(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT106), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n812), .B(new_n813), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n367), .B(KEYINPUT105), .ZN(new_n815));
  INV_X1    g0615(.A(new_n811), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n815), .A2(new_n363), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n715), .B(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n750), .B1(new_n819), .B2(new_n742), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(new_n742), .B2(new_n819), .ZN(new_n821));
  AOI22_X1  g0621(.A1(G143), .A2(new_n773), .B1(new_n777), .B2(G159), .ZN(new_n822));
  INV_X1    g0622(.A(G137), .ZN(new_n823));
  INV_X1    g0623(.A(new_n772), .ZN(new_n824));
  INV_X1    g0624(.A(G150), .ZN(new_n825));
  INV_X1    g0625(.A(new_n776), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n822), .B1(new_n823), .B2(new_n824), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT34), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n827), .A2(new_n828), .ZN(new_n830));
  INV_X1    g0630(.A(new_n802), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n831), .A2(new_n202), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n388), .B1(new_n800), .B2(G132), .ZN(new_n833));
  INV_X1    g0633(.A(G58), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n833), .B1(new_n834), .B2(new_n784), .C1(new_n328), .C2(new_n789), .ZN(new_n835));
  NOR4_X1   g0635(.A1(new_n829), .A2(new_n830), .A3(new_n832), .A4(new_n835), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n798), .A2(new_n826), .B1(new_n824), .B2(new_n502), .ZN(new_n837));
  INV_X1    g0637(.A(new_n777), .ZN(new_n838));
  INV_X1    g0638(.A(new_n773), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n458), .A2(new_n838), .B1(new_n839), .B2(new_n797), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n253), .B1(G311), .B2(new_n800), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n785), .A2(G97), .B1(new_n790), .B2(G87), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n841), .B(new_n842), .C1(new_n831), .C2(new_n221), .ZN(new_n843));
  NOR3_X1   g0643(.A1(new_n837), .A2(new_n840), .A3(new_n843), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT104), .Z(new_n845));
  OAI21_X1  g0645(.A(new_n764), .B1(new_n836), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n764), .A2(new_n761), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT103), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n751), .B1(new_n849), .B2(new_n219), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n846), .B(new_n850), .C1(new_n818), .C2(new_n762), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n821), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(G384));
  NAND4_X1  g0653(.A1(new_n442), .A2(new_n423), .A3(new_n431), .A4(new_n438), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n682), .B1(new_n408), .B2(new_n410), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n441), .A2(new_n855), .A3(new_n429), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(KEYINPUT37), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT37), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n441), .A2(new_n855), .A3(new_n429), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT38), .B1(new_n857), .B2(new_n862), .ZN(new_n863));
  NOR4_X1   g0663(.A1(new_n408), .A2(new_n410), .A3(new_n420), .A4(new_n421), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n392), .A2(new_n281), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n383), .A2(new_n391), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n865), .B1(KEYINPUT16), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n436), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n867), .A2(new_n424), .B1(new_n868), .B2(new_n681), .ZN(new_n869));
  OAI21_X1  g0669(.A(KEYINPUT37), .B1(new_n864), .B2(new_n869), .ZN(new_n870));
  AND2_X1   g0670(.A1(new_n870), .A2(new_n861), .ZN(new_n871));
  INV_X1    g0671(.A(new_n432), .ZN(new_n872));
  AND3_X1   g0672(.A1(new_n442), .A2(new_n443), .A3(new_n438), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n443), .B1(new_n442), .B2(new_n438), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n867), .A2(new_n424), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n682), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n871), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n863), .B1(new_n879), .B2(KEYINPUT38), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT110), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n727), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(new_n733), .B2(new_n688), .ZN(new_n883));
  INV_X1    g0683(.A(new_n734), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n735), .B1(new_n881), .B2(KEYINPUT96), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n717), .ZN(new_n887));
  AND2_X1   g0687(.A1(new_n688), .A2(new_n337), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n371), .A2(new_n372), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n888), .B1(new_n340), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n373), .A2(KEYINPUT108), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT108), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n892), .B(new_n337), .C1(new_n371), .C2(new_n372), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n888), .B1(new_n325), .B2(new_n338), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n891), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n890), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n887), .A2(KEYINPUT40), .A3(new_n818), .A4(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT111), .B1(new_n880), .B2(new_n897), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n887), .A2(new_n818), .A3(new_n896), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n870), .A2(new_n861), .ZN(new_n900));
  OAI211_X1 g0700(.A(KEYINPUT38), .B(new_n900), .C1(new_n445), .C2(new_n877), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n857), .A2(new_n862), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT38), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT111), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n899), .A2(new_n905), .A3(new_n906), .A4(KEYINPUT40), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n898), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n875), .A2(new_n878), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT38), .B1(new_n909), .B2(new_n900), .ZN(new_n910));
  AOI211_X1 g0710(.A(new_n903), .B(new_n871), .C1(new_n875), .C2(new_n878), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n899), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT40), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n908), .A2(new_n914), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n915), .B(KEYINPUT112), .Z(new_n916));
  NAND2_X1  g0716(.A1(new_n447), .A2(new_n887), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(new_n917), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n918), .A2(G330), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(KEYINPUT39), .B1(new_n910), .B2(new_n911), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT39), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n901), .A2(new_n904), .A3(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n921), .A2(KEYINPUT109), .A3(new_n923), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n891), .A2(new_n893), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n925), .A2(new_n688), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n900), .B1(new_n445), .B2(new_n877), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n903), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n901), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT109), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n929), .A2(new_n930), .A3(KEYINPUT39), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n924), .A2(new_n926), .A3(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n636), .A2(new_n682), .ZN(new_n933));
  INV_X1    g0733(.A(new_n896), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n673), .A2(new_n692), .A3(new_n818), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n815), .A2(new_n688), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n933), .B1(new_n937), .B2(new_n929), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n932), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n447), .B(new_n714), .C1(new_n715), .C2(KEYINPUT29), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n645), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n939), .B(new_n941), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n920), .A2(new_n942), .B1(new_n267), .B2(new_n747), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n943), .A2(KEYINPUT113), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n920), .A2(new_n942), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n943), .A2(KEYINPUT113), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n376), .A2(G77), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n212), .A2(new_n948), .B1(G50), .B2(new_n328), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n949), .A2(G1), .A3(new_n290), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT107), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n216), .A2(G116), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(new_n544), .B2(KEYINPUT35), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(KEYINPUT35), .B2(new_n544), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT36), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n951), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(new_n955), .B2(new_n954), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n947), .A2(new_n957), .ZN(G367));
  NAND2_X1  g0758(.A1(new_n576), .A2(new_n490), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n688), .B1(new_n959), .B2(new_n577), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n573), .B1(new_n550), .B2(new_n692), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n577), .B2(new_n692), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n691), .A2(new_n694), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n960), .B1(new_n963), .B2(KEYINPUT42), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(KEYINPUT42), .B2(new_n963), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT43), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n626), .A2(new_n594), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n688), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n669), .B(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n965), .B1(new_n966), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n966), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n970), .B(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n696), .A2(new_n700), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n962), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n972), .B(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n695), .A2(new_n962), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT45), .Z(new_n977));
  NOR2_X1   g0777(.A1(new_n695), .A2(new_n962), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT44), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(new_n973), .ZN(new_n981));
  MUX2_X1   g0781(.A(new_n691), .B(new_n696), .S(new_n693), .Z(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(new_n700), .Z(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n743), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n743), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n703), .B(KEYINPUT41), .Z(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n975), .B1(new_n988), .B2(new_n749), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n784), .A2(new_n328), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(G137), .B2(new_n800), .ZN(new_n991));
  INV_X1    g0791(.A(G143), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n991), .B1(new_n834), .B2(new_n786), .C1(new_n824), .C2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n253), .B1(new_n219), .B2(new_n789), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT114), .Z(new_n995));
  NOR2_X1   g0795(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  AOI22_X1  g0796(.A1(G50), .A2(new_n777), .B1(new_n773), .B2(G150), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n996), .B(new_n997), .C1(new_n380), .C2(new_n826), .ZN(new_n998));
  AOI21_X1  g0798(.A(KEYINPUT46), .B1(new_n787), .B2(G116), .ZN(new_n999));
  INV_X1    g0799(.A(G317), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n388), .B1(new_n780), .B2(new_n1000), .C1(new_n517), .C2(new_n789), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n999), .B(new_n1001), .C1(G107), .C2(new_n785), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n802), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(G283), .A2(new_n777), .B1(new_n773), .B2(G303), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(G294), .A2(new_n776), .B1(new_n772), .B2(G311), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n998), .A2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT47), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n764), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n969), .A2(new_n763), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n765), .B1(new_n208), .B2(new_n355), .C1(new_n236), .C2(new_n758), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1009), .A2(new_n750), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n989), .A2(new_n1012), .ZN(G387));
  OAI22_X1  g0813(.A1(new_n202), .A2(new_n839), .B1(new_n824), .B2(new_n380), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(new_n284), .B2(new_n776), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n786), .A2(new_n219), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n386), .B1(new_n780), .B2(new_n825), .C1(new_n517), .C2(new_n789), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n1016), .B(new_n1017), .C1(new_n356), .C2(new_n785), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1015), .B(new_n1018), .C1(new_n328), .C2(new_n838), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n386), .B1(new_n800), .B2(G326), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n784), .A2(new_n798), .B1(new_n786), .B2(new_n797), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G311), .A2(new_n776), .B1(new_n772), .B2(G322), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1022), .B1(new_n502), .B2(new_n838), .C1(new_n1000), .C2(new_n839), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT48), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1021), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n1024), .B2(new_n1023), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT49), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1020), .B1(new_n458), .B2(new_n789), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  AND2_X1   g0828(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1019), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n764), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n757), .B1(new_n233), .B2(new_n464), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n706), .B2(new_n753), .ZN(new_n1033));
  OR3_X1    g0833(.A1(new_n283), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1034));
  OAI21_X1  g0834(.A(KEYINPUT50), .B1(new_n283), .B2(G50), .ZN(new_n1035));
  AOI21_X1  g0835(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1034), .A2(new_n706), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n1033), .A2(new_n1037), .B1(new_n221), .B2(new_n702), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1031), .B(new_n750), .C1(new_n766), .C2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(new_n696), .B2(new_n763), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT115), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n983), .B2(new_n749), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n984), .A2(new_n703), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n983), .A2(new_n743), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1042), .B1(new_n1043), .B2(new_n1044), .ZN(G393));
  OR2_X1    g0845(.A1(new_n981), .A2(new_n748), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n766), .B1(G97), .B2(new_n702), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n240), .A2(new_n757), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n751), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G150), .A2(new_n772), .B1(new_n773), .B2(G159), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT51), .Z(new_n1051));
  OAI22_X1  g0851(.A1(new_n784), .A2(new_n219), .B1(new_n786), .B2(new_n328), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n386), .B1(new_n780), .B2(new_n992), .C1(new_n414), .C2(new_n789), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n1052), .B(new_n1053), .C1(new_n776), .C2(G50), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1051), .B(new_n1054), .C1(new_n283), .C2(new_n838), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(G311), .A2(new_n773), .B1(new_n772), .B2(G317), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT52), .Z(new_n1057));
  OAI221_X1 g0857(.A(new_n791), .B1(new_n798), .B2(new_n786), .C1(new_n458), .C2(new_n784), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n253), .B(new_n1058), .C1(G322), .C2(new_n800), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(G294), .A2(new_n777), .B1(new_n776), .B2(G303), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1057), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n1055), .A2(new_n1061), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1049), .B1(new_n768), .B2(new_n1062), .C1(new_n962), .C2(new_n807), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n981), .A2(new_n984), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n703), .B1(new_n981), .B2(new_n984), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1046), .B(new_n1063), .C1(new_n1065), .C2(new_n1066), .ZN(G390));
  INV_X1    g0867(.A(G330), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n886), .B2(new_n717), .ZN(new_n1069));
  AND3_X1   g0869(.A1(new_n1069), .A2(new_n818), .A3(new_n896), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n935), .A2(new_n936), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n926), .B1(new_n1071), .B2(new_n896), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(new_n924), .B2(new_n931), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n818), .B(new_n692), .C1(new_n711), .C2(new_n713), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n936), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n896), .ZN(new_n1076));
  OR3_X1    g0876(.A1(new_n925), .A2(KEYINPUT116), .A3(new_n688), .ZN(new_n1077));
  OAI21_X1  g0877(.A(KEYINPUT116), .B1(new_n925), .B2(new_n688), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1076), .A2(new_n1077), .A3(new_n905), .A4(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1070), .B1(new_n1073), .B2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n741), .A2(new_n818), .A3(new_n896), .ZN(new_n1082));
  AOI211_X1 g0882(.A(KEYINPUT109), .B(new_n922), .C1(new_n928), .C2(new_n901), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n930), .B1(new_n929), .B2(KEYINPUT39), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1083), .B1(new_n1084), .B2(new_n923), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1079), .B(new_n1082), .C1(new_n1085), .C2(new_n1072), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n447), .A2(new_n1069), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n940), .A2(new_n645), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n896), .B1(new_n741), .B2(new_n818), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1071), .B1(new_n1089), .B2(new_n1070), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT117), .ZN(new_n1091));
  AND2_X1   g0891(.A1(new_n1069), .A2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n818), .B1(new_n1069), .B2(new_n1091), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n934), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1094), .A2(new_n1082), .A3(new_n936), .A4(new_n1074), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1088), .B1(new_n1090), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1081), .A2(new_n1086), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1096), .B1(new_n1081), .B2(new_n1086), .ZN(new_n1099));
  NOR3_X1   g0899(.A1(new_n1098), .A2(new_n1099), .A3(new_n704), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1081), .A2(new_n1086), .A3(new_n749), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n750), .B1(new_n848), .B2(new_n284), .ZN(new_n1103));
  XOR2_X1   g0903(.A(KEYINPUT54), .B(G143), .Z(new_n1104));
  AOI22_X1  g0904(.A1(G137), .A2(new_n776), .B1(new_n777), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n773), .A2(G132), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n785), .A2(G159), .B1(new_n790), .B2(G50), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n800), .A2(G125), .ZN(new_n1108));
  AND3_X1   g0908(.A1(new_n1107), .A2(new_n253), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT53), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n786), .B2(new_n825), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n787), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n772), .A2(G128), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1105), .A2(new_n1106), .A3(new_n1109), .A4(new_n1113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(G107), .A2(new_n776), .B1(new_n772), .B2(G283), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n517), .B2(new_n838), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT118), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n253), .B1(G294), .B2(new_n800), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n785), .A2(G77), .B1(new_n790), .B2(G68), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1120), .B1(new_n414), .B2(new_n831), .C1(new_n458), .C2(new_n839), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1114), .B1(new_n1117), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1103), .B1(new_n1122), .B2(new_n764), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n1085), .B2(new_n762), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1102), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1101), .A2(new_n1126), .ZN(G378));
  NAND3_X1  g0927(.A1(new_n908), .A2(G330), .A3(new_n914), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n939), .A2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n297), .A2(new_n681), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n635), .A2(new_n343), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(KEYINPUT119), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT119), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n635), .A2(new_n1135), .A3(new_n343), .ZN(new_n1136));
  XOR2_X1   g0936(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n1134), .A2(new_n1136), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1138), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1132), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n1137), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1134), .A2(new_n1136), .A3(new_n1138), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1143), .A2(new_n1131), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(KEYINPUT120), .B1(new_n1141), .B2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1128), .A2(new_n932), .A3(new_n938), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1130), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1146), .B1(new_n1130), .B2(new_n1147), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n749), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1141), .A2(new_n1145), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n761), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n751), .B1(new_n849), .B2(new_n202), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(G125), .A2(new_n772), .B1(new_n773), .B2(G128), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(new_n823), .B2(new_n838), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n785), .A2(G150), .B1(new_n787), .B2(new_n1104), .ZN(new_n1156));
  INV_X1    g0956(.A(G132), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1156), .B1(new_n826), .B2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  OR2_X1    g0960(.A1(new_n1160), .A2(KEYINPUT59), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(KEYINPUT59), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n790), .A2(G159), .ZN(new_n1163));
  AOI211_X1 g0963(.A(G33), .B(G41), .C1(new_n800), .C2(G124), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(G41), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1166), .B(new_n388), .C1(new_n780), .C2(new_n798), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n789), .A2(new_n834), .ZN(new_n1168));
  OR4_X1    g0968(.A1(new_n990), .A2(new_n1167), .A3(new_n1016), .A4(new_n1168), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(G97), .A2(new_n776), .B1(new_n773), .B2(G107), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n458), .B2(new_n824), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1169), .B(new_n1171), .C1(new_n356), .C2(new_n777), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(KEYINPUT58), .ZN(new_n1173));
  AOI21_X1  g0973(.A(G50), .B1(new_n249), .B2(new_n1166), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n386), .B2(G41), .ZN(new_n1175));
  OR2_X1    g0975(.A1(new_n1172), .A2(KEYINPUT58), .ZN(new_n1176));
  AND4_X1   g0976(.A1(new_n1165), .A2(new_n1173), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1152), .B(new_n1153), .C1(new_n768), .C2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1150), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1088), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1097), .A2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT57), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n1183), .A2(KEYINPUT121), .A3(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT121), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT120), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1151), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1147), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1128), .B1(new_n932), .B2(new_n938), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1188), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1130), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1191), .A2(new_n1192), .B1(new_n1181), .B2(new_n1097), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1186), .B1(new_n1193), .B2(KEYINPUT57), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1185), .A2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(KEYINPUT122), .B1(new_n1193), .B2(KEYINPUT57), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT122), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1183), .A2(new_n1197), .A3(new_n1184), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1196), .A2(new_n1198), .A3(new_n703), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1180), .B1(new_n1195), .B2(new_n1199), .ZN(G375));
  INV_X1    g1000(.A(new_n1096), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1090), .A2(new_n1095), .A3(new_n1088), .ZN(new_n1202));
  XOR2_X1   g1002(.A(new_n986), .B(KEYINPUT123), .Z(new_n1203));
  NAND3_X1  g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n748), .B1(new_n1090), .B2(new_n1095), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n934), .A2(new_n761), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n750), .B1(new_n848), .B2(G68), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n776), .A2(G116), .B1(G97), .B2(new_n802), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1208), .B1(new_n798), .B2(new_n839), .C1(new_n797), .C2(new_n824), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n253), .B1(G303), .B2(new_n800), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n785), .A2(new_n356), .B1(new_n790), .B2(G77), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1210), .B(new_n1211), .C1(new_n838), .C2(new_n221), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT124), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n824), .B2(new_n1157), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n772), .A2(KEYINPUT124), .A3(G132), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n777), .A2(G150), .ZN(new_n1216));
  INV_X1    g1016(.A(G128), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n386), .B1(new_n780), .B2(new_n1217), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1168), .B(new_n1218), .C1(G50), .C2(new_n785), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .A4(new_n1219), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(G137), .A2(new_n773), .B1(new_n776), .B2(new_n1104), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n380), .B2(new_n831), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n1209), .A2(new_n1212), .B1(new_n1220), .B2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1207), .B1(new_n1223), .B2(new_n764), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1205), .B1(new_n1206), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1204), .A2(new_n1225), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1226), .B(KEYINPUT125), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(G381));
  INV_X1    g1028(.A(G375), .ZN(new_n1229));
  OR3_X1    g1029(.A1(new_n1100), .A2(KEYINPUT126), .A3(new_n1125), .ZN(new_n1230));
  OAI21_X1  g1030(.A(KEYINPUT126), .B1(new_n1100), .B2(new_n1125), .ZN(new_n1231));
  AND2_X1   g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1229), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(G387), .ZN(new_n1235));
  NOR4_X1   g1035(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1234), .A2(new_n1235), .A3(new_n1227), .A4(new_n1236), .ZN(G407));
  NAND2_X1  g1037(.A1(new_n683), .A2(G213), .ZN(new_n1238));
  OAI211_X1 g1038(.A(G407), .B(G213), .C1(new_n1233), .C2(new_n1238), .ZN(G409));
  OAI211_X1 g1039(.A(G378), .B(new_n1180), .C1(new_n1195), .C2(new_n1199), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1193), .A2(new_n1203), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1230), .B(new_n1231), .C1(new_n1179), .C2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1240), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1238), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1238), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(G2897), .ZN(new_n1246));
  XOR2_X1   g1046(.A(new_n1246), .B(KEYINPUT127), .Z(new_n1247));
  AND2_X1   g1047(.A1(new_n1201), .A2(KEYINPUT60), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1202), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n704), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(new_n1249), .B2(new_n1248), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1251), .A2(G384), .A3(new_n1225), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(G384), .B1(new_n1251), .B2(new_n1225), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1247), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1254), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1247), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1256), .A2(new_n1252), .A3(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1255), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT61), .B1(new_n1244), .B2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT63), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1262), .B1(new_n1244), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1235), .A2(G390), .ZN(new_n1266));
  INV_X1    g1066(.A(G390), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(G387), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(G393), .B(new_n809), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(new_n1269), .B(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1245), .B1(new_n1240), .B2(new_n1242), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1272), .A2(KEYINPUT63), .A3(new_n1263), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1261), .A2(new_n1265), .A3(new_n1271), .A4(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT62), .ZN(new_n1275));
  AND3_X1   g1075(.A1(new_n1272), .A2(new_n1275), .A3(new_n1263), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT61), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1277), .B1(new_n1272), .B2(new_n1259), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1275), .B1(new_n1272), .B2(new_n1263), .ZN(new_n1279));
  NOR3_X1   g1079(.A1(new_n1276), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1274), .B1(new_n1280), .B2(new_n1271), .ZN(G405));
  NAND2_X1  g1081(.A1(G375), .A2(new_n1232), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1282), .A2(new_n1264), .A3(new_n1240), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1264), .B1(new_n1282), .B2(new_n1240), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(new_n1286), .B(new_n1271), .ZN(G402));
endmodule


