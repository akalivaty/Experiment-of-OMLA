//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 0 0 1 0 1 0 0 1 0 0 1 0 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 0 0 0 0 0 0 1 0 1 1 0 1 1 1 0 1 1 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT68), .ZN(new_n188));
  INV_X1    g002(.A(G116), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(G119), .ZN(new_n191));
  INV_X1    g005(.A(G119), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT68), .A3(G116), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n191), .A3(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G113), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT2), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT2), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G113), .ZN(new_n198));
  AND2_X1   g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n194), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n196), .A2(new_n198), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n201), .A2(new_n191), .A3(new_n193), .A4(new_n190), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G134), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(G137), .ZN(new_n205));
  INV_X1    g019(.A(G137), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(G134), .ZN(new_n207));
  OAI21_X1  g021(.A(G131), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT11), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n209), .B1(new_n204), .B2(G137), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n211), .B1(new_n206), .B2(G134), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n206), .A2(KEYINPUT11), .A3(G134), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n204), .A2(KEYINPUT66), .A3(G137), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n210), .A2(new_n212), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n208), .B1(new_n215), .B2(G131), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT67), .ZN(new_n217));
  INV_X1    g031(.A(G143), .ZN(new_n218));
  INV_X1    g032(.A(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT64), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT64), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G146), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n218), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT1), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n217), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT64), .B(G146), .ZN(new_n226));
  OAI211_X1 g040(.A(KEYINPUT67), .B(KEYINPUT1), .C1(new_n226), .C2(new_n218), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n225), .A2(G128), .A3(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n218), .A2(G146), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n220), .A2(new_n222), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(G143), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n228), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT65), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n223), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT65), .B1(new_n226), .B2(new_n218), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n219), .A2(G143), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G128), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(KEYINPUT1), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n235), .A2(new_n236), .A3(new_n238), .A4(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n216), .B1(new_n233), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(KEYINPUT0), .A2(G128), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n235), .A2(new_n236), .A3(new_n244), .A4(new_n238), .ZN(new_n245));
  OR2_X1    g059(.A1(KEYINPUT0), .A2(G128), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n232), .A2(new_n243), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G131), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n215), .B(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n203), .B1(new_n242), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n203), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n215), .B(G131), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(new_n245), .A3(new_n247), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n238), .B1(new_n223), .B2(new_n234), .ZN(new_n256));
  NOR3_X1   g070(.A1(new_n226), .A2(KEYINPUT65), .A3(new_n218), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n232), .A2(new_n228), .B1(new_n258), .B2(new_n240), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n253), .B(new_n255), .C1(new_n259), .C2(new_n216), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n252), .A2(KEYINPUT70), .A3(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n262));
  OAI211_X1 g076(.A(new_n262), .B(new_n203), .C1(new_n242), .C2(new_n251), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n261), .A2(KEYINPUT28), .A3(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n265), .B(G101), .ZN(new_n266));
  INV_X1    g080(.A(G237), .ZN(new_n267));
  INV_X1    g081(.A(G953), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n267), .A2(new_n268), .A3(G210), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n266), .B(new_n269), .ZN(new_n270));
  NOR3_X1   g084(.A1(new_n242), .A2(new_n251), .A3(new_n203), .ZN(new_n271));
  OR2_X1    g085(.A1(new_n271), .A2(KEYINPUT28), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n264), .A2(KEYINPUT29), .A3(new_n270), .A4(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G902), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT29), .ZN(new_n276));
  INV_X1    g090(.A(new_n270), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT30), .B1(new_n242), .B2(new_n251), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT30), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n279), .B(new_n255), .C1(new_n259), .C2(new_n216), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n253), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n277), .B1(new_n281), .B2(new_n271), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT69), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n252), .A2(new_n283), .A3(new_n260), .ZN(new_n284));
  OAI211_X1 g098(.A(KEYINPUT69), .B(new_n203), .C1(new_n242), .C2(new_n251), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n284), .A2(KEYINPUT28), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n272), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n276), .B(new_n282), .C1(new_n287), .C2(new_n277), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n187), .B1(new_n275), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n270), .B1(new_n286), .B2(new_n272), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT31), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n278), .A2(new_n280), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n271), .B1(new_n292), .B2(new_n203), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n291), .B1(new_n293), .B2(new_n270), .ZN(new_n294));
  NOR4_X1   g108(.A1(new_n281), .A2(KEYINPUT31), .A3(new_n277), .A4(new_n271), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n290), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(G472), .A2(G902), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(KEYINPUT32), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n287), .A2(new_n277), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n292), .A2(new_n203), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n301), .A2(new_n270), .A3(new_n260), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT31), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n293), .A2(new_n291), .A3(new_n270), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n300), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT32), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(new_n306), .A3(new_n297), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n289), .B1(new_n299), .B2(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(G125), .B(G140), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT16), .ZN(new_n310));
  INV_X1    g124(.A(G125), .ZN(new_n311));
  OR3_X1    g125(.A1(new_n311), .A2(KEYINPUT16), .A3(G140), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n219), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n310), .A2(G146), .A3(new_n312), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  XOR2_X1   g130(.A(KEYINPUT24), .B(G110), .Z(new_n317));
  XNOR2_X1  g131(.A(G119), .B(G128), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n192), .A2(G128), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT23), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT23), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n322), .B1(new_n192), .B2(G128), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n321), .B(new_n323), .C1(G119), .C2(new_n239), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n324), .B(KEYINPUT71), .ZN(new_n325));
  INV_X1    g139(.A(G110), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n316), .B(new_n319), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n309), .B(KEYINPUT72), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n231), .ZN(new_n329));
  OAI22_X1  g143(.A1(new_n324), .A2(G110), .B1(new_n318), .B2(new_n317), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(new_n330), .A3(new_n315), .ZN(new_n331));
  AND2_X1   g145(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n268), .A2(G221), .A3(G234), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n333), .B(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(KEYINPUT22), .B(G137), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n335), .B(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n332), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n337), .B(KEYINPUT75), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n338), .B(new_n274), .C1(new_n332), .C2(new_n339), .ZN(new_n340));
  XOR2_X1   g154(.A(KEYINPUT76), .B(KEYINPUT25), .Z(new_n341));
  OR2_X1    g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G234), .ZN(new_n343));
  OAI21_X1  g157(.A(G217), .B1(new_n343), .B2(G902), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT25), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n345), .A2(KEYINPUT76), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n344), .B1(new_n340), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n342), .A2(new_n347), .ZN(new_n348));
  OR2_X1    g162(.A1(new_n332), .A2(new_n339), .ZN(new_n349));
  AOI21_X1  g163(.A(G902), .B1(new_n343), .B2(G217), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(new_n338), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n308), .A2(new_n352), .ZN(new_n353));
  XOR2_X1   g167(.A(KEYINPUT9), .B(G234), .Z(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(G221), .B1(new_n355), .B2(G902), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(G214), .B1(G237), .B2(G902), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n190), .A2(new_n193), .A3(KEYINPUT5), .A4(new_n191), .ZN(new_n359));
  NOR3_X1   g173(.A1(new_n189), .A2(KEYINPUT5), .A3(G119), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n360), .A2(new_n195), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(KEYINPUT84), .ZN(new_n363));
  XNOR2_X1  g177(.A(KEYINPUT78), .B(G101), .ZN(new_n364));
  INV_X1    g178(.A(G104), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G107), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT3), .ZN(new_n367));
  INV_X1    g181(.A(G107), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(new_n368), .A3(G104), .ZN(new_n369));
  OAI21_X1  g183(.A(KEYINPUT3), .B1(new_n365), .B2(G107), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n364), .A2(new_n366), .A3(new_n369), .A4(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n368), .A2(G104), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n366), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G101), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT84), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n359), .A2(new_n361), .A3(new_n376), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n363), .A2(new_n202), .A3(new_n375), .A4(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n375), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n362), .A2(new_n202), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(G110), .B(G122), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n382), .B(KEYINPUT8), .ZN(new_n383));
  AND3_X1   g197(.A1(new_n378), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n233), .A2(new_n311), .A3(new_n241), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n248), .A2(G125), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G224), .ZN(new_n388));
  OAI21_X1  g202(.A(KEYINPUT7), .B1(new_n388), .B2(G953), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n384), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n389), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n385), .A2(new_n386), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT87), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n370), .A2(new_n369), .A3(new_n366), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G101), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(KEYINPUT4), .A3(new_n371), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT4), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n395), .A2(new_n398), .A3(G101), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n397), .A2(new_n203), .A3(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT83), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n379), .A2(new_n363), .A3(new_n202), .A4(new_n377), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n397), .A2(KEYINPUT83), .A3(new_n203), .A4(new_n399), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n402), .A2(new_n382), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n385), .A2(KEYINPUT87), .A3(new_n386), .A4(new_n391), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n390), .A2(new_n394), .A3(new_n405), .A4(new_n406), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n407), .A2(new_n274), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT6), .ZN(new_n410));
  INV_X1    g224(.A(new_n382), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT85), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n409), .A2(KEYINPUT85), .A3(new_n410), .A4(new_n411), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n388), .A2(G953), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n417), .B(KEYINPUT86), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n387), .B(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n409), .A2(new_n411), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n420), .A2(KEYINPUT6), .A3(new_n405), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n416), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(G210), .B1(G237), .B2(G902), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n408), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n423), .B1(new_n408), .B2(new_n422), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n358), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n268), .A2(G227), .ZN(new_n427));
  XOR2_X1   g241(.A(new_n427), .B(G140), .Z(new_n428));
  XNOR2_X1  g242(.A(new_n428), .B(KEYINPUT77), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n429), .B(new_n326), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n239), .B1(new_n230), .B2(KEYINPUT1), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n433), .B1(new_n256), .B2(new_n257), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n375), .B1(new_n434), .B2(new_n241), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n435), .B1(new_n259), .B2(new_n375), .ZN(new_n436));
  OAI21_X1  g250(.A(KEYINPUT12), .B1(new_n436), .B2(new_n250), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n233), .A2(new_n241), .A3(new_n375), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n221), .A2(G146), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n219), .A2(KEYINPUT64), .ZN(new_n440));
  OAI21_X1  g254(.A(G143), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n237), .B1(new_n441), .B2(KEYINPUT65), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n432), .B1(new_n442), .B2(new_n235), .ZN(new_n443));
  AND4_X1   g257(.A1(new_n235), .A2(new_n236), .A3(new_n238), .A4(new_n240), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n379), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n438), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT12), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(new_n447), .A3(new_n254), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT79), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT10), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n445), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(KEYINPUT79), .B1(new_n435), .B2(KEYINPUT10), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n397), .A2(new_n399), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n248), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n232), .ZN(new_n456));
  OAI21_X1  g270(.A(KEYINPUT1), .B1(new_n226), .B2(new_n218), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n239), .B1(new_n457), .B2(new_n217), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n456), .B1(new_n458), .B2(new_n227), .ZN(new_n459));
  OAI211_X1 g273(.A(KEYINPUT10), .B(new_n379), .C1(new_n459), .C2(new_n444), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n451), .A2(new_n452), .A3(new_n455), .A4(new_n460), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n437), .B(new_n448), .C1(new_n461), .C2(new_n254), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT80), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n447), .B1(new_n446), .B2(new_n254), .ZN(new_n465));
  AOI211_X1 g279(.A(KEYINPUT12), .B(new_n250), .C1(new_n438), .C2(new_n445), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n375), .B1(new_n233), .B2(new_n241), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n454), .B1(new_n468), .B2(KEYINPUT10), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n469), .A2(new_n250), .A3(new_n452), .A4(new_n451), .ZN(new_n470));
  AOI21_X1  g284(.A(KEYINPUT80), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n431), .B1(new_n464), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n461), .A2(new_n254), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n431), .B1(new_n473), .B2(new_n470), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n472), .A2(new_n274), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(G469), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n473), .A2(new_n470), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n431), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT82), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n470), .A2(new_n430), .A3(new_n437), .A4(new_n448), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  OR2_X1    g296(.A1(new_n481), .A2(new_n480), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT81), .B(G469), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n482), .A2(new_n274), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  AOI211_X1 g299(.A(new_n357), .B(new_n426), .C1(new_n477), .C2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(G475), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n267), .A2(new_n268), .A3(G214), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT89), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n488), .B(KEYINPUT90), .C1(new_n489), .C2(G143), .ZN(new_n490));
  OAI21_X1  g304(.A(KEYINPUT90), .B1(new_n489), .B2(G143), .ZN(new_n491));
  OR2_X1    g305(.A1(KEYINPUT90), .A2(G143), .ZN(new_n492));
  NOR2_X1   g306(.A1(G237), .A2(G953), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n491), .A2(G214), .A3(new_n492), .A4(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n490), .A2(new_n494), .A3(G131), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT91), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n490), .A2(new_n494), .A3(KEYINPUT91), .A4(G131), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n497), .A2(KEYINPUT17), .A3(new_n498), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n314), .A2(new_n315), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT92), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(G131), .B1(new_n490), .B2(new_n494), .ZN(new_n504));
  AOI211_X1 g318(.A(KEYINPUT17), .B(new_n504), .C1(new_n497), .C2(new_n498), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n499), .A2(new_n500), .A3(KEYINPUT92), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n503), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n329), .B1(new_n219), .B2(new_n309), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n490), .A2(new_n494), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT18), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OR2_X1    g326(.A1(new_n495), .A2(new_n511), .ZN(new_n513));
  INV_X1    g327(.A(new_n504), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n509), .A2(new_n512), .A3(new_n513), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n508), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(G113), .B(G122), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(new_n365), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n518), .A2(KEYINPUT93), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(G902), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n508), .A2(new_n515), .A3(new_n519), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n487), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n499), .A2(new_n500), .A3(KEYINPUT92), .ZN(new_n524));
  AOI21_X1  g338(.A(KEYINPUT92), .B1(new_n499), .B2(new_n500), .ZN(new_n525));
  NOR3_X1   g339(.A1(new_n524), .A2(new_n525), .A3(new_n505), .ZN(new_n526));
  INV_X1    g340(.A(new_n515), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n518), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n518), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT19), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n309), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n531), .B1(new_n328), .B2(new_n530), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n231), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n315), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n504), .B1(new_n497), .B2(new_n498), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n515), .B(new_n529), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n528), .A2(new_n487), .A3(new_n274), .A4(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT88), .B(KEYINPUT20), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n536), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n540), .B1(new_n516), .B2(new_n518), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT20), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n541), .A2(new_n542), .A3(new_n487), .A4(new_n274), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n523), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(G478), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n546), .A2(KEYINPUT15), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n354), .A2(G217), .A3(new_n268), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n239), .A2(G143), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n218), .A2(G128), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n550), .A2(new_n551), .A3(new_n204), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT13), .ZN(new_n553));
  OAI21_X1  g367(.A(KEYINPUT95), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n551), .A2(new_n553), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT95), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n556), .A2(new_n218), .A3(KEYINPUT13), .A4(G128), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n554), .A2(new_n550), .A3(new_n555), .A4(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n552), .B1(new_n558), .B2(G134), .ZN(new_n559));
  INV_X1    g373(.A(G122), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(G116), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n189), .A2(G122), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT94), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n561), .A2(new_n562), .A3(KEYINPUT94), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(G107), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n368), .B1(new_n565), .B2(new_n566), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n559), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n189), .A2(KEYINPUT14), .A3(G122), .ZN(new_n571));
  OAI211_X1 g385(.A(G107), .B(new_n571), .C1(new_n563), .C2(KEYINPUT14), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n204), .B1(new_n550), .B2(new_n551), .ZN(new_n573));
  OAI221_X1 g387(.A(new_n572), .B1(new_n573), .B2(new_n552), .C1(new_n567), .C2(G107), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n570), .A2(new_n574), .A3(KEYINPUT96), .ZN(new_n575));
  AOI21_X1  g389(.A(KEYINPUT96), .B1(new_n570), .B2(new_n574), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n549), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n570), .A2(new_n574), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT96), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n548), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n581), .A2(KEYINPUT97), .A3(new_n274), .ZN(new_n582));
  AOI21_X1  g396(.A(G902), .B1(new_n577), .B2(new_n580), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n583), .A2(KEYINPUT97), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n547), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  OAI22_X1  g399(.A1(new_n583), .A2(KEYINPUT97), .B1(KEYINPUT15), .B2(new_n546), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(G952), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n588), .A2(KEYINPUT98), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n588), .A2(KEYINPUT98), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n268), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n591), .B1(G234), .B2(G237), .ZN(new_n592));
  XOR2_X1   g406(.A(KEYINPUT21), .B(G898), .Z(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  AOI211_X1 g408(.A(new_n274), .B(new_n268), .C1(G234), .C2(G237), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n592), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NOR3_X1   g410(.A1(new_n545), .A2(new_n587), .A3(new_n596), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n353), .A2(new_n486), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(new_n364), .ZN(G3));
  AOI21_X1  g413(.A(new_n357), .B1(new_n477), .B2(new_n485), .ZN(new_n600));
  INV_X1    g414(.A(new_n596), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n358), .B(new_n601), .C1(new_n424), .C2(new_n425), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n583), .A2(G478), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT33), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT99), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n578), .B1(new_n605), .B2(new_n549), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n570), .A2(new_n574), .A3(KEYINPUT99), .A4(new_n548), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n604), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AOI211_X1 g422(.A(G902), .B(new_n608), .C1(new_n581), .C2(new_n604), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n603), .B1(new_n609), .B2(G478), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n602), .A2(new_n544), .A3(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n352), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n187), .B1(new_n305), .B2(new_n274), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n294), .A2(new_n295), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n298), .B1(new_n614), .B2(new_n300), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n600), .A2(new_n611), .A3(new_n612), .A4(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT34), .B(G104), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G6));
  XNOR2_X1  g433(.A(new_n537), .B(new_n538), .ZN(new_n620));
  INV_X1    g434(.A(new_n523), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n620), .A2(new_n587), .A3(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n622), .A2(new_n602), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n600), .A2(new_n612), .A3(new_n616), .A4(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT35), .B(G107), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G9));
  INV_X1    g440(.A(KEYINPUT36), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n339), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(new_n332), .ZN(new_n629));
  AOI22_X1  g443(.A1(new_n342), .A2(new_n347), .B1(new_n350), .B2(new_n629), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n613), .A2(new_n615), .A3(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n358), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n408), .A2(new_n422), .ZN(new_n633));
  INV_X1    g447(.A(new_n423), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n408), .A2(new_n422), .A3(new_n423), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n632), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n600), .A2(new_n631), .A3(new_n597), .A4(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT37), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(new_n326), .ZN(G12));
  NAND2_X1  g454(.A1(new_n299), .A2(new_n307), .ZN(new_n641));
  INV_X1    g455(.A(new_n289), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n630), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(G900), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n592), .B1(new_n644), .B2(new_n595), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n622), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n486), .A2(new_n643), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G128), .ZN(G30));
  NOR2_X1   g462(.A1(new_n424), .A2(new_n425), .ZN(new_n649));
  XOR2_X1   g463(.A(new_n649), .B(KEYINPUT38), .Z(new_n650));
  INV_X1    g464(.A(new_n293), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n270), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n261), .A2(new_n263), .ZN(new_n653));
  OAI211_X1 g467(.A(new_n652), .B(new_n274), .C1(new_n270), .C2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(G472), .ZN(new_n655));
  AND2_X1   g469(.A1(new_n641), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n630), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n545), .A2(new_n358), .A3(new_n587), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(G469), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n462), .A2(new_n463), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n467), .A2(KEYINPUT80), .A3(new_n470), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n474), .B1(new_n663), .B2(new_n431), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n660), .B1(new_n664), .B2(new_n274), .ZN(new_n665));
  AND4_X1   g479(.A1(new_n274), .A2(new_n482), .A3(new_n483), .A4(new_n484), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n356), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n645), .B(KEYINPUT39), .ZN(new_n668));
  OR2_X1    g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT100), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n671), .A2(KEYINPUT40), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n671), .A2(KEYINPUT40), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n650), .B(new_n659), .C1(new_n672), .C2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G143), .ZN(G45));
  NOR3_X1   g489(.A1(new_n544), .A2(new_n610), .A3(new_n645), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n486), .A2(new_n643), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G146), .ZN(G48));
  NAND3_X1  g492(.A1(new_n482), .A2(new_n274), .A3(new_n483), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(G469), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n680), .A2(new_n356), .A3(new_n485), .ZN(new_n681));
  AOI211_X1 g495(.A(KEYINPUT32), .B(new_n298), .C1(new_n614), .C2(new_n300), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n306), .B1(new_n305), .B2(new_n297), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n642), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n681), .A2(new_n684), .A3(new_n611), .A4(new_n612), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT41), .B(G113), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G15));
  NAND4_X1  g501(.A1(new_n681), .A2(new_n684), .A3(new_n612), .A4(new_n623), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G116), .ZN(G18));
  NAND4_X1  g503(.A1(new_n680), .A2(new_n637), .A3(new_n356), .A4(new_n485), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n691), .A2(new_n684), .A3(new_n597), .A4(new_n657), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G119), .ZN(G21));
  NOR2_X1   g507(.A1(new_n658), .A2(new_n649), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n264), .A2(new_n272), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n277), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n298), .B1(new_n614), .B2(new_n696), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n613), .A2(new_n352), .A3(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n694), .A2(new_n681), .A3(new_n601), .A4(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(KEYINPUT101), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(new_n560), .ZN(G24));
  OAI21_X1  g515(.A(G472), .B1(new_n296), .B2(G902), .ZN(new_n702));
  INV_X1    g516(.A(new_n697), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n676), .A2(new_n702), .A3(new_n657), .A4(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n704), .A2(new_n690), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(new_n311), .ZN(G27));
  INV_X1    g520(.A(KEYINPUT42), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n635), .A2(new_n358), .A3(new_n636), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n684), .A2(new_n600), .A3(new_n612), .A4(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n676), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n707), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  AOI211_X1 g526(.A(new_n357), .B(new_n708), .C1(new_n477), .C2(new_n485), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n353), .A2(new_n713), .A3(KEYINPUT42), .A4(new_n676), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G131), .ZN(G33));
  INV_X1    g530(.A(new_n646), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n710), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(new_n204), .ZN(G36));
  INV_X1    g533(.A(KEYINPUT45), .ZN(new_n720));
  OR2_X1    g534(.A1(new_n664), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n664), .A2(new_n720), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n721), .A2(G469), .A3(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT102), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n721), .A2(KEYINPUT102), .A3(G469), .A4(new_n722), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n660), .A2(new_n274), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(KEYINPUT46), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT46), .ZN(new_n731));
  AOI211_X1 g545(.A(new_n731), .B(new_n728), .C1(new_n725), .C2(new_n726), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n730), .A2(new_n732), .A3(new_n666), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n733), .A2(new_n357), .A3(new_n668), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n608), .B1(new_n581), .B2(new_n604), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(G478), .A3(new_n274), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n736), .B1(G478), .B2(new_n583), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n544), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT43), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n737), .A2(KEYINPUT104), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT104), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n610), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n740), .A2(new_n742), .A3(new_n544), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n739), .B1(KEYINPUT103), .B2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT103), .ZN(new_n745));
  AOI21_X1  g559(.A(KEYINPUT43), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n747), .B(new_n657), .C1(new_n615), .C2(new_n613), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n734), .A2(new_n750), .ZN(new_n751));
  XOR2_X1   g565(.A(new_n708), .B(KEYINPUT105), .Z(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n753), .B1(new_n748), .B2(new_n749), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(new_n206), .ZN(G39));
  INV_X1    g570(.A(KEYINPUT47), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n757), .B1(new_n733), .B2(new_n357), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n727), .A2(new_n729), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n731), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n727), .A2(KEYINPUT46), .A3(new_n729), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n485), .A3(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n762), .A2(KEYINPUT47), .A3(new_n356), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n758), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n308), .A2(new_n352), .A3(new_n676), .A4(new_n709), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(KEYINPUT106), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G140), .ZN(G42));
  NAND2_X1  g582(.A1(new_n588), .A2(new_n268), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT112), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n747), .A2(new_n592), .A3(new_n681), .A4(new_n698), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n650), .A2(new_n358), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n770), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT50), .ZN(new_n775));
  INV_X1    g589(.A(new_n592), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n612), .A2(new_n702), .A3(new_n703), .ZN(new_n777));
  NOR4_X1   g591(.A1(new_n744), .A2(new_n746), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n778), .A2(KEYINPUT112), .A3(new_n681), .A4(new_n772), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n774), .A2(new_n775), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT113), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT113), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n774), .A2(new_n782), .A3(new_n775), .A4(new_n779), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n771), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n785), .A2(KEYINPUT50), .A3(new_n772), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT114), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT115), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT51), .ZN(new_n789));
  AOI22_X1  g603(.A1(new_n784), .A2(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n744), .A2(new_n776), .A3(new_n746), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n680), .A2(new_n485), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n792), .A2(new_n357), .A3(new_n708), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n791), .A2(KEYINPUT116), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT116), .B1(new_n791), .B2(new_n793), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n613), .A2(new_n697), .A3(new_n630), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n352), .A2(new_n776), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n793), .A2(new_n656), .A3(new_n799), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n800), .A2(new_n545), .A3(new_n737), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n680), .A2(new_n357), .A3(new_n485), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n758), .A2(new_n763), .A3(new_n804), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n778), .A2(new_n753), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n803), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n790), .B1(new_n807), .B2(new_n789), .ZN(new_n808));
  OR3_X1    g622(.A1(new_n800), .A2(new_n544), .A3(new_n610), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n796), .A2(new_n353), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n810), .A2(KEYINPUT48), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(KEYINPUT48), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n591), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n808), .A2(new_n809), .A3(new_n813), .ZN(new_n814));
  AND4_X1   g628(.A1(new_n685), .A2(new_n692), .A3(new_n688), .A4(new_n699), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n715), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n657), .B1(new_n641), .B2(new_n655), .ZN(new_n817));
  INV_X1    g631(.A(new_n645), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n817), .A2(new_n600), .A3(new_n818), .A4(new_n694), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n691), .A2(new_n676), .A3(new_n797), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n647), .A2(new_n819), .A3(new_n677), .A4(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT52), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n637), .B(new_n356), .C1(new_n665), .C2(new_n666), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n824), .A2(new_n308), .A3(new_n630), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n705), .B1(new_n825), .B2(new_n646), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n826), .A2(KEYINPUT52), .A3(new_n677), .A4(new_n819), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n816), .B1(new_n823), .B2(new_n827), .ZN(new_n828));
  AND4_X1   g642(.A1(new_n684), .A2(new_n600), .A3(new_n657), .A4(new_n709), .ZN(new_n829));
  AND4_X1   g643(.A1(new_n585), .A2(new_n620), .A3(new_n586), .A4(new_n621), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n829), .A2(KEYINPUT108), .A3(new_n818), .A4(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n713), .A2(new_n643), .A3(new_n818), .A4(new_n830), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT108), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n713), .ZN(new_n836));
  OAI22_X1  g650(.A1(new_n710), .A2(new_n717), .B1(new_n836), .B2(new_n704), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n544), .A2(new_n587), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n602), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n600), .A2(new_n612), .A3(new_n841), .A4(new_n616), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT107), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n638), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n844), .A2(new_n617), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n843), .B1(new_n638), .B2(new_n842), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n846), .A2(new_n598), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n839), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n828), .A2(new_n849), .A3(KEYINPUT53), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT109), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n823), .A2(new_n827), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n837), .B1(new_n831), .B2(new_n834), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n844), .A2(new_n617), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n855), .A2(new_n598), .A3(new_n846), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n692), .A2(new_n699), .A3(new_n685), .A4(new_n688), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n857), .B1(new_n712), .B2(new_n714), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n853), .A2(new_n854), .A3(new_n856), .A4(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n851), .A2(new_n852), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n852), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n861), .A2(new_n850), .A3(KEYINPUT109), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n860), .A2(KEYINPUT54), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n758), .A2(KEYINPUT111), .A3(new_n763), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(new_n804), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT111), .B1(new_n758), .B2(new_n763), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n806), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n803), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n784), .A2(new_n787), .A3(new_n788), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n789), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT110), .B1(new_n839), .B2(new_n848), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT110), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n856), .A2(new_n873), .A3(new_n854), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n872), .A2(new_n828), .A3(KEYINPUT53), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n861), .ZN(new_n876));
  OR2_X1    g690(.A1(new_n876), .A2(KEYINPUT54), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n814), .A2(new_n863), .A3(new_n871), .A4(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n771), .A2(new_n426), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n769), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n792), .B(KEYINPUT49), .ZN(new_n881));
  NOR4_X1   g695(.A1(new_n881), .A2(new_n632), .A3(new_n650), .A4(new_n738), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n882), .A2(new_n612), .A3(new_n356), .A4(new_n656), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n880), .A2(new_n883), .ZN(G75));
  AOI21_X1  g698(.A(new_n274), .B1(new_n875), .B2(new_n861), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT56), .B1(new_n885), .B2(G210), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n416), .A2(new_n421), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(new_n419), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT55), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n886), .A2(new_n889), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n268), .A2(G952), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(G51));
  NAND2_X1  g707(.A1(new_n876), .A2(KEYINPUT54), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n877), .A2(KEYINPUT117), .A3(new_n894), .ZN(new_n895));
  OR3_X1    g709(.A1(new_n876), .A2(KEYINPUT117), .A3(KEYINPUT54), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n728), .B(KEYINPUT57), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n898), .A2(new_n482), .A3(new_n483), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n885), .A2(new_n725), .A3(new_n726), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n892), .B1(new_n899), .B2(new_n900), .ZN(G54));
  NAND3_X1  g715(.A1(new_n885), .A2(KEYINPUT58), .A3(G475), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n903));
  INV_X1    g717(.A(new_n541), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n892), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n906), .B1(new_n902), .B2(new_n904), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n903), .B1(new_n902), .B2(new_n904), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n905), .A2(new_n907), .A3(new_n908), .ZN(G60));
  NAND2_X1  g723(.A1(G478), .A2(G902), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT59), .Z(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n895), .A2(new_n896), .A3(new_n735), .A4(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n906), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n911), .B1(new_n863), .B2(new_n877), .ZN(new_n915));
  OR3_X1    g729(.A1(new_n915), .A2(KEYINPUT119), .A3(new_n735), .ZN(new_n916));
  OAI21_X1  g730(.A(KEYINPUT119), .B1(new_n915), .B2(new_n735), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(G63));
  NAND2_X1  g732(.A1(G217), .A2(G902), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT60), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT120), .B1(new_n876), .B2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT120), .ZN(new_n923));
  AOI211_X1 g737(.A(new_n923), .B(new_n920), .C1(new_n875), .C2(new_n861), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n349), .A2(new_n338), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n892), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n629), .B1(new_n922), .B2(new_n924), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT121), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI211_X1 g744(.A(KEYINPUT121), .B(new_n629), .C1(new_n922), .C2(new_n924), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n927), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  XNOR2_X1  g746(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n927), .A2(new_n930), .A3(new_n933), .A4(new_n931), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(G66));
  OAI21_X1  g751(.A(G953), .B1(new_n594), .B2(new_n388), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n848), .A2(new_n857), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n938), .B1(new_n939), .B2(G953), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n887), .B1(G898), .B2(new_n268), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(G69));
  OAI21_X1  g756(.A(new_n840), .B1(new_n544), .B2(new_n610), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n671), .A2(new_n353), .A3(new_n709), .A4(new_n943), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(new_n751), .B2(new_n754), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT123), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT62), .ZN(new_n947));
  INV_X1    g761(.A(new_n674), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n826), .A2(new_n677), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n674), .A2(KEYINPUT62), .A3(new_n677), .A4(new_n826), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n292), .B(new_n532), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n946), .A2(new_n952), .A3(new_n767), .A4(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n734), .A2(new_n353), .A3(new_n694), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT124), .Z(new_n957));
  NOR2_X1   g771(.A1(new_n755), .A2(new_n949), .ZN(new_n958));
  INV_X1    g772(.A(new_n715), .ZN(new_n959));
  AOI211_X1 g773(.A(new_n959), .B(new_n718), .C1(new_n764), .C2(new_n766), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n957), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n955), .B(new_n268), .C1(new_n961), .C2(new_n954), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n954), .A2(G227), .A3(G900), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT125), .ZN(new_n964));
  OAI21_X1  g778(.A(G900), .B1(new_n964), .B2(G227), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n953), .B(new_n965), .C1(new_n964), .C2(G900), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n963), .A2(G953), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n962), .A2(new_n967), .ZN(G72));
  NAND4_X1  g782(.A1(new_n957), .A2(new_n960), .A3(new_n939), .A4(new_n958), .ZN(new_n969));
  XNOR2_X1  g783(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n970));
  NAND2_X1  g784(.A1(G472), .A2(G902), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(new_n972));
  AOI211_X1 g786(.A(new_n270), .B(new_n651), .C1(new_n969), .C2(new_n972), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n946), .A2(new_n952), .A3(new_n767), .A4(new_n939), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n652), .B1(new_n974), .B2(new_n972), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n302), .A2(new_n282), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n860), .A2(new_n862), .A3(new_n972), .A4(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n906), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n973), .A2(new_n975), .A3(new_n978), .ZN(G57));
endmodule


