

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U551 ( .A1(n714), .A2(n713), .ZN(n725) );
  NOR2_X2 U552 ( .A1(n607), .A2(n606), .ZN(n657) );
  NOR2_X2 U553 ( .A1(G2105), .A2(n534), .ZN(n860) );
  XNOR2_X1 U554 ( .A(n643), .B(KEYINPUT26), .ZN(n644) );
  INV_X1 U555 ( .A(KEYINPUT30), .ZN(n616) );
  XNOR2_X1 U556 ( .A(n616), .B(KEYINPUT89), .ZN(n617) );
  XNOR2_X1 U557 ( .A(n618), .B(n617), .ZN(n619) );
  NOR2_X1 U558 ( .A1(n546), .A2(n545), .ZN(G160) );
  NOR2_X1 U559 ( .A1(G651), .A2(G543), .ZN(n766) );
  NAND2_X1 U560 ( .A1(n766), .A2(G89), .ZN(n515) );
  XNOR2_X1 U561 ( .A(n515), .B(KEYINPUT4), .ZN(n517) );
  XOR2_X1 U562 ( .A(G543), .B(KEYINPUT0), .Z(n581) );
  INV_X1 U563 ( .A(G651), .ZN(n520) );
  NOR2_X1 U564 ( .A1(n581), .A2(n520), .ZN(n770) );
  NAND2_X1 U565 ( .A1(G76), .A2(n770), .ZN(n516) );
  NAND2_X1 U566 ( .A1(n517), .A2(n516), .ZN(n519) );
  XOR2_X1 U567 ( .A(KEYINPUT5), .B(KEYINPUT69), .Z(n518) );
  XNOR2_X1 U568 ( .A(n519), .B(n518), .ZN(n529) );
  XNOR2_X1 U569 ( .A(KEYINPUT70), .B(KEYINPUT71), .ZN(n527) );
  NOR2_X2 U570 ( .A1(G651), .A2(n581), .ZN(n771) );
  NAND2_X1 U571 ( .A1(n771), .A2(G51), .ZN(n524) );
  NOR2_X1 U572 ( .A1(G543), .A2(n520), .ZN(n521) );
  XOR2_X1 U573 ( .A(KEYINPUT1), .B(n521), .Z(n522) );
  XNOR2_X1 U574 ( .A(KEYINPUT64), .B(n522), .ZN(n767) );
  NAND2_X1 U575 ( .A1(G63), .A2(n767), .ZN(n523) );
  NAND2_X1 U576 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U577 ( .A(n525), .B(KEYINPUT6), .ZN(n526) );
  XNOR2_X1 U578 ( .A(n527), .B(n526), .ZN(n528) );
  NAND2_X1 U579 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U580 ( .A(n530), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U581 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U582 ( .A(G2104), .ZN(n534) );
  NAND2_X1 U583 ( .A1(G102), .A2(n860), .ZN(n533) );
  NOR2_X1 U584 ( .A1(G2104), .A2(G2105), .ZN(n531) );
  XOR2_X2 U585 ( .A(KEYINPUT17), .B(n531), .Z(n861) );
  NAND2_X1 U586 ( .A1(G138), .A2(n861), .ZN(n532) );
  NAND2_X1 U587 ( .A1(n533), .A2(n532), .ZN(n539) );
  INV_X1 U588 ( .A(G2105), .ZN(n535) );
  NOR2_X1 U589 ( .A1(n534), .A2(n535), .ZN(n868) );
  NAND2_X1 U590 ( .A1(G114), .A2(n868), .ZN(n537) );
  NOR2_X1 U591 ( .A1(G2104), .A2(n535), .ZN(n865) );
  NAND2_X1 U592 ( .A1(G126), .A2(n865), .ZN(n536) );
  NAND2_X1 U593 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U594 ( .A1(n539), .A2(n538), .ZN(G164) );
  NAND2_X1 U595 ( .A1(n865), .A2(G125), .ZN(n542) );
  NAND2_X1 U596 ( .A1(G101), .A2(n860), .ZN(n540) );
  XOR2_X1 U597 ( .A(KEYINPUT23), .B(n540), .Z(n541) );
  NAND2_X1 U598 ( .A1(n542), .A2(n541), .ZN(n546) );
  NAND2_X1 U599 ( .A1(G137), .A2(n861), .ZN(n544) );
  NAND2_X1 U600 ( .A1(G113), .A2(n868), .ZN(n543) );
  NAND2_X1 U601 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U602 ( .A1(G85), .A2(n766), .ZN(n548) );
  NAND2_X1 U603 ( .A1(G72), .A2(n770), .ZN(n547) );
  NAND2_X1 U604 ( .A1(n548), .A2(n547), .ZN(n551) );
  NAND2_X1 U605 ( .A1(G60), .A2(n767), .ZN(n549) );
  XNOR2_X1 U606 ( .A(KEYINPUT65), .B(n549), .ZN(n550) );
  NOR2_X1 U607 ( .A1(n551), .A2(n550), .ZN(n553) );
  NAND2_X1 U608 ( .A1(n771), .A2(G47), .ZN(n552) );
  NAND2_X1 U609 ( .A1(n553), .A2(n552), .ZN(G290) );
  NAND2_X1 U610 ( .A1(n766), .A2(G86), .ZN(n555) );
  NAND2_X1 U611 ( .A1(G61), .A2(n767), .ZN(n554) );
  NAND2_X1 U612 ( .A1(n555), .A2(n554), .ZN(n558) );
  NAND2_X1 U613 ( .A1(n770), .A2(G73), .ZN(n556) );
  XOR2_X1 U614 ( .A(KEYINPUT2), .B(n556), .Z(n557) );
  NOR2_X1 U615 ( .A1(n558), .A2(n557), .ZN(n560) );
  NAND2_X1 U616 ( .A1(n771), .A2(G48), .ZN(n559) );
  NAND2_X1 U617 ( .A1(n560), .A2(n559), .ZN(G305) );
  NAND2_X1 U618 ( .A1(n770), .A2(G75), .ZN(n562) );
  NAND2_X1 U619 ( .A1(G62), .A2(n767), .ZN(n561) );
  NAND2_X1 U620 ( .A1(n562), .A2(n561), .ZN(n565) );
  NAND2_X1 U621 ( .A1(G88), .A2(n766), .ZN(n563) );
  XNOR2_X1 U622 ( .A(KEYINPUT77), .B(n563), .ZN(n564) );
  NOR2_X1 U623 ( .A1(n565), .A2(n564), .ZN(n567) );
  NAND2_X1 U624 ( .A1(n771), .A2(G50), .ZN(n566) );
  NAND2_X1 U625 ( .A1(n567), .A2(n566), .ZN(G303) );
  INV_X1 U626 ( .A(G303), .ZN(G166) );
  NAND2_X1 U627 ( .A1(G90), .A2(n766), .ZN(n569) );
  NAND2_X1 U628 ( .A1(G77), .A2(n770), .ZN(n568) );
  NAND2_X1 U629 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U630 ( .A(KEYINPUT9), .B(n570), .ZN(n574) );
  NAND2_X1 U631 ( .A1(n767), .A2(G64), .ZN(n572) );
  NAND2_X1 U632 ( .A1(n771), .A2(G52), .ZN(n571) );
  AND2_X1 U633 ( .A1(n572), .A2(n571), .ZN(n573) );
  NAND2_X1 U634 ( .A1(n574), .A2(n573), .ZN(G301) );
  NAND2_X1 U635 ( .A1(n766), .A2(G91), .ZN(n576) );
  NAND2_X1 U636 ( .A1(G65), .A2(n767), .ZN(n575) );
  NAND2_X1 U637 ( .A1(n576), .A2(n575), .ZN(n580) );
  NAND2_X1 U638 ( .A1(G78), .A2(n770), .ZN(n578) );
  NAND2_X1 U639 ( .A1(G53), .A2(n771), .ZN(n577) );
  NAND2_X1 U640 ( .A1(n578), .A2(n577), .ZN(n579) );
  OR2_X1 U641 ( .A1(n580), .A2(n579), .ZN(G299) );
  NAND2_X1 U642 ( .A1(G87), .A2(n581), .ZN(n583) );
  NAND2_X1 U643 ( .A1(G74), .A2(G651), .ZN(n582) );
  NAND2_X1 U644 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U645 ( .A1(n767), .A2(n584), .ZN(n586) );
  NAND2_X1 U646 ( .A1(n771), .A2(G49), .ZN(n585) );
  NAND2_X1 U647 ( .A1(n586), .A2(n585), .ZN(G288) );
  NOR2_X1 U648 ( .A1(G164), .A2(G1384), .ZN(n605) );
  NAND2_X1 U649 ( .A1(G160), .A2(G40), .ZN(n606) );
  NOR2_X1 U650 ( .A1(n605), .A2(n606), .ZN(n737) );
  NAND2_X1 U651 ( .A1(G95), .A2(n860), .ZN(n588) );
  NAND2_X1 U652 ( .A1(G107), .A2(n868), .ZN(n587) );
  NAND2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U654 ( .A1(G131), .A2(n861), .ZN(n589) );
  XNOR2_X1 U655 ( .A(KEYINPUT83), .B(n589), .ZN(n590) );
  NOR2_X1 U656 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U657 ( .A1(n865), .A2(G119), .ZN(n592) );
  NAND2_X1 U658 ( .A1(n593), .A2(n592), .ZN(n844) );
  NAND2_X1 U659 ( .A1(G1991), .A2(n844), .ZN(n603) );
  NAND2_X1 U660 ( .A1(G117), .A2(n868), .ZN(n595) );
  NAND2_X1 U661 ( .A1(G129), .A2(n865), .ZN(n594) );
  NAND2_X1 U662 ( .A1(n595), .A2(n594), .ZN(n598) );
  NAND2_X1 U663 ( .A1(n860), .A2(G105), .ZN(n596) );
  XOR2_X1 U664 ( .A(KEYINPUT38), .B(n596), .Z(n597) );
  NOR2_X1 U665 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U666 ( .A(n599), .B(KEYINPUT84), .ZN(n601) );
  NAND2_X1 U667 ( .A1(G141), .A2(n861), .ZN(n600) );
  NAND2_X1 U668 ( .A1(n601), .A2(n600), .ZN(n849) );
  NAND2_X1 U669 ( .A1(G1996), .A2(n849), .ZN(n602) );
  NAND2_X1 U670 ( .A1(n603), .A2(n602), .ZN(n985) );
  NAND2_X1 U671 ( .A1(n737), .A2(n985), .ZN(n729) );
  XNOR2_X1 U672 ( .A(G1986), .B(G290), .ZN(n929) );
  NAND2_X1 U673 ( .A1(n737), .A2(n929), .ZN(n604) );
  NAND2_X1 U674 ( .A1(n729), .A2(n604), .ZN(n714) );
  OR2_X1 U675 ( .A1(G305), .A2(G1981), .ZN(n697) );
  XOR2_X1 U676 ( .A(KEYINPUT24), .B(n697), .Z(n608) );
  INV_X1 U677 ( .A(n605), .ZN(n607) );
  INV_X1 U678 ( .A(n657), .ZN(n675) );
  NAND2_X1 U679 ( .A1(n675), .A2(G8), .ZN(n614) );
  INV_X1 U680 ( .A(n614), .ZN(n704) );
  NAND2_X1 U681 ( .A1(n608), .A2(n704), .ZN(n695) );
  NAND2_X1 U682 ( .A1(G8), .A2(G166), .ZN(n609) );
  NOR2_X1 U683 ( .A1(G2090), .A2(n609), .ZN(n610) );
  XNOR2_X1 U684 ( .A(n610), .B(KEYINPUT95), .ZN(n692) );
  NAND2_X1 U685 ( .A1(G1961), .A2(n675), .ZN(n612) );
  XOR2_X1 U686 ( .A(G2078), .B(KEYINPUT25), .Z(n907) );
  NAND2_X1 U687 ( .A1(n657), .A2(n907), .ZN(n611) );
  NAND2_X1 U688 ( .A1(n612), .A2(n611), .ZN(n670) );
  NAND2_X1 U689 ( .A1(G301), .A2(n670), .ZN(n613) );
  XNOR2_X1 U690 ( .A(KEYINPUT91), .B(n613), .ZN(n622) );
  NOR2_X1 U691 ( .A1(G1966), .A2(n614), .ZN(n687) );
  NOR2_X1 U692 ( .A1(G2084), .A2(n675), .ZN(n684) );
  NOR2_X1 U693 ( .A1(n687), .A2(n684), .ZN(n615) );
  NAND2_X1 U694 ( .A1(G8), .A2(n615), .ZN(n618) );
  NOR2_X1 U695 ( .A1(G168), .A2(n619), .ZN(n620) );
  XNOR2_X1 U696 ( .A(n620), .B(KEYINPUT90), .ZN(n621) );
  NOR2_X1 U697 ( .A1(n622), .A2(n621), .ZN(n624) );
  XOR2_X1 U698 ( .A(KEYINPUT92), .B(KEYINPUT31), .Z(n623) );
  XNOR2_X1 U699 ( .A(n624), .B(n623), .ZN(n674) );
  XNOR2_X1 U700 ( .A(KEYINPUT29), .B(KEYINPUT88), .ZN(n669) );
  NAND2_X1 U701 ( .A1(n767), .A2(G66), .ZN(n625) );
  XNOR2_X1 U702 ( .A(n625), .B(KEYINPUT66), .ZN(n632) );
  NAND2_X1 U703 ( .A1(G92), .A2(n766), .ZN(n627) );
  NAND2_X1 U704 ( .A1(G79), .A2(n770), .ZN(n626) );
  NAND2_X1 U705 ( .A1(n627), .A2(n626), .ZN(n630) );
  NAND2_X1 U706 ( .A1(G54), .A2(n771), .ZN(n628) );
  XNOR2_X1 U707 ( .A(KEYINPUT67), .B(n628), .ZN(n629) );
  NOR2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U709 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U710 ( .A(KEYINPUT15), .B(n633), .ZN(n928) );
  NAND2_X1 U711 ( .A1(n767), .A2(G56), .ZN(n634) );
  XOR2_X1 U712 ( .A(KEYINPUT14), .B(n634), .Z(n640) );
  NAND2_X1 U713 ( .A1(n766), .A2(G81), .ZN(n635) );
  XNOR2_X1 U714 ( .A(n635), .B(KEYINPUT12), .ZN(n637) );
  NAND2_X1 U715 ( .A1(G68), .A2(n770), .ZN(n636) );
  NAND2_X1 U716 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U717 ( .A(KEYINPUT13), .B(n638), .Z(n639) );
  NOR2_X1 U718 ( .A1(n640), .A2(n639), .ZN(n642) );
  NAND2_X1 U719 ( .A1(n771), .A2(G43), .ZN(n641) );
  NAND2_X1 U720 ( .A1(n642), .A2(n641), .ZN(n940) );
  AND2_X1 U721 ( .A1(n657), .A2(G1996), .ZN(n643) );
  INV_X1 U722 ( .A(n644), .ZN(n646) );
  NAND2_X1 U723 ( .A1(n675), .A2(G1341), .ZN(n645) );
  NAND2_X1 U724 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U725 ( .A1(n940), .A2(n647), .ZN(n648) );
  OR2_X1 U726 ( .A1(n928), .A2(n648), .ZN(n655) );
  NAND2_X1 U727 ( .A1(n928), .A2(n648), .ZN(n653) );
  AND2_X1 U728 ( .A1(n657), .A2(G2067), .ZN(n649) );
  XNOR2_X1 U729 ( .A(n649), .B(KEYINPUT85), .ZN(n651) );
  NAND2_X1 U730 ( .A1(n675), .A2(G1348), .ZN(n650) );
  NAND2_X1 U731 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U732 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U733 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U734 ( .A(KEYINPUT86), .B(n656), .Z(n663) );
  NAND2_X1 U735 ( .A1(n657), .A2(G2072), .ZN(n658) );
  XOR2_X1 U736 ( .A(KEYINPUT27), .B(n658), .Z(n660) );
  NAND2_X1 U737 ( .A1(G1956), .A2(n675), .ZN(n659) );
  NAND2_X1 U738 ( .A1(n660), .A2(n659), .ZN(n664) );
  NOR2_X1 U739 ( .A1(G299), .A2(n664), .ZN(n661) );
  XOR2_X1 U740 ( .A(KEYINPUT87), .B(n661), .Z(n662) );
  NOR2_X1 U741 ( .A1(n663), .A2(n662), .ZN(n667) );
  NAND2_X1 U742 ( .A1(G299), .A2(n664), .ZN(n665) );
  XOR2_X1 U743 ( .A(KEYINPUT28), .B(n665), .Z(n666) );
  NOR2_X1 U744 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U745 ( .A(n669), .B(n668), .ZN(n672) );
  OR2_X1 U746 ( .A1(n670), .A2(G301), .ZN(n671) );
  NAND2_X1 U747 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U748 ( .A1(n674), .A2(n673), .ZN(n685) );
  NAND2_X1 U749 ( .A1(n685), .A2(G286), .ZN(n681) );
  NOR2_X1 U750 ( .A1(G1971), .A2(n614), .ZN(n677) );
  NOR2_X1 U751 ( .A1(G2090), .A2(n675), .ZN(n676) );
  NOR2_X1 U752 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U753 ( .A1(n678), .A2(G303), .ZN(n679) );
  XOR2_X1 U754 ( .A(KEYINPUT93), .B(n679), .Z(n680) );
  NAND2_X1 U755 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U756 ( .A1(n682), .A2(G8), .ZN(n683) );
  XNOR2_X1 U757 ( .A(n683), .B(KEYINPUT32), .ZN(n691) );
  NAND2_X1 U758 ( .A1(G8), .A2(n684), .ZN(n689) );
  INV_X1 U759 ( .A(n685), .ZN(n686) );
  NOR2_X1 U760 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U761 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U762 ( .A1(n691), .A2(n690), .ZN(n699) );
  NAND2_X1 U763 ( .A1(n692), .A2(n699), .ZN(n693) );
  NAND2_X1 U764 ( .A1(n614), .A2(n693), .ZN(n694) );
  NAND2_X1 U765 ( .A1(n695), .A2(n694), .ZN(n712) );
  NAND2_X1 U766 ( .A1(G1981), .A2(G305), .ZN(n696) );
  NAND2_X1 U767 ( .A1(n697), .A2(n696), .ZN(n942) );
  NOR2_X1 U768 ( .A1(G1976), .A2(G288), .ZN(n703) );
  NOR2_X1 U769 ( .A1(G1971), .A2(G303), .ZN(n698) );
  NOR2_X1 U770 ( .A1(n703), .A2(n698), .ZN(n927) );
  NAND2_X1 U771 ( .A1(n699), .A2(n927), .ZN(n701) );
  AND2_X1 U772 ( .A1(G1976), .A2(G288), .ZN(n930) );
  NOR2_X1 U773 ( .A1(n930), .A2(n614), .ZN(n700) );
  NAND2_X1 U774 ( .A1(n701), .A2(n700), .ZN(n702) );
  INV_X1 U775 ( .A(KEYINPUT33), .ZN(n706) );
  NAND2_X1 U776 ( .A1(n702), .A2(n706), .ZN(n709) );
  NAND2_X1 U777 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U778 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U779 ( .A(n707), .B(KEYINPUT94), .Z(n708) );
  NAND2_X1 U780 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U781 ( .A1(n942), .A2(n710), .ZN(n711) );
  NOR2_X1 U782 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U783 ( .A(G2067), .B(KEYINPUT37), .ZN(n735) );
  NAND2_X1 U784 ( .A1(n860), .A2(G104), .ZN(n715) );
  XNOR2_X1 U785 ( .A(n715), .B(KEYINPUT82), .ZN(n717) );
  NAND2_X1 U786 ( .A1(G140), .A2(n861), .ZN(n716) );
  NAND2_X1 U787 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U788 ( .A(KEYINPUT34), .B(n718), .ZN(n723) );
  NAND2_X1 U789 ( .A1(G116), .A2(n868), .ZN(n720) );
  NAND2_X1 U790 ( .A1(G128), .A2(n865), .ZN(n719) );
  NAND2_X1 U791 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U792 ( .A(KEYINPUT35), .B(n721), .Z(n722) );
  NOR2_X1 U793 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U794 ( .A(KEYINPUT36), .B(n724), .ZN(n875) );
  NOR2_X1 U795 ( .A1(n735), .A2(n875), .ZN(n988) );
  NAND2_X1 U796 ( .A1(n737), .A2(n988), .ZN(n734) );
  NAND2_X1 U797 ( .A1(n725), .A2(n734), .ZN(n726) );
  XNOR2_X1 U798 ( .A(n726), .B(KEYINPUT96), .ZN(n740) );
  NOR2_X1 U799 ( .A1(G1986), .A2(G290), .ZN(n727) );
  NOR2_X1 U800 ( .A1(G1991), .A2(n844), .ZN(n982) );
  NOR2_X1 U801 ( .A1(n727), .A2(n982), .ZN(n728) );
  XNOR2_X1 U802 ( .A(n728), .B(KEYINPUT97), .ZN(n730) );
  NAND2_X1 U803 ( .A1(n730), .A2(n729), .ZN(n731) );
  OR2_X1 U804 ( .A1(n849), .A2(G1996), .ZN(n979) );
  NAND2_X1 U805 ( .A1(n731), .A2(n979), .ZN(n732) );
  XOR2_X1 U806 ( .A(KEYINPUT39), .B(n732), .Z(n733) );
  NAND2_X1 U807 ( .A1(n734), .A2(n733), .ZN(n736) );
  NAND2_X1 U808 ( .A1(n735), .A2(n875), .ZN(n992) );
  NAND2_X1 U809 ( .A1(n736), .A2(n992), .ZN(n738) );
  NAND2_X1 U810 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U811 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U812 ( .A(n741), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U813 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U814 ( .A(G132), .ZN(G219) );
  INV_X1 U815 ( .A(G82), .ZN(G220) );
  INV_X1 U816 ( .A(G120), .ZN(G236) );
  INV_X1 U817 ( .A(G69), .ZN(G235) );
  INV_X1 U818 ( .A(G57), .ZN(G237) );
  NAND2_X1 U819 ( .A1(G7), .A2(G661), .ZN(n742) );
  XNOR2_X1 U820 ( .A(n742), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U821 ( .A(G223), .ZN(n809) );
  NAND2_X1 U822 ( .A1(n809), .A2(G567), .ZN(n743) );
  XOR2_X1 U823 ( .A(KEYINPUT11), .B(n743), .Z(G234) );
  INV_X1 U824 ( .A(G860), .ZN(n778) );
  OR2_X1 U825 ( .A1(n940), .A2(n778), .ZN(G153) );
  INV_X1 U826 ( .A(G868), .ZN(n790) );
  AND2_X1 U827 ( .A1(n790), .A2(n928), .ZN(n745) );
  NOR2_X1 U828 ( .A1(n790), .A2(G301), .ZN(n744) );
  NOR2_X1 U829 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U830 ( .A(KEYINPUT68), .B(n746), .ZN(G284) );
  NOR2_X1 U831 ( .A1(G286), .A2(n790), .ZN(n748) );
  NOR2_X1 U832 ( .A1(G868), .A2(G299), .ZN(n747) );
  NOR2_X1 U833 ( .A1(n748), .A2(n747), .ZN(G297) );
  NAND2_X1 U834 ( .A1(n778), .A2(G559), .ZN(n749) );
  NAND2_X1 U835 ( .A1(n749), .A2(n928), .ZN(n750) );
  XNOR2_X1 U836 ( .A(n750), .B(KEYINPUT16), .ZN(n751) );
  XNOR2_X1 U837 ( .A(KEYINPUT72), .B(n751), .ZN(G148) );
  NOR2_X1 U838 ( .A1(G559), .A2(n790), .ZN(n752) );
  NAND2_X1 U839 ( .A1(n928), .A2(n752), .ZN(n753) );
  XNOR2_X1 U840 ( .A(n753), .B(KEYINPUT73), .ZN(n755) );
  NOR2_X1 U841 ( .A1(n940), .A2(G868), .ZN(n754) );
  NOR2_X1 U842 ( .A1(n755), .A2(n754), .ZN(G282) );
  NAND2_X1 U843 ( .A1(G99), .A2(n860), .ZN(n757) );
  NAND2_X1 U844 ( .A1(G111), .A2(n868), .ZN(n756) );
  NAND2_X1 U845 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U846 ( .A(KEYINPUT74), .B(n758), .ZN(n763) );
  NAND2_X1 U847 ( .A1(G123), .A2(n865), .ZN(n759) );
  XNOR2_X1 U848 ( .A(n759), .B(KEYINPUT18), .ZN(n761) );
  NAND2_X1 U849 ( .A1(n861), .A2(G135), .ZN(n760) );
  NAND2_X1 U850 ( .A1(n761), .A2(n760), .ZN(n762) );
  NOR2_X1 U851 ( .A1(n763), .A2(n762), .ZN(n981) );
  XNOR2_X1 U852 ( .A(n981), .B(G2096), .ZN(n765) );
  INV_X1 U853 ( .A(G2100), .ZN(n764) );
  NAND2_X1 U854 ( .A1(n765), .A2(n764), .ZN(G156) );
  NAND2_X1 U855 ( .A1(n766), .A2(G93), .ZN(n769) );
  NAND2_X1 U856 ( .A1(G67), .A2(n767), .ZN(n768) );
  NAND2_X1 U857 ( .A1(n769), .A2(n768), .ZN(n775) );
  NAND2_X1 U858 ( .A1(G80), .A2(n770), .ZN(n773) );
  NAND2_X1 U859 ( .A1(G55), .A2(n771), .ZN(n772) );
  NAND2_X1 U860 ( .A1(n773), .A2(n772), .ZN(n774) );
  OR2_X1 U861 ( .A1(n775), .A2(n774), .ZN(n789) );
  XNOR2_X1 U862 ( .A(n789), .B(KEYINPUT76), .ZN(n780) );
  XNOR2_X1 U863 ( .A(n940), .B(KEYINPUT75), .ZN(n777) );
  NAND2_X1 U864 ( .A1(n928), .A2(G559), .ZN(n776) );
  XNOR2_X1 U865 ( .A(n777), .B(n776), .ZN(n787) );
  NAND2_X1 U866 ( .A1(n787), .A2(n778), .ZN(n779) );
  XNOR2_X1 U867 ( .A(n780), .B(n779), .ZN(G145) );
  XOR2_X1 U868 ( .A(KEYINPUT78), .B(KEYINPUT19), .Z(n781) );
  XNOR2_X1 U869 ( .A(G288), .B(n781), .ZN(n782) );
  XOR2_X1 U870 ( .A(n789), .B(n782), .Z(n784) );
  XOR2_X1 U871 ( .A(G290), .B(G305), .Z(n783) );
  XNOR2_X1 U872 ( .A(n784), .B(n783), .ZN(n785) );
  XNOR2_X1 U873 ( .A(G166), .B(n785), .ZN(n786) );
  XNOR2_X1 U874 ( .A(n786), .B(G299), .ZN(n881) );
  XNOR2_X1 U875 ( .A(n881), .B(n787), .ZN(n788) );
  NAND2_X1 U876 ( .A1(n788), .A2(G868), .ZN(n792) );
  NAND2_X1 U877 ( .A1(n790), .A2(n789), .ZN(n791) );
  NAND2_X1 U878 ( .A1(n792), .A2(n791), .ZN(G295) );
  NAND2_X1 U879 ( .A1(G2078), .A2(G2084), .ZN(n793) );
  XOR2_X1 U880 ( .A(KEYINPUT20), .B(n793), .Z(n794) );
  NAND2_X1 U881 ( .A1(G2090), .A2(n794), .ZN(n795) );
  XNOR2_X1 U882 ( .A(KEYINPUT21), .B(n795), .ZN(n796) );
  NAND2_X1 U883 ( .A1(n796), .A2(G2072), .ZN(n797) );
  XOR2_X1 U884 ( .A(KEYINPUT79), .B(n797), .Z(G158) );
  XNOR2_X1 U885 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U886 ( .A1(G235), .A2(G236), .ZN(n798) );
  XOR2_X1 U887 ( .A(KEYINPUT80), .B(n798), .Z(n799) );
  NOR2_X1 U888 ( .A1(G237), .A2(n799), .ZN(n800) );
  NAND2_X1 U889 ( .A1(G108), .A2(n800), .ZN(n901) );
  NAND2_X1 U890 ( .A1(G567), .A2(n901), .ZN(n805) );
  NOR2_X1 U891 ( .A1(G220), .A2(G219), .ZN(n801) );
  XOR2_X1 U892 ( .A(KEYINPUT22), .B(n801), .Z(n802) );
  NOR2_X1 U893 ( .A1(G218), .A2(n802), .ZN(n803) );
  NAND2_X1 U894 ( .A1(G96), .A2(n803), .ZN(n902) );
  NAND2_X1 U895 ( .A1(G2106), .A2(n902), .ZN(n804) );
  NAND2_X1 U896 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U897 ( .A(KEYINPUT81), .B(n806), .ZN(G319) );
  INV_X1 U898 ( .A(G319), .ZN(n808) );
  NAND2_X1 U899 ( .A1(G661), .A2(G483), .ZN(n807) );
  NOR2_X1 U900 ( .A1(n808), .A2(n807), .ZN(n814) );
  NAND2_X1 U901 ( .A1(n814), .A2(G36), .ZN(G176) );
  INV_X1 U902 ( .A(G301), .ZN(G171) );
  NAND2_X1 U903 ( .A1(G2106), .A2(n809), .ZN(G217) );
  INV_X1 U904 ( .A(G661), .ZN(n811) );
  NAND2_X1 U905 ( .A1(G2), .A2(G15), .ZN(n810) );
  NOR2_X1 U906 ( .A1(n811), .A2(n810), .ZN(n812) );
  XOR2_X1 U907 ( .A(KEYINPUT100), .B(n812), .Z(G259) );
  NAND2_X1 U908 ( .A1(G3), .A2(G1), .ZN(n813) );
  NAND2_X1 U909 ( .A1(n814), .A2(n813), .ZN(G188) );
  XOR2_X1 U910 ( .A(KEYINPUT42), .B(G2090), .Z(n816) );
  XNOR2_X1 U911 ( .A(G2078), .B(G2072), .ZN(n815) );
  XNOR2_X1 U912 ( .A(n816), .B(n815), .ZN(n817) );
  XOR2_X1 U913 ( .A(n817), .B(G2100), .Z(n819) );
  XNOR2_X1 U914 ( .A(G2067), .B(G2084), .ZN(n818) );
  XNOR2_X1 U915 ( .A(n819), .B(n818), .ZN(n823) );
  XOR2_X1 U916 ( .A(G2096), .B(KEYINPUT43), .Z(n821) );
  XNOR2_X1 U917 ( .A(KEYINPUT101), .B(G2678), .ZN(n820) );
  XNOR2_X1 U918 ( .A(n821), .B(n820), .ZN(n822) );
  XOR2_X1 U919 ( .A(n823), .B(n822), .Z(G227) );
  XOR2_X1 U920 ( .A(G1976), .B(G1971), .Z(n825) );
  XNOR2_X1 U921 ( .A(G1986), .B(G1956), .ZN(n824) );
  XNOR2_X1 U922 ( .A(n825), .B(n824), .ZN(n835) );
  XOR2_X1 U923 ( .A(KEYINPUT104), .B(KEYINPUT102), .Z(n827) );
  XNOR2_X1 U924 ( .A(G1996), .B(G2474), .ZN(n826) );
  XNOR2_X1 U925 ( .A(n827), .B(n826), .ZN(n831) );
  XOR2_X1 U926 ( .A(G1981), .B(G1961), .Z(n829) );
  XNOR2_X1 U927 ( .A(G1991), .B(G1966), .ZN(n828) );
  XNOR2_X1 U928 ( .A(n829), .B(n828), .ZN(n830) );
  XOR2_X1 U929 ( .A(n831), .B(n830), .Z(n833) );
  XNOR2_X1 U930 ( .A(KEYINPUT103), .B(KEYINPUT41), .ZN(n832) );
  XNOR2_X1 U931 ( .A(n833), .B(n832), .ZN(n834) );
  XNOR2_X1 U932 ( .A(n835), .B(n834), .ZN(G229) );
  NAND2_X1 U933 ( .A1(G124), .A2(n865), .ZN(n836) );
  XNOR2_X1 U934 ( .A(n836), .B(KEYINPUT44), .ZN(n838) );
  NAND2_X1 U935 ( .A1(n860), .A2(G100), .ZN(n837) );
  NAND2_X1 U936 ( .A1(n838), .A2(n837), .ZN(n842) );
  NAND2_X1 U937 ( .A1(G136), .A2(n861), .ZN(n840) );
  NAND2_X1 U938 ( .A1(G112), .A2(n868), .ZN(n839) );
  NAND2_X1 U939 ( .A1(n840), .A2(n839), .ZN(n841) );
  NOR2_X1 U940 ( .A1(n842), .A2(n841), .ZN(G162) );
  XOR2_X1 U941 ( .A(G162), .B(n981), .Z(n851) );
  XOR2_X1 U942 ( .A(KEYINPUT106), .B(KEYINPUT108), .Z(n843) );
  XNOR2_X1 U943 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U944 ( .A(n845), .B(KEYINPUT48), .Z(n847) );
  XNOR2_X1 U945 ( .A(G164), .B(KEYINPUT46), .ZN(n846) );
  XNOR2_X1 U946 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U947 ( .A(n849), .B(n848), .Z(n850) );
  XNOR2_X1 U948 ( .A(n851), .B(n850), .ZN(n877) );
  NAND2_X1 U949 ( .A1(G103), .A2(n860), .ZN(n853) );
  NAND2_X1 U950 ( .A1(G139), .A2(n861), .ZN(n852) );
  NAND2_X1 U951 ( .A1(n853), .A2(n852), .ZN(n859) );
  NAND2_X1 U952 ( .A1(G115), .A2(n868), .ZN(n855) );
  NAND2_X1 U953 ( .A1(G127), .A2(n865), .ZN(n854) );
  NAND2_X1 U954 ( .A1(n855), .A2(n854), .ZN(n856) );
  XNOR2_X1 U955 ( .A(KEYINPUT47), .B(n856), .ZN(n857) );
  XNOR2_X1 U956 ( .A(KEYINPUT107), .B(n857), .ZN(n858) );
  NOR2_X1 U957 ( .A1(n859), .A2(n858), .ZN(n993) );
  XNOR2_X1 U958 ( .A(G160), .B(n993), .ZN(n873) );
  NAND2_X1 U959 ( .A1(G106), .A2(n860), .ZN(n863) );
  NAND2_X1 U960 ( .A1(G142), .A2(n861), .ZN(n862) );
  NAND2_X1 U961 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U962 ( .A(n864), .B(KEYINPUT45), .ZN(n867) );
  NAND2_X1 U963 ( .A1(G130), .A2(n865), .ZN(n866) );
  NAND2_X1 U964 ( .A1(n867), .A2(n866), .ZN(n871) );
  NAND2_X1 U965 ( .A1(G118), .A2(n868), .ZN(n869) );
  XNOR2_X1 U966 ( .A(KEYINPUT105), .B(n869), .ZN(n870) );
  NOR2_X1 U967 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U968 ( .A(n873), .B(n872), .ZN(n874) );
  XNOR2_X1 U969 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U970 ( .A(n877), .B(n876), .ZN(n878) );
  NOR2_X1 U971 ( .A1(G37), .A2(n878), .ZN(G395) );
  XNOR2_X1 U972 ( .A(n940), .B(G286), .ZN(n880) );
  XNOR2_X1 U973 ( .A(G171), .B(n928), .ZN(n879) );
  XNOR2_X1 U974 ( .A(n880), .B(n879), .ZN(n882) );
  XNOR2_X1 U975 ( .A(n882), .B(n881), .ZN(n883) );
  NOR2_X1 U976 ( .A1(G37), .A2(n883), .ZN(n884) );
  XOR2_X1 U977 ( .A(KEYINPUT109), .B(n884), .Z(G397) );
  XNOR2_X1 U978 ( .A(G2451), .B(G2446), .ZN(n894) );
  XOR2_X1 U979 ( .A(G2430), .B(G2443), .Z(n886) );
  XNOR2_X1 U980 ( .A(G2454), .B(G2435), .ZN(n885) );
  XNOR2_X1 U981 ( .A(n886), .B(n885), .ZN(n890) );
  XOR2_X1 U982 ( .A(G2438), .B(KEYINPUT98), .Z(n888) );
  XNOR2_X1 U983 ( .A(G1341), .B(G1348), .ZN(n887) );
  XNOR2_X1 U984 ( .A(n888), .B(n887), .ZN(n889) );
  XOR2_X1 U985 ( .A(n890), .B(n889), .Z(n892) );
  XNOR2_X1 U986 ( .A(KEYINPUT99), .B(G2427), .ZN(n891) );
  XNOR2_X1 U987 ( .A(n892), .B(n891), .ZN(n893) );
  XNOR2_X1 U988 ( .A(n894), .B(n893), .ZN(n895) );
  NAND2_X1 U989 ( .A1(n895), .A2(G14), .ZN(n903) );
  NAND2_X1 U990 ( .A1(G319), .A2(n903), .ZN(n898) );
  NOR2_X1 U991 ( .A1(G227), .A2(G229), .ZN(n896) );
  XNOR2_X1 U992 ( .A(KEYINPUT49), .B(n896), .ZN(n897) );
  NOR2_X1 U993 ( .A1(n898), .A2(n897), .ZN(n900) );
  NOR2_X1 U994 ( .A1(G395), .A2(G397), .ZN(n899) );
  NAND2_X1 U995 ( .A1(n900), .A2(n899), .ZN(G225) );
  XOR2_X1 U996 ( .A(KEYINPUT110), .B(G225), .Z(G308) );
  XNOR2_X1 U997 ( .A(G108), .B(KEYINPUT111), .ZN(G238) );
  INV_X1 U999 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1000 ( .A1(n902), .A2(n901), .ZN(G325) );
  INV_X1 U1001 ( .A(G325), .ZN(G261) );
  INV_X1 U1002 ( .A(n903), .ZN(G401) );
  XOR2_X1 U1003 ( .A(G2084), .B(G34), .Z(n904) );
  XNOR2_X1 U1004 ( .A(KEYINPUT54), .B(n904), .ZN(n921) );
  XNOR2_X1 U1005 ( .A(G2090), .B(G35), .ZN(n919) );
  XOR2_X1 U1006 ( .A(G1991), .B(G25), .Z(n905) );
  NAND2_X1 U1007 ( .A1(G28), .A2(n905), .ZN(n906) );
  XNOR2_X1 U1008 ( .A(n906), .B(KEYINPUT117), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(G1996), .B(G32), .ZN(n909) );
  XNOR2_X1 U1010 ( .A(n907), .B(G27), .ZN(n908) );
  NOR2_X1 U1011 ( .A1(n909), .A2(n908), .ZN(n910) );
  NAND2_X1 U1012 ( .A1(n911), .A2(n910), .ZN(n916) );
  XNOR2_X1 U1013 ( .A(G2067), .B(G26), .ZN(n913) );
  XNOR2_X1 U1014 ( .A(G2072), .B(G33), .ZN(n912) );
  NOR2_X1 U1015 ( .A1(n913), .A2(n912), .ZN(n914) );
  XOR2_X1 U1016 ( .A(KEYINPUT118), .B(n914), .Z(n915) );
  NOR2_X1 U1017 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1018 ( .A(KEYINPUT53), .B(n917), .ZN(n918) );
  NOR2_X1 U1019 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(n922), .B(KEYINPUT119), .ZN(n923) );
  XNOR2_X1 U1022 ( .A(KEYINPUT55), .B(n923), .ZN(n924) );
  INV_X1 U1023 ( .A(G29), .ZN(n1006) );
  NAND2_X1 U1024 ( .A1(n924), .A2(n1006), .ZN(n925) );
  NAND2_X1 U1025 ( .A1(n925), .A2(G11), .ZN(n1012) );
  XNOR2_X1 U1026 ( .A(KEYINPUT56), .B(G16), .ZN(n949) );
  XOR2_X1 U1027 ( .A(G1956), .B(G299), .Z(n926) );
  NAND2_X1 U1028 ( .A1(n927), .A2(n926), .ZN(n938) );
  XNOR2_X1 U1029 ( .A(n928), .B(G1348), .ZN(n936) );
  NOR2_X1 U1030 ( .A1(n930), .A2(n929), .ZN(n932) );
  NAND2_X1 U1031 ( .A1(G1971), .A2(G303), .ZN(n931) );
  NAND2_X1 U1032 ( .A1(n932), .A2(n931), .ZN(n934) );
  XNOR2_X1 U1033 ( .A(G1961), .B(G301), .ZN(n933) );
  NOR2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1036 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1037 ( .A(KEYINPUT120), .B(n939), .ZN(n947) );
  XNOR2_X1 U1038 ( .A(n940), .B(G1341), .ZN(n945) );
  XOR2_X1 U1039 ( .A(G1966), .B(G168), .Z(n941) );
  NOR2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1041 ( .A(KEYINPUT57), .B(n943), .ZN(n944) );
  NOR2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1044 ( .A1(n949), .A2(n948), .ZN(n1010) );
  XOR2_X1 U1045 ( .A(G16), .B(KEYINPUT121), .Z(n975) );
  XNOR2_X1 U1046 ( .A(KEYINPUT124), .B(KEYINPUT125), .ZN(n950) );
  XNOR2_X1 U1047 ( .A(n950), .B(KEYINPUT61), .ZN(n973) );
  XNOR2_X1 U1048 ( .A(KEYINPUT123), .B(G1966), .ZN(n951) );
  XNOR2_X1 U1049 ( .A(n951), .B(G21), .ZN(n964) );
  XOR2_X1 U1050 ( .A(G1348), .B(KEYINPUT59), .Z(n952) );
  XNOR2_X1 U1051 ( .A(G4), .B(n952), .ZN(n959) );
  XOR2_X1 U1052 ( .A(G1956), .B(G20), .Z(n954) );
  XOR2_X1 U1053 ( .A(G1981), .B(G6), .Z(n953) );
  NAND2_X1 U1054 ( .A1(n954), .A2(n953), .ZN(n956) );
  XNOR2_X1 U1055 ( .A(G19), .B(G1341), .ZN(n955) );
  NOR2_X1 U1056 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1057 ( .A(KEYINPUT122), .B(n957), .Z(n958) );
  NOR2_X1 U1058 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1059 ( .A(KEYINPUT60), .B(n960), .Z(n962) );
  XNOR2_X1 U1060 ( .A(G1961), .B(G5), .ZN(n961) );
  NOR2_X1 U1061 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1062 ( .A1(n964), .A2(n963), .ZN(n971) );
  XNOR2_X1 U1063 ( .A(G1971), .B(G22), .ZN(n966) );
  XNOR2_X1 U1064 ( .A(G23), .B(G1976), .ZN(n965) );
  NOR2_X1 U1065 ( .A1(n966), .A2(n965), .ZN(n968) );
  XOR2_X1 U1066 ( .A(G1986), .B(G24), .Z(n967) );
  NAND2_X1 U1067 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1068 ( .A(KEYINPUT58), .B(n969), .ZN(n970) );
  NOR2_X1 U1069 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1070 ( .A(n973), .B(n972), .ZN(n974) );
  NOR2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1072 ( .A(KEYINPUT126), .B(n976), .ZN(n1008) );
  XNOR2_X1 U1073 ( .A(G2090), .B(G162), .ZN(n977) );
  XNOR2_X1 U1074 ( .A(n977), .B(KEYINPUT114), .ZN(n978) );
  NAND2_X1 U1075 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1076 ( .A(n980), .B(KEYINPUT51), .ZN(n1001) );
  NOR2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n987) );
  XOR2_X1 U1078 ( .A(G160), .B(G2084), .Z(n983) );
  XNOR2_X1 U1079 ( .A(KEYINPUT112), .B(n983), .ZN(n984) );
  NOR2_X1 U1080 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n989) );
  NOR2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n990) );
  XOR2_X1 U1083 ( .A(KEYINPUT113), .B(n990), .Z(n991) );
  NAND2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n999) );
  XNOR2_X1 U1085 ( .A(G2072), .B(n993), .ZN(n995) );
  XNOR2_X1 U1086 ( .A(G164), .B(G2078), .ZN(n994) );
  NAND2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1088 ( .A(KEYINPUT50), .B(n996), .Z(n997) );
  XNOR2_X1 U1089 ( .A(KEYINPUT115), .B(n997), .ZN(n998) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(n1002), .B(KEYINPUT116), .ZN(n1003) );
  XNOR2_X1 U1093 ( .A(KEYINPUT52), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1094 ( .A1(KEYINPUT55), .A2(n1004), .ZN(n1005) );
  NOR2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1099 ( .A(KEYINPUT62), .B(n1013), .Z(n1014) );
  XNOR2_X1 U1100 ( .A(KEYINPUT127), .B(n1014), .ZN(G311) );
  INV_X1 U1101 ( .A(G311), .ZN(G150) );
endmodule

