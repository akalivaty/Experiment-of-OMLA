//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 0 0 0 0 1 0 0 1 0 0 0 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 0 1 0 1 1 0 0 0 1 1 1 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:54 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1230, new_n1231,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND3_X1  g0009(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n203), .A2(G50), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n212), .B1(new_n202), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n217));
  INV_X1    g0017(.A(G77), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  INV_X1    g0019(.A(G107), .ZN(new_n220));
  INV_X1    g0020(.A(G264), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n206), .B1(new_n216), .B2(new_n222), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n209), .B1(new_n210), .B2(new_n211), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT64), .ZN(G361));
  XOR2_X1   g0026(.A(G250), .B(G257), .Z(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT65), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G264), .B(G270), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n230), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G50), .B(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT66), .ZN(new_n238));
  XOR2_X1   g0038(.A(G58), .B(G77), .Z(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT67), .ZN(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n240), .B(new_n244), .ZN(G351));
  OAI21_X1  g0045(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n246));
  INV_X1    g0046(.A(G150), .ZN(new_n247));
  NOR2_X1   g0047(.A1(G20), .A2(G33), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT8), .B(G58), .ZN(new_n250));
  INV_X1    g0050(.A(G20), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G33), .ZN(new_n252));
  OAI221_X1 g0052(.A(new_n246), .B1(new_n247), .B2(new_n249), .C1(new_n250), .C2(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G1), .A2(G13), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G50), .ZN(new_n257));
  OR2_X1    g0057(.A1(KEYINPUT68), .A2(G1), .ZN(new_n258));
  NAND2_X1  g0058(.A1(KEYINPUT68), .A2(G1), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n258), .A2(G13), .A3(G20), .A4(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n253), .A2(new_n256), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n256), .ZN(new_n263));
  AND2_X1   g0063(.A1(KEYINPUT68), .A2(G1), .ZN(new_n264));
  NOR2_X1   g0064(.A1(KEYINPUT68), .A2(G1), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G20), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n263), .A2(G50), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT3), .B(G33), .ZN(new_n270));
  NOR2_X1   g0070(.A1(G222), .A2(G1698), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G223), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n270), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n255), .B1(G33), .B2(G41), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n274), .B(new_n275), .C1(G77), .C2(new_n270), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G41), .A2(G45), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n275), .B1(new_n266), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G226), .ZN(new_n280));
  INV_X1    g0080(.A(G33), .ZN(new_n281));
  INV_X1    g0081(.A(G41), .ZN(new_n282));
  OAI211_X1 g0082(.A(G1), .B(G13), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G1), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n283), .A2(new_n284), .A3(G274), .A4(new_n278), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n276), .A2(new_n280), .A3(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G169), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n269), .B(new_n288), .C1(G179), .C2(new_n286), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G190), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n286), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT70), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n286), .A2(G200), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n269), .A2(KEYINPUT9), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n269), .A2(KEYINPUT9), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n293), .B(new_n294), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(KEYINPUT10), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT69), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n300), .B1(new_n296), .B2(new_n297), .ZN(new_n301));
  INV_X1    g0101(.A(new_n297), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n302), .A2(KEYINPUT69), .A3(new_n295), .ZN(new_n303));
  AOI21_X1  g0103(.A(KEYINPUT10), .B1(new_n286), .B2(G200), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n301), .A2(new_n303), .A3(new_n293), .A4(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n290), .B1(new_n299), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n202), .A2(G20), .ZN(new_n307));
  OAI221_X1 g0107(.A(new_n307), .B1(new_n252), .B2(new_n218), .C1(new_n249), .C2(new_n257), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n256), .ZN(new_n309));
  XOR2_X1   g0109(.A(new_n309), .B(KEYINPUT11), .Z(new_n310));
  OAI21_X1  g0110(.A(KEYINPUT12), .B1(new_n260), .B2(G68), .ZN(new_n311));
  OR3_X1    g0111(.A1(new_n260), .A2(KEYINPUT12), .A3(G68), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n263), .A2(G68), .A3(new_n267), .ZN(new_n314));
  XOR2_X1   g0114(.A(new_n314), .B(KEYINPUT71), .Z(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n232), .A2(G1698), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n270), .B(new_n317), .C1(G226), .C2(G1698), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G33), .A2(G97), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n283), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT68), .B(G1), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n283), .B1(new_n321), .B2(new_n277), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n285), .B1(new_n322), .B2(new_n213), .ZN(new_n323));
  OR3_X1    g0123(.A1(new_n320), .A2(new_n323), .A3(KEYINPUT13), .ZN(new_n324));
  OAI21_X1  g0124(.A(KEYINPUT13), .B1(new_n320), .B2(new_n323), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT72), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT14), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n326), .A2(G169), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n324), .A2(G179), .A3(new_n325), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n328), .B1(new_n326), .B2(G169), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n316), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n326), .A2(G200), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n324), .A2(G190), .A3(new_n325), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n313), .A2(new_n334), .A3(new_n315), .A4(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n250), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n339), .A2(new_n248), .B1(G20), .B2(G77), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT15), .B(G87), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n340), .B1(new_n252), .B2(new_n341), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n342), .A2(new_n256), .B1(new_n261), .B2(new_n218), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n263), .A2(G77), .A3(new_n267), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n279), .A2(G244), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n285), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n270), .A2(G238), .A3(G1698), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n270), .A2(G232), .A3(new_n272), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n348), .B(new_n349), .C1(new_n220), .C2(new_n270), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n347), .B1(new_n275), .B2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n345), .B1(new_n351), .B2(G190), .ZN(new_n352));
  INV_X1    g0152(.A(G200), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n352), .B1(new_n353), .B2(new_n351), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n345), .B1(new_n351), .B2(G169), .ZN(new_n355));
  INV_X1    g0155(.A(G179), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n351), .A2(new_n356), .ZN(new_n357));
  OR2_X1    g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n306), .A2(new_n338), .A3(new_n354), .A4(new_n358), .ZN(new_n359));
  OAI211_X1 g0159(.A(G232), .B(new_n283), .C1(new_n321), .C2(new_n277), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n285), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT77), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OR2_X1    g0163(.A1(G223), .A2(G1698), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(G226), .B2(new_n272), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT3), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n366), .A2(KEYINPUT73), .A3(G33), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(G33), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n281), .A2(KEYINPUT3), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT73), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n365), .B1(new_n367), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n281), .A2(new_n214), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n275), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n360), .A2(KEYINPUT77), .A3(new_n285), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n363), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n353), .ZN(new_n377));
  AND3_X1   g0177(.A1(new_n360), .A2(KEYINPUT77), .A3(new_n285), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT77), .B1(new_n360), .B2(new_n285), .ZN(new_n379));
  OAI21_X1  g0179(.A(KEYINPUT78), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT78), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n363), .A2(new_n381), .A3(new_n375), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n374), .A2(new_n291), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n377), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT75), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G58), .A2(G68), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n203), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n386), .B1(new_n388), .B2(new_n251), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n248), .A2(G159), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n203), .A2(new_n387), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n391), .A2(KEYINPUT75), .A3(G20), .ZN(new_n392));
  AND3_X1   g0192(.A1(new_n389), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  AND3_X1   g0193(.A1(new_n371), .A2(KEYINPUT74), .A3(new_n367), .ZN(new_n394));
  AOI21_X1  g0194(.A(KEYINPUT74), .B1(new_n371), .B2(new_n367), .ZN(new_n395));
  NOR2_X1   g0195(.A1(KEYINPUT7), .A2(G20), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NOR3_X1   g0197(.A1(new_n394), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n371), .A2(new_n251), .A3(new_n367), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT7), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(G68), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n393), .B(KEYINPUT16), .C1(new_n398), .C2(new_n401), .ZN(new_n402));
  XNOR2_X1  g0202(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n389), .A2(new_n390), .A3(new_n392), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT7), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(new_n270), .B2(G20), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n368), .A2(new_n369), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n407), .A2(KEYINPUT7), .A3(new_n251), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n202), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n403), .B1(new_n404), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n402), .A2(new_n410), .A3(new_n256), .ZN(new_n411));
  INV_X1    g0211(.A(new_n256), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n267), .A2(new_n412), .A3(new_n339), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(new_n260), .B2(new_n339), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n385), .A2(new_n411), .A3(new_n415), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n416), .B(KEYINPUT17), .ZN(new_n417));
  AND3_X1   g0217(.A1(new_n366), .A2(KEYINPUT73), .A3(G33), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n418), .B1(new_n270), .B2(new_n370), .ZN(new_n419));
  OAI22_X1  g0219(.A1(new_n419), .A2(new_n365), .B1(new_n281), .B2(new_n214), .ZN(new_n420));
  AOI21_X1  g0220(.A(G179), .B1(new_n420), .B2(new_n275), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n380), .A2(new_n382), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n376), .A2(new_n287), .ZN(new_n423));
  AND2_X1   g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n411), .A2(new_n415), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT18), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n424), .A2(new_n425), .A3(KEYINPUT18), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n417), .A2(new_n430), .ZN(new_n431));
  OR3_X1    g0231(.A1(new_n359), .A2(KEYINPUT79), .A3(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(KEYINPUT79), .B1(new_n359), .B2(new_n431), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT6), .ZN(new_n435));
  AND2_X1   g0235(.A1(G97), .A2(G107), .ZN(new_n436));
  NOR2_X1   g0236(.A1(G97), .A2(G107), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(KEYINPUT6), .A2(G97), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT80), .B1(new_n439), .B2(G107), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT80), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n441), .A2(new_n220), .A3(KEYINPUT6), .A4(G97), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n438), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(KEYINPUT81), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT81), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n438), .A2(new_n440), .A3(new_n445), .A4(new_n442), .ZN(new_n446));
  AND3_X1   g0246(.A1(new_n444), .A2(G20), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(KEYINPUT7), .B1(new_n407), .B2(new_n251), .ZN(new_n448));
  AOI211_X1 g0248(.A(new_n405), .B(G20), .C1(new_n368), .C2(new_n369), .ZN(new_n449));
  OAI21_X1  g0249(.A(G107), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n248), .A2(G77), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n256), .B1(new_n447), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n258), .A2(G33), .A3(new_n259), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n260), .A2(new_n412), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G97), .ZN(new_n456));
  INV_X1    g0256(.A(G97), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n260), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT82), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n456), .A2(KEYINPUT82), .A3(new_n458), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n453), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT5), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G41), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n258), .A2(new_n466), .A3(G45), .A4(new_n259), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT84), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT84), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n266), .A2(new_n469), .A3(G45), .A4(new_n466), .ZN(new_n470));
  INV_X1    g0270(.A(G274), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n275), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n282), .A2(KEYINPUT5), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n468), .A2(new_n470), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n468), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n473), .B1(new_n467), .B2(KEYINPUT84), .ZN(new_n476));
  OAI211_X1 g0276(.A(G257), .B(new_n283), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n368), .A2(new_n369), .A3(G250), .A4(G1698), .ZN(new_n478));
  AND2_X1   g0278(.A1(KEYINPUT4), .A2(G244), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n368), .A2(new_n369), .A3(new_n479), .A4(new_n272), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G33), .A2(G283), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n371), .A2(new_n367), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n483), .A2(G244), .A3(new_n272), .ZN(new_n484));
  XNOR2_X1  g0284(.A(KEYINPUT83), .B(KEYINPUT4), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n482), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n474), .B(new_n477), .C1(new_n486), .C2(new_n283), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n287), .ZN(new_n488));
  INV_X1    g0288(.A(new_n485), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n219), .B1(new_n371), .B2(new_n367), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n489), .B1(new_n490), .B2(new_n272), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n275), .B1(new_n491), .B2(new_n482), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n492), .A2(new_n356), .A3(new_n474), .A4(new_n477), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n464), .A2(new_n488), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n444), .A2(new_n446), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n451), .B(new_n450), .C1(new_n495), .C2(new_n251), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n496), .A2(new_n256), .B1(new_n461), .B2(new_n462), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n487), .A2(G200), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n492), .A2(G190), .A3(new_n474), .A4(new_n477), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n341), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(new_n260), .ZN(new_n502));
  AOI21_X1  g0302(.A(G20), .B1(new_n371), .B2(new_n367), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(G68), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT19), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n251), .B1(new_n319), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n437), .A2(new_n214), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n251), .A2(G33), .A3(G97), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n506), .A2(new_n507), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n502), .B1(new_n510), .B2(new_n256), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n341), .B2(new_n455), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n490), .A2(G1698), .B1(G33), .B2(G116), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n483), .A2(G238), .A3(new_n272), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n283), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(G45), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n215), .B1(new_n321), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n266), .A2(G45), .A3(new_n471), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n517), .A2(new_n518), .A3(new_n283), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n287), .B1(new_n515), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n483), .A2(G244), .A3(G1698), .ZN(new_n522));
  NAND2_X1  g0322(.A1(G33), .A2(G116), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n514), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n275), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n525), .A2(new_n356), .A3(new_n519), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n512), .A2(new_n521), .A3(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(G200), .B1(new_n515), .B2(new_n520), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n525), .A2(G190), .A3(new_n519), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n455), .A2(new_n214), .ZN(new_n530));
  AOI211_X1 g0330(.A(new_n502), .B(new_n530), .C1(new_n510), .C2(new_n256), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n528), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  AND4_X1   g0332(.A1(new_n494), .A2(new_n500), .A3(new_n527), .A4(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT24), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT22), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n535), .B1(new_n503), .B2(G87), .ZN(new_n536));
  NOR3_X1   g0336(.A1(new_n214), .A2(KEYINPUT22), .A3(G20), .ZN(new_n537));
  AOI21_X1  g0337(.A(KEYINPUT88), .B1(new_n270), .B2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n270), .A2(KEYINPUT88), .A3(new_n537), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(KEYINPUT89), .B1(new_n536), .B2(new_n541), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n270), .A2(KEYINPUT88), .A3(new_n537), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n543), .A2(new_n538), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT89), .ZN(new_n545));
  AOI211_X1 g0345(.A(G20), .B(new_n214), .C1(new_n371), .C2(new_n367), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n544), .B(new_n545), .C1(new_n546), .C2(new_n535), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n220), .A2(KEYINPUT23), .A3(G20), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(KEYINPUT23), .B1(new_n220), .B2(G20), .ZN(new_n551));
  INV_X1    g0351(.A(G116), .ZN(new_n552));
  OAI22_X1  g0352(.A1(new_n550), .A2(new_n551), .B1(new_n552), .B2(new_n252), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n534), .B1(new_n548), .B2(new_n554), .ZN(new_n555));
  AOI211_X1 g0355(.A(KEYINPUT24), .B(new_n553), .C1(new_n542), .C2(new_n547), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n256), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT25), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n260), .B2(G107), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n261), .A2(KEYINPUT25), .A3(new_n220), .ZN(new_n560));
  INV_X1    g0360(.A(new_n455), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n559), .A2(new_n560), .B1(new_n561), .B2(G107), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G33), .A2(G294), .ZN(new_n563));
  NAND2_X1  g0363(.A1(G257), .A2(G1698), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n563), .B1(new_n419), .B2(new_n564), .ZN(new_n565));
  AOI211_X1 g0365(.A(new_n215), .B(G1698), .C1(new_n371), .C2(new_n367), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n275), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n468), .A2(new_n470), .A3(new_n473), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n568), .A2(G264), .A3(new_n283), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n474), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n353), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(G190), .B2(new_n570), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n557), .A2(new_n562), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n533), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n568), .A2(G270), .A3(new_n283), .ZN(new_n576));
  OR2_X1    g0376(.A1(G257), .A2(G1698), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n221), .A2(G1698), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n579), .B1(new_n371), .B2(new_n367), .ZN(new_n580));
  XNOR2_X1  g0380(.A(KEYINPUT85), .B(G303), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n407), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n275), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n474), .ZN(new_n584));
  OAI21_X1  g0384(.A(G169), .B1(new_n576), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n261), .A2(new_n552), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(new_n552), .B2(new_n455), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n481), .B(new_n251), .C1(G33), .C2(new_n457), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT86), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n552), .A2(G20), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n256), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n589), .B1(new_n256), .B2(new_n590), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n588), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT20), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(KEYINPUT20), .B(new_n588), .C1(new_n591), .C2(new_n592), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n587), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(KEYINPUT87), .B1(new_n585), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(KEYINPUT21), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT21), .ZN(new_n600));
  OAI211_X1 g0400(.A(KEYINPUT87), .B(new_n600), .C1(new_n585), .C2(new_n597), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n568), .A2(G270), .A3(new_n283), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n602), .A2(G179), .A3(new_n474), .A4(new_n583), .ZN(new_n603));
  OR2_X1    g0403(.A1(new_n603), .A2(new_n597), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n599), .A2(new_n601), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n557), .A2(new_n562), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n570), .A2(G169), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(KEYINPUT90), .ZN(new_n608));
  OR2_X1    g0408(.A1(new_n570), .A2(new_n356), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n570), .A2(new_n356), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT90), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n605), .B1(new_n606), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n576), .A2(new_n584), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G190), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n616), .B(new_n597), .C1(new_n353), .C2(new_n615), .ZN(new_n617));
  AND4_X1   g0417(.A1(new_n434), .A2(new_n575), .A3(new_n614), .A4(new_n617), .ZN(G372));
  INV_X1    g0418(.A(new_n527), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT26), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n527), .A2(new_n532), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n620), .B1(new_n621), .B2(new_n494), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n464), .A2(new_n488), .A3(new_n493), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n623), .A2(KEYINPUT26), .A3(new_n527), .A4(new_n532), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n619), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n625), .B1(new_n614), .B2(new_n574), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n434), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n333), .A2(new_n358), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n417), .A2(new_n628), .A3(new_n336), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT74), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n483), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n371), .A2(KEYINPUT74), .A3(new_n367), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n631), .A2(new_n632), .A3(new_n396), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n202), .B1(new_n399), .B2(KEYINPUT7), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n404), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n412), .B1(new_n635), .B2(KEYINPUT16), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n414), .B1(new_n636), .B2(new_n410), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n422), .A2(new_n423), .ZN(new_n638));
  OAI21_X1  g0438(.A(KEYINPUT91), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT91), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n424), .A2(new_n425), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n427), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n639), .A2(KEYINPUT18), .A3(new_n641), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n629), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n299), .A2(new_n305), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n290), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n627), .A2(new_n648), .ZN(G369));
  INV_X1    g0449(.A(new_n605), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n251), .A2(G13), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n266), .A2(new_n651), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(G213), .A3(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(G343), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n658), .A2(new_n597), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n659), .B(KEYINPUT92), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n650), .A2(new_n617), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(new_n650), .B2(new_n660), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(G330), .ZN(new_n663));
  INV_X1    g0463(.A(new_n606), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n573), .B1(new_n664), .B2(new_n658), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n557), .A2(new_n562), .B1(new_n610), .B2(new_n612), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n666), .A2(new_n658), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n663), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n669), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n650), .A2(new_n657), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n673), .B1(new_n668), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n672), .A2(new_n675), .ZN(G399));
  NOR2_X1   g0476(.A1(new_n507), .A2(G116), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n207), .A2(new_n282), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(G1), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n211), .B2(new_n678), .ZN(new_n680));
  XOR2_X1   g0480(.A(new_n680), .B(KEYINPUT93), .Z(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT28), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT94), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT30), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n525), .A2(new_n569), .A3(new_n567), .A4(new_n519), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n685), .A2(new_n603), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n683), .B(new_n684), .C1(new_n686), .C2(new_n487), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n685), .A2(new_n603), .A3(new_n487), .ZN(new_n688));
  OAI21_X1  g0488(.A(KEYINPUT30), .B1(new_n688), .B2(KEYINPUT94), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n615), .A2(G179), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n525), .A2(new_n519), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n690), .A2(new_n570), .A3(new_n487), .A4(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n687), .A2(new_n689), .A3(new_n692), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n693), .A2(KEYINPUT31), .A3(new_n657), .ZN(new_n694));
  AOI21_X1  g0494(.A(KEYINPUT31), .B1(new_n693), .B2(new_n657), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n575), .A2(new_n614), .A3(new_n617), .A4(new_n658), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(G330), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OAI211_X1 g0501(.A(new_n573), .B(new_n533), .C1(new_n666), .C2(new_n605), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n657), .B1(new_n702), .B2(new_n625), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT29), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n682), .B1(new_n707), .B2(new_n284), .ZN(new_n708));
  XOR2_X1   g0508(.A(new_n708), .B(KEYINPUT95), .Z(G364));
  INV_X1    g0509(.A(new_n663), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n284), .B1(new_n651), .B2(G45), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n678), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(G330), .B2(new_n662), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n270), .A2(new_n207), .ZN(new_n716));
  INV_X1    g0516(.A(G355), .ZN(new_n717));
  OAI22_X1  g0517(.A1(new_n716), .A2(new_n717), .B1(G116), .B2(new_n207), .ZN(new_n718));
  XOR2_X1   g0518(.A(new_n718), .B(KEYINPUT96), .Z(new_n719));
  OR2_X1    g0519(.A1(new_n240), .A2(new_n516), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n394), .A2(new_n395), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n207), .ZN(new_n722));
  INV_X1    g0522(.A(new_n211), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n722), .B1(new_n516), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n719), .B1(new_n720), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(G13), .A2(G33), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(G20), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n255), .B1(G20), .B2(new_n287), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n713), .B1(new_n725), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n251), .A2(new_n356), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n733), .A2(new_n291), .A3(G200), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(G317), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(KEYINPUT33), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n736), .A2(KEYINPUT33), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n735), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(G294), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n291), .A2(G179), .A3(G200), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n251), .ZN(new_n742));
  INV_X1    g0542(.A(G303), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n251), .A2(new_n353), .A3(G179), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G190), .ZN(new_n745));
  OAI221_X1 g0545(.A(new_n739), .B1(new_n740), .B2(new_n742), .C1(new_n743), .C2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G190), .A2(G200), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n747), .A2(G20), .A3(new_n356), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n270), .B1(new_n749), .B2(G329), .ZN(new_n750));
  NOR4_X1   g0550(.A1(new_n251), .A2(new_n356), .A3(new_n291), .A4(G200), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(G322), .ZN(new_n753));
  INV_X1    g0553(.A(G311), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n733), .A2(new_n747), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI221_X1 g0556(.A(new_n750), .B1(new_n752), .B2(new_n753), .C1(new_n754), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n744), .A2(new_n291), .ZN(new_n758));
  INV_X1    g0558(.A(G283), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n733), .A2(G190), .A3(G200), .ZN(new_n760));
  INV_X1    g0560(.A(G326), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n758), .A2(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n746), .A2(new_n757), .A3(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n270), .B1(new_n756), .B2(new_n218), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n745), .A2(new_n214), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT32), .ZN(new_n766));
  INV_X1    g0566(.A(G159), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n748), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n765), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n742), .ZN(new_n770));
  INV_X1    g0570(.A(new_n760), .ZN(new_n771));
  AOI22_X1  g0571(.A1(G97), .A2(new_n770), .B1(new_n771), .B2(G50), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n764), .B(new_n773), .C1(G58), .C2(new_n751), .ZN(new_n774));
  INV_X1    g0574(.A(new_n758), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n775), .A2(G107), .B1(new_n735), .B2(G68), .ZN(new_n776));
  OAI211_X1 g0576(.A(new_n774), .B(new_n776), .C1(new_n766), .C2(new_n768), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT97), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n763), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(new_n778), .B2(new_n777), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n732), .B1(new_n780), .B2(new_n729), .ZN(new_n781));
  INV_X1    g0581(.A(new_n728), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n781), .B1(new_n662), .B2(new_n782), .ZN(new_n783));
  AND2_X1   g0583(.A1(new_n715), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(G396));
  NOR2_X1   g0585(.A1(new_n358), .A2(new_n657), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n345), .A2(new_n657), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n354), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n786), .B1(new_n788), .B2(new_n358), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n626), .A2(new_n658), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(KEYINPUT98), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n703), .A2(new_n789), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n791), .B(new_n792), .Z(new_n793));
  INV_X1    g0593(.A(new_n701), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n795), .B(new_n796), .C1(new_n678), .C2(new_n711), .ZN(new_n797));
  INV_X1    g0597(.A(new_n789), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(new_n726), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n729), .A2(new_n726), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(G77), .ZN(new_n802));
  AOI22_X1  g0602(.A1(G159), .A2(new_n755), .B1(new_n751), .B2(G143), .ZN(new_n803));
  INV_X1    g0603(.A(G137), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n803), .B1(new_n804), .B2(new_n760), .C1(new_n247), .C2(new_n734), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT34), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n721), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n758), .A2(new_n202), .ZN(new_n809));
  INV_X1    g0609(.A(G132), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n745), .A2(new_n257), .B1(new_n810), .B2(new_n748), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n809), .B(new_n811), .C1(G58), .C2(new_n770), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n807), .A2(new_n808), .A3(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n805), .A2(new_n806), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n775), .A2(G87), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n815), .B1(new_n743), .B2(new_n760), .C1(new_n220), .C2(new_n745), .ZN(new_n816));
  AOI22_X1  g0616(.A1(G97), .A2(new_n770), .B1(new_n735), .B2(G283), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n270), .B1(new_n751), .B2(G294), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n755), .A2(G116), .B1(new_n749), .B2(G311), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n813), .A2(new_n814), .B1(new_n816), .B2(new_n820), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n712), .B(new_n802), .C1(new_n821), .C2(new_n729), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n797), .B1(new_n799), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(G384));
  NOR2_X1   g0624(.A1(new_n210), .A2(new_n552), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT35), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n825), .B1(new_n495), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(new_n826), .B2(new_n495), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT36), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n723), .A2(G77), .A3(new_n387), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n257), .A2(G68), .ZN(new_n831));
  AOI211_X1 g0631(.A(G13), .B(new_n266), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT38), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT101), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n637), .B2(new_n655), .ZN(new_n836));
  INV_X1    g0636(.A(new_n655), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n425), .A2(KEYINPUT101), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(new_n645), .B2(new_n417), .ZN(new_n840));
  AOI21_X1  g0640(.A(KEYINPUT101), .B1(new_n425), .B2(new_n837), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n835), .B(new_n655), .C1(new_n411), .C2(new_n415), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT37), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n426), .A2(new_n416), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n642), .A2(new_n839), .A3(new_n416), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n846), .B1(new_n847), .B2(KEYINPUT37), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n834), .B1(new_n840), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n403), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n402), .B(new_n256), .C1(new_n850), .C2(new_n635), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n655), .B1(new_n851), .B2(new_n415), .ZN(new_n852));
  INV_X1    g0652(.A(new_n430), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT17), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n416), .B(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n852), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n851), .A2(new_n415), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n857), .A2(new_n424), .B1(new_n637), .B2(new_n385), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n852), .B1(new_n858), .B2(KEYINPUT100), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT100), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n385), .A2(new_n411), .A3(new_n415), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n638), .B1(new_n415), .B2(new_n851), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n844), .B1(new_n859), .B2(new_n863), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n856), .B(KEYINPUT38), .C1(new_n864), .C2(new_n846), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT39), .B1(new_n849), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n857), .A2(new_n424), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n868), .A2(KEYINPUT100), .A3(new_n416), .ZN(new_n869));
  INV_X1    g0669(.A(new_n852), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n863), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n846), .B1(new_n871), .B2(KEYINPUT37), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n870), .B1(new_n417), .B2(new_n430), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n834), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n874), .A2(KEYINPUT39), .A3(new_n865), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  OR2_X1    g0676(.A1(new_n333), .A2(new_n657), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n867), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n786), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n790), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n316), .A2(new_n657), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n333), .A2(new_n336), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n882), .B1(new_n333), .B2(new_n336), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n881), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT99), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n881), .A2(KEYINPUT99), .A3(new_n886), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n874), .A2(new_n865), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n643), .A2(new_n644), .A3(new_n655), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n879), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n434), .A2(new_n705), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n895), .A2(new_n648), .ZN(new_n896));
  XOR2_X1   g0696(.A(new_n894), .B(new_n896), .Z(new_n897));
  OAI21_X1  g0697(.A(new_n789), .B1(new_n883), .B2(new_n884), .ZN(new_n898));
  AOI211_X1 g0698(.A(KEYINPUT40), .B(new_n898), .C1(new_n696), .C2(new_n697), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n891), .ZN(new_n900));
  INV_X1    g0700(.A(new_n898), .ZN(new_n901));
  INV_X1    g0701(.A(new_n695), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n693), .A2(KEYINPUT31), .A3(new_n657), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AND4_X1   g0704(.A1(new_n575), .A2(new_n614), .A3(new_n617), .A4(new_n658), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n901), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n906), .B1(new_n865), .B2(new_n849), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT40), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n900), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(new_n434), .A3(new_n698), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n639), .A2(KEYINPUT18), .A3(new_n641), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT18), .B1(new_n639), .B2(new_n641), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n417), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NOR3_X1   g0713(.A1(new_n637), .A2(KEYINPUT91), .A3(new_n638), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n640), .B1(new_n424), .B2(new_n425), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n416), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT37), .B1(new_n916), .B2(new_n843), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n843), .A2(new_n845), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n843), .A2(new_n913), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n865), .B1(new_n919), .B2(KEYINPUT38), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n898), .B1(new_n696), .B2(new_n697), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n922), .A2(KEYINPUT40), .B1(new_n891), .B2(new_n899), .ZN(new_n923));
  INV_X1    g0723(.A(new_n434), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n923), .B1(new_n924), .B2(new_n699), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n910), .A2(new_n925), .A3(G330), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n897), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n266), .B2(new_n651), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n897), .A2(new_n926), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n833), .B1(new_n928), .B2(new_n929), .ZN(G367));
  OR2_X1    g0730(.A1(new_n531), .A2(new_n658), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n931), .A2(new_n527), .A3(new_n532), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT102), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n932), .A2(new_n933), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n931), .A2(new_n527), .ZN(new_n936));
  NOR3_X1   g0736(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT43), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n674), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n670), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT42), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n494), .B(new_n500), .C1(new_n497), .C2(new_n658), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n623), .A2(new_n657), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n941), .A2(new_n942), .A3(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT103), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n946), .B(new_n947), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n667), .A2(new_n943), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n657), .B1(new_n949), .B2(new_n494), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n941), .A2(new_n945), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n950), .B1(new_n951), .B2(KEYINPUT42), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n939), .B1(new_n948), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n937), .A2(new_n938), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n671), .A2(new_n945), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n953), .A2(new_n954), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n956), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n959), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n957), .B1(new_n961), .B2(new_n955), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n678), .B(KEYINPUT41), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n673), .B1(new_n667), .B2(new_n665), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n674), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n670), .A2(new_n940), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n663), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AND3_X1   g0767(.A1(new_n965), .A2(new_n663), .A3(new_n966), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n706), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n675), .A2(new_n945), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(KEYINPUT104), .B2(KEYINPUT44), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT104), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT44), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n972), .B(new_n973), .C1(new_n675), .C2(new_n945), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n971), .B(new_n974), .C1(new_n972), .C2(new_n973), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n675), .A2(new_n945), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT45), .Z(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n671), .A2(KEYINPUT105), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n969), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n975), .A2(new_n977), .A3(new_n979), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n963), .B1(new_n983), .B2(new_n706), .ZN(new_n984));
  INV_X1    g0784(.A(new_n711), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n960), .B(new_n962), .C1(new_n984), .C2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n937), .A2(new_n728), .ZN(new_n987));
  INV_X1    g0787(.A(new_n745), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(G116), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT46), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n721), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n775), .A2(G97), .B1(new_n771), .B2(G311), .ZN(new_n992));
  AOI22_X1  g0792(.A1(G107), .A2(new_n770), .B1(new_n735), .B2(G294), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n755), .A2(G283), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n751), .A2(new_n581), .B1(new_n749), .B2(G317), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n992), .A2(new_n993), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n775), .A2(G77), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n997), .B1(new_n767), .B2(new_n734), .C1(new_n201), .C2(new_n745), .ZN(new_n998));
  AOI22_X1  g0798(.A1(G68), .A2(new_n770), .B1(new_n771), .B2(G143), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n407), .B1(new_n749), .B2(G137), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(G50), .A2(new_n755), .B1(new_n751), .B2(G150), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n991), .A2(new_n996), .B1(new_n998), .B2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(KEYINPUT106), .B(KEYINPUT47), .Z(new_n1004));
  XNOR2_X1  g0804(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n729), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n730), .B1(new_n207), .B2(new_n341), .C1(new_n230), .C2(new_n722), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n987), .A2(new_n713), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n986), .A2(new_n1008), .ZN(G387));
  NOR2_X1   g0809(.A1(new_n968), .A2(new_n967), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n707), .A2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n678), .B(KEYINPUT109), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1011), .A2(new_n969), .A3(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n964), .A2(new_n782), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n716), .A2(new_n677), .B1(G107), .B2(new_n207), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n235), .A2(new_n516), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n677), .ZN(new_n1017));
  AOI211_X1 g0817(.A(G45), .B(new_n1017), .C1(G68), .C2(G77), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n250), .A2(G50), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT50), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n722), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1015), .B1(new_n1016), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n770), .A2(new_n501), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n734), .B2(new_n250), .C1(new_n767), .C2(new_n760), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n755), .A2(G68), .B1(new_n749), .B2(G150), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n257), .B2(new_n752), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n218), .A2(new_n745), .B1(new_n758), .B2(new_n457), .ZN(new_n1027));
  NOR4_X1   g0827(.A1(new_n1024), .A2(new_n1026), .A3(new_n721), .A4(new_n1027), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n758), .A2(new_n552), .B1(new_n761), .B2(new_n748), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n745), .A2(new_n740), .B1(new_n742), .B2(new_n759), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n581), .A2(new_n755), .B1(new_n751), .B2(G317), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n1031), .B1(new_n754), .B2(new_n734), .C1(new_n753), .C2(new_n760), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT48), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1030), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n1033), .B2(new_n1032), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT107), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n808), .B(new_n1029), .C1(new_n1036), .C2(KEYINPUT49), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1036), .A2(KEYINPUT49), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1028), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n729), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n713), .B1(new_n731), .B2(new_n1022), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT108), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1013), .B1(new_n711), .B2(new_n1010), .C1(new_n1014), .C2(new_n1042), .ZN(G393));
  NOR2_X1   g0843(.A1(new_n978), .A2(new_n671), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n672), .B1(new_n975), .B2(new_n977), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n969), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1046), .A2(new_n983), .A3(new_n1012), .ZN(new_n1047));
  OR3_X1    g0847(.A1(new_n1044), .A2(new_n711), .A3(new_n1045), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n730), .B1(new_n457), .B2(new_n207), .C1(new_n244), .C2(new_n722), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n713), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n771), .A2(G150), .B1(new_n751), .B2(G159), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT110), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n1052), .A2(KEYINPUT51), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(KEYINPUT51), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n988), .A2(G68), .B1(new_n735), .B2(G50), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n755), .A2(new_n339), .B1(new_n749), .B2(G143), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n770), .A2(G77), .ZN(new_n1057));
  AND4_X1   g0857(.A1(new_n815), .A2(new_n1055), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1053), .A2(new_n808), .A3(new_n1054), .A4(new_n1058), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n771), .A2(G317), .B1(new_n751), .B2(G311), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT52), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n988), .A2(G283), .B1(new_n770), .B2(G116), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n775), .A2(G107), .B1(new_n735), .B2(new_n581), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n407), .B1(new_n748), .B2(new_n753), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(G294), .B2(new_n755), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1062), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1059), .B1(new_n1061), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1050), .B1(new_n1067), .B2(new_n729), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n945), .B2(new_n782), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1047), .A2(new_n1048), .A3(new_n1069), .ZN(G390));
  INV_X1    g0870(.A(KEYINPUT113), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n698), .A2(G330), .A3(new_n789), .A4(new_n886), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n786), .B1(new_n703), .B2(new_n789), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n877), .B1(new_n1073), .B2(new_n885), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n866), .B2(new_n875), .ZN(new_n1075));
  AND4_X1   g0875(.A1(KEYINPUT111), .A2(new_n887), .A3(new_n877), .A4(new_n920), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n878), .B1(new_n881), .B2(new_n886), .ZN(new_n1077));
  AOI21_X1  g0877(.A(KEYINPUT111), .B1(new_n1077), .B2(new_n920), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1072), .B(new_n1075), .C1(new_n1076), .C2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT111), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n913), .A2(new_n843), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n917), .A2(new_n918), .ZN(new_n1083));
  AOI21_X1  g0883(.A(KEYINPUT38), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NOR3_X1   g0884(.A1(new_n872), .A2(new_n834), .A3(new_n873), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1081), .B1(new_n1074), .B2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1077), .A2(KEYINPUT111), .A3(new_n920), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1072), .B1(new_n1089), .B2(new_n1075), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1071), .B1(new_n1080), .B2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1075), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1072), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1094), .A2(KEYINPUT113), .A3(new_n1079), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT112), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1072), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n1073), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n698), .A2(G330), .A3(new_n789), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n885), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n1072), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1100), .A2(KEYINPUT112), .A3(new_n1073), .A4(new_n1072), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n701), .A2(new_n434), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1105), .A2(new_n895), .A3(new_n648), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1104), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1091), .A2(new_n1095), .A3(new_n1108), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1094), .A2(new_n1079), .A3(new_n1104), .A4(new_n1107), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT114), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1109), .A2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1091), .A2(new_n1095), .A3(new_n1111), .A4(new_n1108), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1113), .A2(new_n1012), .A3(new_n1114), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1057), .B1(new_n734), .B2(new_n220), .C1(new_n759), .C2(new_n760), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n751), .A2(G116), .B1(new_n749), .B2(G294), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1117), .B(new_n407), .C1(new_n457), .C2(new_n756), .ZN(new_n1118));
  NOR4_X1   g0918(.A1(new_n1116), .A2(new_n1118), .A3(new_n765), .A4(new_n809), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n771), .A2(G128), .B1(new_n751), .B2(G132), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT117), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n745), .A2(new_n247), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT53), .ZN(new_n1123));
  INV_X1    g0923(.A(G125), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n1122), .A2(new_n1123), .B1(new_n1124), .B2(new_n748), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(new_n1123), .B2(new_n1122), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n270), .B1(new_n758), .B2(new_n257), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT116), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n1121), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(KEYINPUT54), .B(G143), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n770), .A2(G159), .B1(new_n755), .B2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n804), .B2(new_n734), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT115), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1119), .B1(new_n1129), .B2(new_n1134), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n713), .B1(new_n339), .B2(new_n801), .C1(new_n1135), .C2(new_n1040), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n867), .A2(new_n876), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1136), .B1(new_n1137), .B2(new_n726), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1080), .A2(new_n1090), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1138), .B1(new_n1139), .B2(new_n985), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1115), .A2(new_n1140), .ZN(G378));
  INV_X1    g0941(.A(KEYINPUT120), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n923), .B2(new_n700), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n900), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n908), .B1(new_n920), .B2(new_n921), .ZN(new_n1145));
  OAI211_X1 g0945(.A(KEYINPUT120), .B(G330), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n269), .A2(new_n837), .ZN(new_n1147));
  XOR2_X1   g0947(.A(new_n306), .B(new_n1147), .Z(new_n1148));
  XNOR2_X1  g0948(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1149));
  XOR2_X1   g0949(.A(new_n1148), .B(new_n1149), .Z(new_n1150));
  NAND3_X1  g0950(.A1(new_n1143), .A2(new_n1146), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n894), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1150), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1142), .B(new_n1153), .C1(new_n923), .C2(new_n700), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n1151), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1152), .B1(new_n1151), .B2(new_n1154), .ZN(new_n1156));
  NOR3_X1   g0956(.A1(new_n1155), .A2(new_n1156), .A3(new_n711), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1150), .A2(new_n726), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n713), .B1(new_n801), .B2(G50), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n756), .A2(new_n804), .B1(new_n810), .B2(new_n734), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT119), .ZN(new_n1161));
  INV_X1    g0961(.A(G128), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n752), .A2(new_n1162), .B1(new_n247), .B2(new_n742), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n745), .A2(new_n1130), .B1(new_n760), .B2(new_n1124), .ZN(new_n1164));
  NOR3_X1   g0964(.A1(new_n1161), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  OR2_X1    g0966(.A1(new_n1166), .A2(KEYINPUT59), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(KEYINPUT59), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n775), .A2(G159), .ZN(new_n1169));
  AOI211_X1 g0969(.A(G33), .B(G41), .C1(new_n749), .C2(G124), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n758), .A2(new_n201), .ZN(new_n1172));
  XOR2_X1   g0972(.A(new_n1172), .B(KEYINPUT118), .Z(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n721), .ZN(new_n1174));
  AOI21_X1  g0974(.A(G41), .B1(new_n749), .B2(G283), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1175), .B1(new_n752), .B2(new_n220), .C1(new_n341), .C2(new_n756), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(G97), .A2(new_n735), .B1(new_n771), .B2(G116), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1177), .B1(new_n202), .B2(new_n742), .C1(new_n218), .C2(new_n745), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n1174), .A2(new_n1176), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(KEYINPUT58), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n282), .B1(new_n721), .B2(new_n281), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n257), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n1179), .A2(KEYINPUT58), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1171), .A2(new_n1180), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1159), .B1(new_n1184), .B2(new_n729), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1158), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(KEYINPUT121), .B1(new_n1157), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n894), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1151), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1190), .A2(new_n985), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT121), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1192), .A2(new_n1193), .A3(new_n1186), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1188), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1110), .A2(new_n1107), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1196), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT57), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1196), .A2(new_n1190), .A3(KEYINPUT57), .A4(new_n1191), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1199), .A2(new_n1012), .A3(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1195), .A2(new_n1201), .ZN(G375));
  INV_X1    g1002(.A(new_n963), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1102), .A2(new_n1103), .A3(new_n1106), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1108), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n885), .A2(new_n726), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n713), .B1(new_n801), .B2(G68), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n220), .A2(new_n756), .B1(new_n752), .B2(new_n759), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n270), .B(new_n1208), .C1(G303), .C2(new_n749), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n734), .A2(new_n552), .B1(new_n760), .B2(new_n740), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(G97), .B2(new_n988), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1209), .A2(new_n997), .A3(new_n1023), .A4(new_n1211), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n756), .A2(new_n247), .B1(new_n748), .B2(new_n1162), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(G137), .B2(new_n751), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n988), .A2(G159), .B1(new_n735), .B2(new_n1131), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(G50), .A2(new_n770), .B1(new_n771), .B2(G132), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1173), .A2(new_n808), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1212), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1207), .B1(new_n1219), .B2(new_n729), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n1104), .A2(new_n985), .B1(new_n1206), .B2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1205), .A2(new_n1221), .ZN(G381));
  INV_X1    g1022(.A(KEYINPUT122), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(new_n1115), .B2(new_n1140), .ZN(new_n1224));
  AND3_X1   g1024(.A1(new_n1115), .A2(new_n1223), .A3(new_n1140), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(G375), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  OR2_X1    g1026(.A1(G393), .A2(G396), .ZN(new_n1227));
  NOR4_X1   g1027(.A1(G384), .A2(new_n1227), .A3(G390), .A4(G381), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1226), .A2(new_n986), .A3(new_n1008), .A4(new_n1228), .ZN(G407));
  NAND3_X1  g1029(.A1(new_n1226), .A2(G213), .A3(new_n656), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(G407), .A2(G213), .A3(new_n1230), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1231), .B(KEYINPUT123), .ZN(G409));
  NAND2_X1  g1032(.A1(new_n656), .A2(G213), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT60), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1012), .B1(new_n1204), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1204), .A2(new_n1234), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n1108), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(KEYINPUT124), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT124), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1236), .A2(new_n1108), .A3(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1235), .B1(new_n1238), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1221), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n823), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NOR3_X1   g1044(.A1(new_n1241), .A2(new_n823), .A3(new_n1242), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1196), .A2(new_n1190), .A3(new_n1203), .A4(new_n1191), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1247), .A2(new_n1192), .A3(new_n1186), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1225), .A2(new_n1224), .A3(new_n1249), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1195), .A2(G378), .A3(new_n1201), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1233), .B(new_n1246), .C1(new_n1250), .C2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(KEYINPUT62), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1233), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1254));
  INV_X1    g1054(.A(G2897), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1233), .A2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1246), .A2(new_n1256), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n1244), .A2(new_n1245), .B1(new_n1255), .B2(new_n1233), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1254), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT61), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(G378), .A2(KEYINPUT122), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1115), .A2(new_n1223), .A3(new_n1140), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1262), .A2(new_n1248), .A3(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1195), .A2(G378), .A3(new_n1201), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT62), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1266), .A2(new_n1267), .A3(new_n1233), .A4(new_n1246), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1253), .A2(new_n1260), .A3(new_n1261), .A4(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(G390), .B1(new_n986), .B2(new_n1008), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(G393), .A2(G396), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n986), .A2(new_n1008), .A3(G390), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1271), .A2(new_n1227), .A3(new_n1272), .A4(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1227), .A2(new_n1272), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1273), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1275), .B1(new_n1276), .B2(new_n1270), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1274), .A2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1269), .A2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1274), .A2(new_n1277), .A3(new_n1261), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT63), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1280), .B1(new_n1252), .B2(new_n1281), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1266), .A2(KEYINPUT63), .A3(new_n1233), .A4(new_n1246), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT125), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1259), .B1(new_n1254), .B2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT125), .B1(new_n1266), .B2(new_n1233), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1282), .B(new_n1283), .C1(new_n1285), .C2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1279), .A2(new_n1287), .ZN(G405));
  OR3_X1    g1088(.A1(new_n1244), .A2(KEYINPUT127), .A3(new_n1245), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(new_n1278), .B(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(G375), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1292));
  OR2_X1    g1092(.A1(new_n1292), .A2(KEYINPUT126), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(KEYINPUT126), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1293), .A2(new_n1265), .A3(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1291), .A2(new_n1295), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1290), .A2(new_n1265), .A3(new_n1294), .A4(new_n1293), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(G402));
endmodule


