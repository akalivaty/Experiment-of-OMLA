//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1 1 0 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 1 1 1 0 1 0 0 1 0 0 0 0 1 1 1 0 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1241, new_n1242, new_n1243,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XNOR2_X1  g0005(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n205), .B(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(G68), .ZN(new_n208));
  INV_X1    g0008(.A(G238), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G87), .ZN(new_n211));
  INV_X1    g0011(.A(G250), .ZN(new_n212));
  INV_X1    g0012(.A(G97), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  OAI22_X1  g0014(.A1(new_n211), .A2(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n210), .B(new_n215), .C1(G107), .C2(G264), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G50), .A2(G226), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G77), .A2(G244), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G116), .A2(G270), .ZN(new_n219));
  NAND4_X1  g0019(.A1(new_n216), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G58), .ZN(new_n221));
  INV_X1    g0021(.A(G232), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n203), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n221), .A2(new_n208), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G50), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n207), .B(new_n225), .C1(new_n228), .C2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G264), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n235), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  INV_X1    g0043(.A(G107), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(G97), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n213), .A2(G107), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n243), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(KEYINPUT7), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT3), .B(G33), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n251), .B1(new_n252), .B2(G20), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(KEYINPUT7), .A3(new_n227), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n253), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G68), .ZN(new_n261));
  AND3_X1   g0061(.A1(new_n227), .A2(new_n254), .A3(KEYINPUT66), .ZN(new_n262));
  AOI21_X1  g0062(.A(KEYINPUT66), .B1(new_n227), .B2(new_n254), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G159), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G58), .A2(G68), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n227), .B1(new_n229), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n261), .A2(new_n267), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT16), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n226), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n261), .A2(KEYINPUT16), .A3(new_n267), .A4(new_n270), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n273), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G1698), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT65), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT65), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G1698), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n282), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n283));
  OAI22_X1  g0083(.A1(new_n283), .A2(new_n258), .B1(new_n254), .B2(new_n211), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G33), .A2(G41), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(G1), .A3(G13), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G1), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n289), .B1(G41), .B2(G45), .ZN(new_n290));
  INV_X1    g0090(.A(G274), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n286), .A2(new_n290), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G232), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n288), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G200), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n288), .A2(G190), .A3(new_n293), .A4(new_n295), .ZN(new_n298));
  XNOR2_X1  g0098(.A(KEYINPUT8), .B(G58), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n227), .A2(G1), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n289), .A2(G13), .A3(G20), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n303), .A2(new_n275), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n301), .A2(new_n304), .B1(new_n303), .B2(new_n299), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n277), .A2(new_n297), .A3(new_n298), .A4(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT17), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n305), .ZN(new_n309));
  INV_X1    g0109(.A(new_n275), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n310), .B1(new_n271), .B2(new_n272), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n309), .B1(new_n311), .B2(new_n276), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n312), .A2(KEYINPUT17), .A3(new_n297), .A4(new_n298), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n308), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(G33), .A2(G97), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT69), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n315), .B(new_n316), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT65), .B(G1698), .ZN(new_n318));
  INV_X1    g0118(.A(G226), .ZN(new_n319));
  OAI22_X1  g0119(.A1(new_n318), .A2(new_n319), .B1(new_n222), .B2(new_n278), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n317), .B1(new_n320), .B2(new_n252), .ZN(new_n321));
  OR2_X1    g0121(.A1(new_n321), .A2(new_n286), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n292), .B1(new_n294), .B2(G238), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT70), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n322), .A2(new_n323), .B1(new_n324), .B2(KEYINPUT13), .ZN(new_n325));
  OAI211_X1 g0125(.A(KEYINPUT13), .B(new_n323), .C1(new_n321), .C2(new_n286), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n326), .A2(KEYINPUT70), .ZN(new_n327));
  OAI21_X1  g0127(.A(G190), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n303), .A2(KEYINPUT12), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n302), .A2(KEYINPUT68), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT68), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n331), .A2(new_n289), .A3(G13), .A4(G20), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n310), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(KEYINPUT12), .B1(new_n333), .B2(new_n300), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n329), .B1(new_n334), .B2(G68), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n330), .A2(new_n332), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(KEYINPUT12), .A3(new_n208), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n208), .A2(G20), .ZN(new_n338));
  INV_X1    g0138(.A(G77), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n254), .A2(G20), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G50), .ZN(new_n342));
  OAI221_X1 g0142(.A(new_n338), .B1(new_n339), .B2(new_n341), .C1(new_n264), .C2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT11), .ZN(new_n344));
  AND3_X1   g0144(.A1(new_n343), .A2(new_n344), .A3(new_n275), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n344), .B1(new_n343), .B2(new_n275), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n335), .B(new_n337), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT13), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n321), .A2(new_n286), .ZN(new_n350));
  INV_X1    g0150(.A(new_n323), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n349), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n352), .A2(G200), .A3(new_n326), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n328), .A2(new_n348), .A3(KEYINPUT71), .A4(new_n353), .ZN(new_n354));
  XOR2_X1   g0154(.A(KEYINPUT15), .B(G87), .Z(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n340), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT67), .ZN(new_n357));
  XNOR2_X1  g0157(.A(new_n356), .B(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n264), .ZN(new_n359));
  INV_X1    g0159(.A(new_n299), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(G20), .A2(G77), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n358), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n275), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n336), .A2(new_n339), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n333), .A2(new_n300), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(G77), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n364), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  OAI221_X1 g0168(.A(new_n252), .B1(new_n209), .B2(new_n278), .C1(new_n318), .C2(new_n222), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n369), .B(new_n287), .C1(G107), .C2(new_n252), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n294), .A2(G244), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(new_n293), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(G169), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OR2_X1    g0174(.A1(new_n372), .A2(G179), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n368), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  AND2_X1   g0176(.A1(new_n354), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n208), .B1(new_n253), .B2(new_n259), .ZN(new_n378));
  NOR3_X1   g0178(.A1(new_n378), .A2(new_n266), .A3(new_n269), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n275), .B1(new_n379), .B2(KEYINPUT16), .ZN(new_n380));
  INV_X1    g0180(.A(new_n276), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n305), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n296), .A2(G169), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n288), .A2(G179), .A3(new_n293), .A4(new_n295), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(KEYINPUT18), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n382), .A2(new_n385), .A3(KEYINPUT18), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(G190), .ZN(new_n390));
  OR2_X1    g0190(.A1(new_n372), .A2(new_n390), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n363), .A2(new_n275), .B1(G77), .B2(new_n366), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n372), .A2(G200), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n391), .A2(new_n392), .A3(new_n393), .A4(new_n365), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n314), .A2(new_n377), .A3(new_n389), .A4(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n352), .A2(G169), .A3(new_n326), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT14), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n397), .A2(KEYINPUT72), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(G179), .B1(new_n325), .B2(new_n327), .ZN(new_n400));
  INV_X1    g0200(.A(new_n398), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n352), .A2(G169), .A3(new_n326), .A4(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n399), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  AND2_X1   g0203(.A1(new_n403), .A2(new_n347), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n395), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G223), .A2(G1698), .ZN(new_n406));
  INV_X1    g0206(.A(G222), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n252), .B(new_n406), .C1(new_n318), .C2(new_n407), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n408), .B(new_n287), .C1(G77), .C2(new_n252), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n294), .A2(G226), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n409), .A2(new_n410), .A3(new_n293), .ZN(new_n411));
  OR2_X1    g0211(.A1(new_n411), .A2(G179), .ZN(new_n412));
  OAI21_X1  g0212(.A(G20), .B1(new_n229), .B2(G50), .ZN(new_n413));
  INV_X1    g0213(.A(G150), .ZN(new_n414));
  OAI221_X1 g0214(.A(new_n413), .B1(new_n299), .B2(new_n341), .C1(new_n264), .C2(new_n414), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n415), .A2(new_n275), .B1(new_n342), .B2(new_n303), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n304), .B(G50), .C1(G1), .C2(new_n227), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n411), .A2(new_n373), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n412), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n411), .A2(G200), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT9), .ZN(new_n423));
  OAI221_X1 g0223(.A(new_n422), .B1(new_n390), .B2(new_n411), .C1(new_n418), .C2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n418), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n425), .A2(KEYINPUT9), .ZN(new_n426));
  OR3_X1    g0226(.A1(new_n424), .A2(KEYINPUT10), .A3(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(KEYINPUT10), .B1(new_n424), .B2(new_n426), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n421), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n328), .A2(new_n353), .A3(new_n348), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT71), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT73), .B1(new_n405), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT73), .ZN(new_n436));
  NOR4_X1   g0236(.A1(new_n433), .A2(new_n395), .A3(new_n436), .A4(new_n404), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT24), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT23), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n227), .B2(G107), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n244), .A2(KEYINPUT23), .A3(G20), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(G116), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n254), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n227), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n255), .A2(new_n257), .A3(new_n227), .A4(G87), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT22), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT22), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n252), .A2(new_n450), .A3(new_n227), .A4(G87), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n447), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT79), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n439), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n449), .A2(new_n451), .ZN(new_n455));
  INV_X1    g0255(.A(new_n447), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT79), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n457), .A2(KEYINPUT79), .A3(new_n439), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n459), .A2(new_n275), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(G13), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n462), .A2(G1), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n463), .A2(G20), .A3(new_n244), .ZN(new_n464));
  XNOR2_X1  g0264(.A(new_n464), .B(KEYINPUT25), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n254), .A2(G1), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n303), .A2(new_n275), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n465), .B1(G107), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n461), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g0269(.A(KEYINPUT5), .B(G41), .ZN(new_n470));
  INV_X1    g0270(.A(G45), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(G1), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n470), .A2(G274), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(G294), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n254), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n214), .A2(new_n278), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n477), .B1(new_n318), .B2(new_n212), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n475), .B1(new_n478), .B2(new_n252), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n473), .B1(new_n479), .B2(new_n286), .ZN(new_n480));
  INV_X1    g0280(.A(G179), .ZN(new_n481));
  AND2_X1   g0281(.A1(KEYINPUT5), .A2(G41), .ZN(new_n482));
  NOR2_X1   g0282(.A1(KEYINPUT5), .A2(G41), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n472), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n484), .A2(G264), .A3(new_n286), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT80), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n484), .A2(KEYINPUT80), .A3(G264), .A4(new_n286), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NOR3_X1   g0289(.A1(new_n480), .A2(new_n481), .A3(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n212), .B1(new_n279), .B2(new_n281), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n252), .B1(new_n492), .B2(new_n476), .ZN(new_n493));
  INV_X1    g0293(.A(new_n475), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n286), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n473), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n489), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G169), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n491), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n469), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n333), .A2(G116), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n330), .B(new_n332), .C1(new_n444), .C2(new_n466), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G283), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n506), .B(new_n227), .C1(G33), .C2(new_n213), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n444), .A2(G20), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n507), .A2(new_n275), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT20), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n507), .A2(KEYINPUT20), .A3(new_n275), .A4(new_n508), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n505), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G179), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G264), .A2(G1698), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n252), .B(new_n516), .C1(new_n318), .C2(new_n214), .ZN(new_n517));
  INV_X1    g0317(.A(G303), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n286), .B1(new_n258), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n226), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n470), .A2(new_n472), .B1(new_n521), .B2(new_n285), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G270), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n520), .A2(new_n523), .A3(new_n473), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n515), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n373), .B1(new_n505), .B2(new_n513), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT78), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n519), .A2(new_n517), .B1(new_n522), .B2(G270), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n529), .A2(KEYINPUT78), .A3(new_n473), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n526), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(KEYINPUT21), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT21), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n526), .A2(new_n528), .A3(new_n530), .A4(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n525), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(KEYINPUT78), .B1(new_n529), .B2(new_n473), .ZN(new_n536));
  AND4_X1   g0336(.A1(KEYINPUT78), .A2(new_n520), .A3(new_n523), .A4(new_n473), .ZN(new_n537));
  OAI21_X1  g0337(.A(G190), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n514), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n528), .A2(new_n530), .A3(G200), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n502), .A2(new_n535), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n282), .A2(new_n252), .A3(G244), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT4), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n255), .A2(new_n257), .A3(G250), .A4(G1698), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n546), .A2(new_n506), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n282), .A2(new_n252), .A3(KEYINPUT4), .A4(G244), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n545), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n287), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n484), .A2(new_n286), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n473), .B1(new_n551), .B2(new_n214), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n550), .A2(G190), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(G200), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n552), .B1(new_n549), .B2(new_n287), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n481), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(G169), .B2(new_n556), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n302), .A2(G97), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n467), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n562), .A2(new_n213), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n244), .B1(new_n253), .B2(new_n259), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n264), .A2(new_n339), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT6), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n213), .A2(new_n244), .ZN(new_n568));
  NOR2_X1   g0368(.A1(G97), .A2(G107), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n244), .A2(KEYINPUT6), .A3(G97), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n227), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NOR3_X1   g0372(.A1(new_n565), .A2(new_n566), .A3(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n561), .B(new_n564), .C1(new_n573), .C2(new_n310), .ZN(new_n574));
  MUX2_X1   g0374(.A(new_n557), .B(new_n559), .S(new_n574), .Z(new_n575));
  NAND4_X1  g0375(.A1(new_n255), .A2(new_n257), .A3(G244), .A4(G1698), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(KEYINPUT75), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT75), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n252), .A2(new_n578), .A3(G244), .A4(G1698), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n282), .A2(new_n252), .A3(G238), .ZN(new_n580));
  INV_X1    g0380(.A(new_n445), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n577), .A2(new_n579), .A3(new_n580), .A4(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT76), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n582), .A2(new_n583), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n287), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n472), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n587), .A2(G250), .A3(new_n286), .ZN(new_n588));
  XNOR2_X1  g0388(.A(new_n588), .B(KEYINPUT74), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n472), .A2(G274), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n586), .A2(new_n481), .A3(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n258), .A2(new_n318), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n445), .B1(new_n594), .B2(G238), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n595), .A2(KEYINPUT76), .A3(new_n577), .A4(new_n579), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n582), .A2(new_n583), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n286), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n373), .B1(new_n598), .B2(new_n591), .ZN(new_n599));
  INV_X1    g0399(.A(new_n355), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n336), .ZN(new_n601));
  AOI21_X1  g0401(.A(KEYINPUT19), .B1(new_n340), .B2(G97), .ZN(new_n602));
  NOR3_X1   g0402(.A1(new_n258), .A2(G20), .A3(new_n208), .ZN(new_n603));
  XNOR2_X1  g0403(.A(new_n315), .B(KEYINPUT69), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT19), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n227), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  XNOR2_X1  g0406(.A(KEYINPUT77), .B(G87), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n569), .ZN(new_n608));
  AOI211_X1 g0408(.A(new_n602), .B(new_n603), .C1(new_n606), .C2(new_n608), .ZN(new_n609));
  OAI221_X1 g0409(.A(new_n601), .B1(new_n600), .B2(new_n562), .C1(new_n609), .C2(new_n310), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n593), .A2(new_n599), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n586), .A2(G190), .A3(new_n592), .ZN(new_n612));
  OAI21_X1  g0412(.A(G200), .B1(new_n598), .B2(new_n591), .ZN(new_n613));
  INV_X1    g0413(.A(new_n601), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n562), .A2(new_n211), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n602), .B1(new_n606), .B2(new_n608), .ZN(new_n616));
  INV_X1    g0416(.A(new_n603), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI211_X1 g0418(.A(new_n614), .B(new_n615), .C1(new_n618), .C2(new_n275), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n612), .A2(new_n613), .A3(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n555), .B1(new_n480), .B2(new_n489), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n489), .A2(new_n495), .A3(new_n496), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n621), .A2(KEYINPUT81), .B1(new_n622), .B2(new_n390), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT81), .ZN(new_n624));
  NOR4_X1   g0424(.A1(new_n480), .A2(new_n489), .A3(new_n624), .A4(G190), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n461), .B(new_n468), .C1(new_n623), .C2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n575), .A2(new_n611), .A3(new_n620), .A4(new_n626), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n438), .A2(new_n542), .A3(new_n627), .ZN(G372));
  INV_X1    g0428(.A(new_n376), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n404), .B1(new_n430), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n308), .A2(new_n313), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n389), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n427), .A2(new_n428), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n421), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n502), .A2(new_n535), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n635), .A2(new_n575), .A3(new_n620), .A4(new_n626), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n611), .A2(new_n620), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n550), .A2(new_n553), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n373), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n639), .A2(new_n574), .A3(new_n558), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT26), .B1(new_n637), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(KEYINPUT82), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT82), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n639), .A2(new_n574), .A3(new_n643), .A4(new_n558), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n645), .A2(new_n646), .A3(new_n611), .A4(new_n620), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n636), .A2(new_n641), .A3(new_n647), .A4(new_n611), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n634), .B1(new_n438), .B2(new_n649), .ZN(new_n650));
  XNOR2_X1  g0450(.A(new_n650), .B(KEYINPUT83), .ZN(G369));
  AOI22_X1  g0451(.A1(new_n461), .A2(new_n468), .B1(new_n491), .B2(new_n500), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n463), .A2(new_n227), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(G213), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(G343), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n469), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n652), .B1(new_n626), .B2(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n502), .A2(new_n658), .ZN(new_n661));
  OAI21_X1  g0461(.A(KEYINPUT84), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT84), .ZN(new_n663));
  INV_X1    g0463(.A(new_n658), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n652), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n664), .B1(new_n461), .B2(new_n468), .ZN(new_n666));
  INV_X1    g0466(.A(new_n625), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n624), .B1(new_n499), .B2(new_n555), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n499), .A2(G190), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n469), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n666), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n663), .B(new_n665), .C1(new_n672), .C2(new_n652), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n662), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(G330), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n539), .A2(new_n664), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n535), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n535), .A2(new_n541), .A3(new_n678), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n676), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n675), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n535), .A2(new_n658), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n662), .A2(new_n673), .A3(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n682), .A2(new_n665), .A3(new_n684), .ZN(G399));
  INV_X1    g0485(.A(new_n204), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(G41), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n607), .A2(new_n444), .A3(new_n569), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n688), .A2(G1), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n230), .B2(new_n688), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT28), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n642), .A2(new_n644), .ZN(new_n694));
  OAI21_X1  g0494(.A(KEYINPUT26), .B1(new_n694), .B2(new_n637), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n611), .A2(new_n620), .ZN(new_n696));
  INV_X1    g0496(.A(new_n640), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(new_n646), .A3(new_n697), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n695), .A2(new_n698), .A3(new_n611), .A4(new_n636), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n664), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(KEYINPUT29), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT29), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n648), .A2(new_n702), .A3(new_n664), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n542), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n640), .B1(new_n574), .B2(new_n557), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n706), .B1(new_n671), .B2(new_n670), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n705), .A2(new_n707), .A3(new_n696), .A4(new_n664), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT31), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n586), .A2(new_n592), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n556), .A2(new_n536), .A3(new_n537), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n710), .A2(new_n711), .A3(new_n481), .A4(new_n499), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT30), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n622), .A2(G179), .A3(new_n529), .A4(new_n556), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n713), .B1(new_n710), .B2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n598), .A2(new_n591), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n556), .A2(new_n529), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n716), .A2(KEYINPUT30), .A3(new_n490), .A4(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n712), .A2(new_n715), .A3(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n709), .B1(new_n719), .B2(new_n658), .ZN(new_n720));
  AND3_X1   g0520(.A1(new_n719), .A2(new_n709), .A3(new_n658), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n708), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G330), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(KEYINPUT85), .B1(new_n704), .B2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT85), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n701), .A2(new_n726), .A3(new_n723), .A4(new_n703), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n693), .B1(new_n728), .B2(G1), .ZN(G364));
  AOI21_X1  g0529(.A(new_n226), .B1(G20), .B2(new_n373), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n481), .A2(new_n555), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n227), .A2(G190), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(G317), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(KEYINPUT33), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n735), .A2(KEYINPUT33), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n734), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n555), .A2(G179), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n732), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(G283), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n258), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n227), .A2(new_n390), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n731), .A2(new_n743), .ZN(new_n744));
  XOR2_X1   g0544(.A(new_n744), .B(KEYINPUT90), .Z(new_n745));
  NOR2_X1   g0545(.A1(G179), .A2(G200), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n227), .B1(new_n746), .B2(G190), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  AOI22_X1  g0548(.A1(new_n745), .A2(G326), .B1(G294), .B2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT91), .ZN(new_n750));
  OR2_X1    g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  INV_X1    g0552(.A(G311), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n481), .A2(G200), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n732), .A2(new_n754), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n751), .B(new_n752), .C1(new_n753), .C2(new_n755), .ZN(new_n756));
  XOR2_X1   g0556(.A(new_n756), .B(KEYINPUT92), .Z(new_n757));
  NAND2_X1  g0557(.A1(new_n732), .A2(new_n746), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI211_X1 g0559(.A(new_n742), .B(new_n757), .C1(G329), .C2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n743), .A2(new_n739), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G303), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n743), .A2(new_n754), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G322), .ZN(new_n766));
  AND4_X1   g0566(.A1(new_n738), .A2(new_n760), .A3(new_n763), .A4(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n747), .A2(new_n213), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  XOR2_X1   g0569(.A(new_n764), .B(KEYINPUT89), .Z(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  OAI221_X1 g0571(.A(new_n769), .B1(new_n607), .B2(new_n761), .C1(new_n771), .C2(new_n221), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n733), .A2(new_n208), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n740), .A2(new_n244), .ZN(new_n774));
  INV_X1    g0574(.A(new_n755), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n774), .B1(G77), .B2(new_n775), .ZN(new_n776));
  OAI211_X1 g0576(.A(new_n776), .B(new_n252), .C1(new_n342), .C2(new_n744), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n759), .A2(G159), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT32), .ZN(new_n779));
  NOR4_X1   g0579(.A1(new_n772), .A2(new_n773), .A3(new_n777), .A4(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n730), .B1(new_n767), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G13), .A2(G33), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT87), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(new_n227), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT88), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n730), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n231), .A2(new_n471), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n686), .A2(new_n252), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n788), .B(new_n789), .C1(new_n243), .C2(new_n471), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n252), .A2(G355), .A3(new_n204), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n790), .B(new_n791), .C1(G116), .C2(new_n204), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n787), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n462), .A2(G20), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G45), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n795), .A2(KEYINPUT86), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(KEYINPUT86), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n796), .A2(G1), .A3(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n687), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n679), .A2(new_n680), .A3(new_n786), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n781), .A2(new_n793), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n681), .ZN(new_n802));
  INV_X1    g0602(.A(new_n799), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n679), .A2(new_n676), .A3(new_n680), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n801), .A2(new_n805), .ZN(G396));
  INV_X1    g0606(.A(new_n744), .ZN(new_n807));
  AOI22_X1  g0607(.A1(G137), .A2(new_n807), .B1(new_n734), .B2(G150), .ZN(new_n808));
  INV_X1    g0608(.A(G143), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n808), .B1(new_n265), .B2(new_n755), .C1(new_n771), .C2(new_n809), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT34), .Z(new_n811));
  AOI21_X1  g0611(.A(new_n258), .B1(new_n759), .B2(G132), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(KEYINPUT93), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n740), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n812), .A2(KEYINPUT93), .B1(G68), .B2(new_n815), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n814), .B(new_n816), .C1(new_n342), .C2(new_n761), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(G58), .B2(new_n748), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n740), .A2(new_n211), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n769), .B1(new_n244), .B2(new_n761), .C1(new_n518), .C2(new_n744), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n819), .B(new_n820), .C1(G311), .C2(new_n759), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n252), .B1(new_n775), .B2(G116), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n821), .B(new_n822), .C1(new_n741), .C2(new_n733), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(G294), .B2(new_n765), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n730), .B1(new_n818), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n783), .A2(new_n730), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n339), .ZN(new_n827));
  AND4_X1   g0627(.A1(new_n368), .A2(new_n374), .A3(new_n375), .A4(new_n664), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n368), .A2(new_n658), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n394), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n828), .B1(new_n376), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n783), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n825), .A2(new_n799), .A3(new_n827), .A4(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n832), .B1(new_n649), .B2(new_n658), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n648), .A2(new_n664), .A3(new_n831), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(new_n723), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n834), .B1(new_n838), .B2(new_n799), .ZN(G384));
  INV_X1    g0639(.A(new_n656), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n382), .B1(new_n385), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT37), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n841), .A2(new_n842), .A3(new_n306), .ZN(new_n843));
  INV_X1    g0643(.A(new_n306), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n271), .A2(KEYINPUT95), .A3(new_n272), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n272), .A2(KEYINPUT95), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n379), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n845), .A2(new_n275), .A3(new_n847), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n848), .A2(new_n305), .B1(new_n383), .B2(new_n384), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n656), .B1(new_n848), .B2(new_n305), .ZN(new_n850));
  NOR3_X1   g0650(.A1(new_n844), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n843), .B1(new_n851), .B2(new_n842), .ZN(new_n852));
  AND3_X1   g0652(.A1(new_n382), .A2(new_n385), .A3(KEYINPUT18), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n853), .A2(new_n386), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n850), .B1(new_n854), .B2(new_n631), .ZN(new_n855));
  AND3_X1   g0655(.A1(new_n852), .A2(KEYINPUT38), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT38), .B1(new_n852), .B2(new_n855), .ZN(new_n857));
  OAI21_X1  g0657(.A(KEYINPUT39), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT38), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n841), .A2(new_n306), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n860), .B(new_n842), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n382), .A2(new_n840), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(new_n314), .B2(new_n389), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n859), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n852), .A2(new_n855), .A3(KEYINPUT38), .ZN(new_n865));
  XNOR2_X1  g0665(.A(KEYINPUT96), .B(KEYINPUT39), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n858), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n404), .A2(new_n664), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n828), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n836), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n403), .A2(new_n658), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n658), .A2(KEYINPUT71), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n399), .A2(new_n400), .A3(new_n402), .A4(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n874), .A2(new_n347), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n430), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n873), .B(new_n879), .C1(new_n857), .C2(new_n856), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n854), .A2(new_n656), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n871), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n704), .B1(new_n435), .B2(new_n437), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n634), .ZN(new_n884));
  XOR2_X1   g0684(.A(new_n882), .B(new_n884), .Z(new_n885));
  INV_X1    g0685(.A(KEYINPUT40), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n856), .A2(new_n857), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n877), .A2(new_n430), .A3(new_n831), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n722), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n886), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n864), .A2(new_n865), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n891), .A2(KEYINPUT40), .A3(new_n722), .A4(new_n888), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n722), .B1(new_n435), .B2(new_n437), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n893), .B(new_n894), .Z(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(G330), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n885), .B(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n289), .B2(new_n794), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n570), .A2(new_n571), .ZN(new_n899));
  OAI211_X1 g0699(.A(G116), .B(new_n228), .C1(new_n899), .C2(KEYINPUT35), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT94), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n899), .A2(KEYINPUT35), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n903), .B(KEYINPUT36), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n268), .A2(G77), .ZN(new_n905));
  OAI22_X1  g0705(.A1(new_n230), .A2(new_n905), .B1(G50), .B2(new_n208), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n906), .A2(G1), .A3(new_n462), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n898), .A2(new_n904), .A3(new_n907), .ZN(G367));
  INV_X1    g0708(.A(new_n574), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n575), .B1(new_n909), .B2(new_n664), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n697), .A2(new_n658), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  OR2_X1    g0713(.A1(new_n684), .A2(new_n913), .ZN(new_n914));
  OR2_X1    g0714(.A1(new_n914), .A2(KEYINPUT42), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n640), .B1(new_n910), .B2(new_n502), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n664), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n914), .A2(KEYINPUT42), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n915), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  OAI221_X1 g0719(.A(new_n601), .B1(new_n211), .B2(new_n562), .C1(new_n609), .C2(new_n310), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n658), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n696), .A2(new_n921), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n922), .B(KEYINPUT97), .Z(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n611), .B2(new_n921), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(KEYINPUT43), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n919), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n682), .A2(new_n913), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n926), .B(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n924), .A2(KEYINPUT43), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT98), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n928), .B(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n687), .B(KEYINPUT41), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n684), .A2(new_n665), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n913), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(KEYINPUT99), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT99), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n934), .A2(new_n937), .A3(new_n913), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n936), .A2(KEYINPUT44), .A3(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT44), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n937), .B1(new_n934), .B2(new_n913), .ZN(new_n941));
  AOI211_X1 g0741(.A(KEYINPUT99), .B(new_n912), .C1(new_n684), .C2(new_n665), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n684), .A2(new_n665), .A3(new_n912), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT45), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n944), .B(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n939), .A2(new_n943), .A3(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n682), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n939), .A2(new_n943), .A3(new_n682), .A4(new_n946), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n674), .A2(new_n802), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n682), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n683), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n682), .A2(new_n683), .A3(new_n951), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(new_n725), .B2(new_n727), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n949), .A2(new_n950), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(KEYINPUT100), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT100), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n949), .A2(new_n957), .A3(new_n960), .A4(new_n950), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n933), .B1(new_n962), .B2(new_n728), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n931), .B1(new_n963), .B2(new_n798), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n764), .A2(new_n414), .B1(new_n740), .B2(new_n339), .ZN(new_n965));
  AOI22_X1  g0765(.A1(G50), .A2(new_n775), .B1(new_n759), .B2(G137), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n221), .B2(new_n761), .ZN(new_n967));
  AOI211_X1 g0767(.A(new_n965), .B(new_n967), .C1(G159), .C2(new_n734), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n748), .A2(G68), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n745), .A2(G143), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n968), .A2(new_n252), .A3(new_n969), .A4(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n771), .A2(new_n518), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n762), .A2(KEYINPUT46), .A3(G116), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n973), .B(new_n258), .C1(new_n244), .C2(new_n747), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n213), .A2(new_n740), .B1(new_n755), .B2(new_n741), .ZN(new_n975));
  AOI21_X1  g0775(.A(KEYINPUT46), .B1(new_n762), .B2(G116), .ZN(new_n976));
  NOR3_X1   g0776(.A1(new_n974), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  AOI22_X1  g0777(.A1(G294), .A2(new_n734), .B1(new_n759), .B2(G317), .ZN(new_n978));
  INV_X1    g0778(.A(new_n745), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n977), .B(new_n978), .C1(new_n753), .C2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n971), .B1(new_n972), .B2(new_n980), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT47), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n730), .ZN(new_n983));
  INV_X1    g0783(.A(new_n789), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n787), .B1(new_n204), .B2(new_n600), .C1(new_n235), .C2(new_n984), .ZN(new_n985));
  AND3_X1   g0785(.A1(new_n983), .A2(new_n799), .A3(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n924), .B2(new_n785), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n964), .A2(new_n987), .ZN(G387));
  AOI21_X1  g0788(.A(new_n803), .B1(new_n674), .B2(new_n786), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n690), .B(new_n471), .C1(new_n208), .C2(new_n339), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT101), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n360), .A2(new_n342), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT50), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n789), .B1(new_n471), .B2(new_n239), .C1(new_n991), .C2(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n689), .A2(new_n204), .A3(new_n252), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n994), .B(new_n995), .C1(G107), .C2(new_n204), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT102), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n787), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n762), .A2(G294), .B1(new_n748), .B2(G283), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n770), .A2(G317), .B1(G311), .B2(new_n734), .ZN(new_n1000));
  INV_X1    g0800(.A(G322), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1000), .B1(new_n518), .B2(new_n755), .C1(new_n1001), .C2(new_n979), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT48), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n999), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT103), .Z(new_n1005));
  NAND2_X1  g0805(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT49), .Z(new_n1008));
  AOI21_X1  g0808(.A(new_n252), .B1(new_n759), .B2(G326), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n444), .B2(new_n740), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n758), .A2(new_n414), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n600), .A2(new_n747), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(G50), .B2(new_n765), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n258), .B1(new_n734), .B2(new_n360), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(G159), .A2(new_n807), .B1(new_n762), .B2(G77), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G68), .A2(new_n775), .B1(new_n815), .B2(G97), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n1008), .A2(new_n1010), .B1(new_n1011), .B2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT104), .Z(new_n1019));
  INV_X1    g0819(.A(new_n730), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n989), .B(new_n998), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n956), .A2(new_n725), .A3(new_n727), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT105), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n688), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n957), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1024), .B(new_n1025), .C1(new_n1023), .C2(new_n1022), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n798), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1021), .B(new_n1026), .C1(new_n1027), .C2(new_n956), .ZN(G393));
  INV_X1    g0828(.A(KEYINPUT109), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n957), .B1(new_n949), .B2(new_n950), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n688), .B(new_n1030), .C1(new_n959), .C2(new_n961), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n949), .A2(new_n798), .A3(new_n950), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n744), .A2(new_n414), .B1(new_n764), .B2(new_n265), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT51), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(G68), .A2(new_n762), .B1(new_n775), .B2(new_n360), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1034), .B(new_n1035), .C1(new_n342), .C2(new_n733), .ZN(new_n1036));
  NOR3_X1   g0836(.A1(new_n1036), .A2(new_n258), .A3(new_n819), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n748), .A2(G77), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1037), .B(new_n1038), .C1(new_n809), .C2(new_n758), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT106), .Z(new_n1040));
  OAI22_X1  g0840(.A1(new_n744), .A2(new_n735), .B1(new_n764), .B2(new_n753), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(KEYINPUT107), .B(KEYINPUT52), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1041), .B(new_n1042), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n252), .B(new_n1043), .C1(G116), .C2(new_n748), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n733), .A2(new_n518), .B1(new_n758), .B2(new_n1001), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1045), .A2(new_n774), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1044), .B(new_n1046), .C1(new_n474), .C2(new_n755), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(G283), .B2(new_n762), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n730), .B1(new_n1040), .B2(new_n1048), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n787), .B1(new_n213), .B2(new_n204), .C1(new_n249), .C2(new_n984), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1049), .A2(new_n799), .A3(new_n1050), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT108), .Z(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n785), .B2(new_n912), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1032), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1029), .B1(new_n1031), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1030), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n962), .A2(new_n1056), .A3(new_n687), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1054), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1057), .A2(KEYINPUT109), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1055), .A2(new_n1059), .ZN(G390));
  NOR2_X1   g0860(.A1(new_n721), .A2(new_n720), .ZN(new_n1061));
  NOR3_X1   g0861(.A1(new_n627), .A2(new_n542), .A3(new_n658), .ZN(new_n1062));
  OAI211_X1 g0862(.A(G330), .B(new_n831), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n878), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT111), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n888), .B(G330), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1063), .A2(KEYINPUT111), .A3(new_n878), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n873), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1067), .A2(KEYINPUT110), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT110), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n722), .A2(new_n1072), .A3(G330), .A4(new_n888), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n830), .A2(new_n376), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n699), .A2(new_n664), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n872), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(new_n878), .B2(new_n1063), .ZN(new_n1078));
  AOI21_X1  g0878(.A(KEYINPUT112), .B1(new_n1074), .B2(new_n1078), .ZN(new_n1079));
  AND4_X1   g0879(.A1(new_n646), .A2(new_n611), .A3(new_n620), .A4(new_n697), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n645), .A2(new_n611), .A3(new_n620), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1080), .B1(KEYINPUT26), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n611), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n920), .B1(new_n716), .B2(G190), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n502), .A2(new_n535), .B1(new_n1084), .B2(new_n613), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1083), .B1(new_n707), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n658), .B1(new_n1082), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n828), .B1(new_n1087), .B2(new_n1075), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1071), .A2(new_n1064), .A3(new_n1073), .A4(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT112), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1070), .B1(new_n1079), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n870), .B1(new_n873), .B2(new_n879), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n878), .B1(new_n1076), .B2(new_n872), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n891), .A2(new_n869), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n1093), .A2(new_n868), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n1067), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n1098), .B1(new_n1095), .B2(new_n1094), .C1(new_n1093), .C2(new_n868), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  OAI211_X1 g0900(.A(G330), .B(new_n722), .C1(new_n435), .C2(new_n437), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n883), .A2(new_n634), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1092), .A2(new_n1100), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n687), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT113), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1100), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1074), .A2(new_n1078), .A3(KEYINPUT112), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1109), .A2(new_n1110), .B1(new_n873), .B2(new_n1069), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT114), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n1111), .A2(new_n1112), .A3(new_n1102), .ZN(new_n1113));
  AOI21_X1  g0913(.A(KEYINPUT114), .B1(new_n1092), .B2(new_n1103), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1108), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1104), .A2(KEYINPUT113), .A3(new_n687), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1107), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1100), .A2(new_n798), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n858), .A2(new_n867), .A3(new_n783), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(G283), .A2(new_n807), .B1(new_n815), .B2(G68), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(new_n211), .B2(new_n761), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n1038), .B1(new_n444), .B2(new_n764), .C1(new_n474), .C2(new_n758), .ZN(new_n1122));
  NOR3_X1   g0922(.A1(new_n1121), .A2(new_n1122), .A3(new_n252), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n1123), .B1(new_n213), .B2(new_n755), .C1(new_n244), .C2(new_n733), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n747), .A2(new_n265), .ZN(new_n1125));
  XOR2_X1   g0925(.A(KEYINPUT54), .B(G143), .Z(new_n1126));
  AOI21_X1  g0926(.A(new_n258), .B1(new_n775), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(G132), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n1127), .B1(new_n342), .B2(new_n740), .C1(new_n1128), .C2(new_n764), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(G125), .B2(new_n759), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n761), .A2(new_n414), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT53), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(G128), .A2(new_n807), .B1(new_n734), .B2(G137), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1130), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1124), .B1(new_n1125), .B2(new_n1134), .ZN(new_n1135));
  XOR2_X1   g0935(.A(new_n1135), .B(KEYINPUT115), .Z(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n730), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n826), .A2(new_n299), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1119), .A2(new_n799), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1118), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1117), .A2(new_n1141), .ZN(G378));
  INV_X1    g0942(.A(KEYINPUT57), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1102), .B(KEYINPUT120), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1102), .B1(new_n1145), .B2(new_n1070), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1144), .B1(new_n1100), .B2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n890), .A2(new_n892), .A3(G330), .ZN(new_n1148));
  XOR2_X1   g0948(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n429), .A2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n429), .A2(new_n1150), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n425), .A2(new_n656), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  OR3_X1    g0954(.A1(new_n1151), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1154), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1148), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1148), .A2(new_n1157), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n882), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1160), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n882), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(new_n1163), .A3(new_n1158), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1161), .A2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1143), .B1(new_n1147), .B2(new_n1165), .ZN(new_n1166));
  XOR2_X1   g0966(.A(new_n1102), .B(KEYINPUT120), .Z(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(new_n1104), .ZN(new_n1168));
  AND2_X1   g0968(.A1(new_n1161), .A2(new_n1164), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1168), .A2(new_n1169), .A3(KEYINPUT57), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1166), .A2(new_n687), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1169), .A2(new_n798), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1157), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n783), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n826), .A2(new_n342), .ZN(new_n1175));
  INV_X1    g0975(.A(G41), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n254), .A2(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT116), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1178), .B(new_n342), .C1(G41), .C2(new_n252), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n734), .A2(G97), .B1(new_n775), .B2(new_n355), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1180), .B(KEYINPUT117), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1181), .B(new_n969), .C1(new_n741), .C2(new_n758), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n740), .A2(new_n221), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1176), .B(new_n258), .C1(new_n764), .C2(new_n244), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n744), .A2(new_n444), .B1(new_n761), .B2(new_n339), .ZN(new_n1185));
  NOR4_X1   g0985(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .A4(new_n1185), .ZN(new_n1186));
  XOR2_X1   g0986(.A(KEYINPUT118), .B(KEYINPUT58), .Z(new_n1187));
  XNOR2_X1  g0987(.A(new_n1186), .B(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1126), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1189), .A2(new_n761), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n807), .A2(G125), .B1(new_n748), .B2(G150), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT119), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1190), .B(new_n1192), .C1(G137), .C2(new_n775), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n1128), .B2(new_n733), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G128), .B2(new_n765), .ZN(new_n1195));
  XOR2_X1   g0995(.A(new_n1195), .B(KEYINPUT59), .Z(new_n1196));
  AOI21_X1  g0996(.A(new_n1178), .B1(G124), .B2(new_n759), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n265), .B2(new_n740), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1179), .B(new_n1188), .C1(new_n1196), .C2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(new_n730), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1174), .A2(new_n799), .A3(new_n1175), .A4(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1172), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1171), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT121), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1204), .B(new_n1205), .ZN(G375));
  NAND2_X1  g1006(.A1(new_n826), .A2(new_n208), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n252), .B1(new_n747), .B2(new_n342), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1183), .B(new_n1208), .C1(G128), .C2(new_n759), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1209), .B1(new_n414), .B2(new_n755), .C1(new_n265), .C2(new_n761), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT122), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n770), .A2(G137), .B1(G132), .B2(new_n807), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1211), .B(new_n1212), .C1(new_n733), .C2(new_n1189), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n258), .B1(new_n755), .B2(new_n244), .C1(new_n213), .C2(new_n761), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n744), .A2(new_n474), .B1(new_n740), .B2(new_n339), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n758), .A2(new_n518), .ZN(new_n1216));
  NOR4_X1   g1016(.A1(new_n1214), .A2(new_n1012), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n444), .B2(new_n733), .C1(new_n741), .C2(new_n764), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1020), .B1(new_n1213), .B2(new_n1218), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n803), .B(new_n1219), .C1(new_n878), .C2(new_n783), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n1092), .A2(new_n798), .B1(new_n1207), .B2(new_n1220), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1070), .B(new_n1102), .C1(new_n1079), .C2(new_n1091), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1221), .B1(new_n1223), .B2(new_n933), .ZN(G381));
  INV_X1    g1024(.A(KEYINPUT123), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1106), .B(new_n688), .C1(new_n1146), .C2(new_n1100), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1112), .B1(new_n1111), .B2(new_n1102), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1092), .A2(KEYINPUT114), .A3(new_n1103), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1100), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(KEYINPUT113), .B1(new_n1104), .B2(new_n687), .ZN(new_n1230));
  NOR3_X1   g1030(.A1(new_n1226), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1225), .B1(new_n1231), .B2(new_n1140), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1117), .A2(new_n1141), .A3(KEYINPUT123), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(G375), .A2(new_n1235), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n964), .A2(new_n1055), .A3(new_n987), .A4(new_n1059), .ZN(new_n1237));
  NOR3_X1   g1037(.A1(new_n1237), .A2(G381), .A3(G384), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(G393), .A2(G396), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1236), .A2(new_n1238), .A3(new_n1239), .ZN(G407));
  NAND2_X1  g1040(.A1(new_n657), .A2(G213), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1241), .B(KEYINPUT124), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1236), .A2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(G407), .A2(G213), .A3(new_n1243), .ZN(G409));
  XOR2_X1   g1044(.A(G393), .B(G396), .Z(new_n1245));
  AND4_X1   g1045(.A1(new_n964), .A2(new_n1055), .A3(new_n987), .A4(new_n1059), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n964), .A2(new_n987), .B1(new_n1055), .B2(new_n1059), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1245), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(G387), .A2(G390), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1245), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1249), .A2(new_n1250), .A3(new_n1237), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1248), .A2(new_n1251), .ZN(new_n1252));
  OR2_X1    g1052(.A1(G384), .A2(KEYINPUT126), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1146), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT125), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(new_n1111), .B2(new_n1102), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT60), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1254), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1222), .A2(KEYINPUT125), .A3(new_n1257), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n687), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1221), .B(new_n1253), .C1(new_n1258), .C2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(G384), .A2(KEYINPUT126), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1261), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1222), .ZN(new_n1265));
  OAI21_X1  g1065(.A(KEYINPUT60), .B1(new_n1265), .B2(new_n1255), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1266), .A2(new_n687), .A3(new_n1254), .A4(new_n1259), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1267), .A2(new_n1221), .A3(new_n1253), .A4(new_n1262), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1264), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1147), .A2(new_n1165), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n932), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1203), .A2(new_n1272), .ZN(new_n1273));
  AND3_X1   g1073(.A1(new_n1117), .A2(KEYINPUT123), .A3(new_n1141), .ZN(new_n1274));
  AOI21_X1  g1074(.A(KEYINPUT123), .B1(new_n1117), .B2(new_n1141), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1273), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(G378), .A2(new_n1171), .A3(new_n1203), .ZN(new_n1277));
  AOI211_X1 g1077(.A(new_n1242), .B(new_n1270), .C1(new_n1276), .C2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1252), .B1(KEYINPUT63), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1242), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1202), .B1(new_n932), .B2(new_n1271), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1281), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1277), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1280), .B(new_n1269), .C1(new_n1282), .C2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1242), .A2(G2897), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1264), .A2(new_n1268), .A3(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1285), .B1(new_n1264), .B2(new_n1268), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1288), .B1(new_n1289), .B2(new_n1280), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT63), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1284), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT61), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1279), .A2(new_n1292), .A3(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1284), .A2(KEYINPUT62), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1280), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1288), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1295), .A2(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1293), .B1(new_n1284), .B2(KEYINPUT62), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1252), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1294), .A2(new_n1301), .ZN(G405));
  NOR2_X1   g1102(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1303));
  AOI21_X1  g1103(.A(KEYINPUT121), .B1(new_n1171), .B2(new_n1203), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1234), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1270), .B1(new_n1305), .B2(new_n1277), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1252), .A2(KEYINPUT127), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1305), .A2(new_n1277), .A3(new_n1270), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT127), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1248), .A2(new_n1310), .A3(new_n1251), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1307), .A2(new_n1308), .A3(new_n1309), .A4(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1309), .ZN(new_n1313));
  OAI211_X1 g1113(.A(KEYINPUT127), .B(new_n1252), .C1(new_n1313), .C2(new_n1306), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1312), .A2(new_n1314), .ZN(G402));
endmodule


