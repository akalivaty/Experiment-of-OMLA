//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 1 0 1 1 1 1 1 0 1 1 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n757, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n831, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958;
  INV_X1    g000(.A(G22gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G228gat), .A2(G233gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT22), .ZN(new_n204));
  INV_X1    g003(.A(G211gat), .ZN(new_n205));
  INV_X1    g004(.A(G218gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT71), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT71), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n209), .B(new_n204), .C1(new_n205), .C2(new_n206), .ZN(new_n210));
  XNOR2_X1  g009(.A(G197gat), .B(G204gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n208), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  XOR2_X1   g011(.A(G211gat), .B(G218gat), .Z(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n213), .ZN(new_n215));
  NAND4_X1  g014(.A1(new_n215), .A2(new_n208), .A3(new_n210), .A4(new_n211), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AND2_X1   g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G148gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT76), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT76), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(G148gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n222), .A2(new_n224), .A3(G141gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n221), .A2(G141gat), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n220), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G155gat), .A2(G162gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT2), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT77), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT77), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n229), .A2(new_n232), .A3(KEYINPUT2), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT2), .ZN(new_n235));
  INV_X1    g034(.A(G141gat), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n236), .A2(G148gat), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n235), .B1(new_n226), .B2(new_n237), .ZN(new_n238));
  AOI22_X1  g037(.A1(new_n228), .A2(new_n234), .B1(new_n220), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT29), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n217), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT83), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n225), .A2(new_n227), .ZN(new_n246));
  INV_X1    g045(.A(new_n220), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n246), .A2(new_n234), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n238), .A2(new_n220), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT29), .B1(new_n214), .B2(new_n216), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n250), .B1(new_n251), .B2(KEYINPUT3), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n252), .B1(new_n243), .B2(new_n244), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n203), .B1(new_n245), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT84), .ZN(new_n255));
  AND2_X1   g054(.A1(new_n251), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n240), .B1(new_n251), .B2(new_n255), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n250), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT85), .ZN(new_n259));
  AOI221_X4 g058(.A(KEYINPUT3), .B1(new_n238), .B2(new_n220), .C1(new_n228), .C2(new_n234), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n259), .B1(new_n260), .B2(KEYINPUT29), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n241), .A2(KEYINPUT85), .A3(new_n242), .ZN(new_n262));
  INV_X1    g061(.A(new_n217), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n258), .A2(G228gat), .A3(G233gat), .A4(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n202), .B1(new_n254), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n254), .A2(new_n265), .A3(new_n202), .ZN(new_n268));
  XNOR2_X1  g067(.A(G78gat), .B(G106gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(KEYINPUT31), .B(G50gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n267), .A2(new_n268), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n271), .ZN(new_n273));
  INV_X1    g072(.A(new_n268), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n273), .B1(new_n274), .B2(new_n266), .ZN(new_n275));
  AND2_X1   g074(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G57gat), .B(G85gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(KEYINPUT80), .ZN(new_n278));
  XOR2_X1   g077(.A(KEYINPUT79), .B(KEYINPUT0), .Z(new_n279));
  OR2_X1    g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n279), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G1gat), .B(G29gat), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n280), .A2(new_n283), .A3(new_n281), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G225gat), .A2(G233gat), .ZN(new_n288));
  INV_X1    g087(.A(G120gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(G113gat), .ZN(new_n290));
  INV_X1    g089(.A(G113gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(G120gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT1), .ZN(new_n294));
  XNOR2_X1  g093(.A(G127gat), .B(G134gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT68), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n293), .B(new_n294), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G134gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(G127gat), .ZN(new_n299));
  INV_X1    g098(.A(G127gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(G134gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n296), .A2(new_n294), .ZN(new_n303));
  XNOR2_X1  g102(.A(G113gat), .B(G120gat), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n302), .B(new_n303), .C1(new_n304), .C2(KEYINPUT1), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n297), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n306), .B1(new_n239), .B2(new_n240), .ZN(new_n307));
  OAI21_X1  g106(.A(KEYINPUT78), .B1(new_n307), .B2(new_n260), .ZN(new_n308));
  AND2_X1   g107(.A1(new_n297), .A2(new_n305), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n309), .B1(new_n250), .B2(KEYINPUT3), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT78), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n310), .A2(new_n311), .A3(new_n241), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT4), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n314), .B1(new_n250), .B2(new_n306), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n239), .A2(new_n309), .A3(KEYINPUT4), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n288), .B1(new_n313), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT39), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n287), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n250), .A2(new_n306), .ZN(new_n321));
  AOI22_X1  g120(.A1(new_n248), .A2(new_n249), .B1(new_n297), .B2(new_n305), .ZN(new_n322));
  OR2_X1    g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n288), .ZN(new_n324));
  OAI21_X1  g123(.A(KEYINPUT39), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n320), .B1(new_n318), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT40), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n324), .B1(new_n321), .B2(new_n322), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT5), .ZN(new_n330));
  AND3_X1   g129(.A1(new_n315), .A2(new_n288), .A3(new_n316), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n330), .B1(new_n313), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT5), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n315), .A2(new_n333), .A3(new_n288), .A4(new_n316), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n334), .B1(new_n308), .B2(new_n312), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n287), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n320), .B(KEYINPUT40), .C1(new_n318), .C2(new_n325), .ZN(new_n337));
  AND3_X1   g136(.A1(new_n328), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(G183gat), .ZN(new_n339));
  INV_X1    g138(.A(G190gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OR2_X1    g142(.A1(KEYINPUT66), .A2(KEYINPUT24), .ZN(new_n344));
  NAND2_X1  g143(.A1(G183gat), .A2(G190gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(KEYINPUT66), .A2(KEYINPUT24), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(G169gat), .A2(G176gat), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT64), .B(KEYINPUT23), .ZN(new_n351));
  INV_X1    g150(.A(G169gat), .ZN(new_n352));
  INV_X1    g151(.A(G176gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n350), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n352), .A2(new_n353), .A3(KEYINPUT65), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT65), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n357), .B1(G169gat), .B2(G176gat), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n356), .A2(new_n358), .A3(KEYINPUT23), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n348), .A2(new_n355), .A3(KEYINPUT25), .A4(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT24), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n362), .A2(new_n341), .A3(new_n342), .ZN(new_n363));
  AND2_X1   g162(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n364));
  NOR2_X1   g163(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n354), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n352), .A2(new_n353), .A3(KEYINPUT23), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n363), .A2(new_n366), .A3(new_n349), .A4(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT25), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n360), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n339), .A2(KEYINPUT27), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT27), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(G183gat), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n372), .A2(new_n374), .A3(new_n340), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT28), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT27), .B(G183gat), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n378), .A2(KEYINPUT28), .A3(new_n340), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT26), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n356), .A2(new_n358), .A3(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n383), .A2(new_n349), .ZN(new_n384));
  AOI22_X1  g183(.A1(new_n382), .A2(new_n384), .B1(G183gat), .B2(G190gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n242), .ZN(new_n388));
  NAND2_X1  g187(.A1(G226gat), .A2(G233gat), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n263), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT67), .ZN(new_n391));
  AND3_X1   g190(.A1(new_n380), .A2(new_n385), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n391), .B1(new_n380), .B2(new_n385), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n371), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT72), .ZN(new_n395));
  INV_X1    g194(.A(new_n389), .ZN(new_n396));
  AND3_X1   g195(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n395), .B1(new_n394), .B2(new_n396), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n390), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  XOR2_X1   g198(.A(G8gat), .B(G36gat), .Z(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(KEYINPUT73), .ZN(new_n401));
  XNOR2_X1  g200(.A(G64gat), .B(G92gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n396), .A2(KEYINPUT29), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n360), .A2(new_n370), .B1(new_n380), .B2(new_n385), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n394), .A2(new_n404), .B1(new_n405), .B2(new_n396), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n263), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n399), .A2(new_n403), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT75), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT30), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n399), .A2(KEYINPUT75), .A3(new_n407), .A4(new_n403), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n399), .A2(new_n403), .A3(new_n407), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n407), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n403), .B(KEYINPUT74), .ZN(new_n416));
  AOI22_X1  g215(.A1(new_n414), .A2(KEYINPUT30), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n276), .B1(new_n338), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT82), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT6), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n420), .B1(new_n336), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n311), .B1(new_n310), .B2(new_n241), .ZN(new_n423));
  NOR3_X1   g222(.A1(new_n307), .A2(KEYINPUT78), .A3(new_n260), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n331), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n330), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n334), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n287), .B1(new_n313), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT6), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n336), .ZN(new_n431));
  INV_X1    g230(.A(new_n335), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n427), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n433), .A2(KEYINPUT82), .A3(KEYINPUT6), .A4(new_n287), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n422), .A2(new_n431), .A3(new_n434), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n415), .A2(KEYINPUT37), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n217), .B1(new_n388), .B2(new_n389), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n437), .B1(new_n397), .B2(new_n398), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT37), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n439), .B1(new_n406), .B2(new_n217), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT38), .ZN(new_n442));
  AND2_X1   g241(.A1(new_n416), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n410), .B(new_n412), .C1(new_n436), .C2(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n435), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n403), .B1(new_n415), .B2(KEYINPUT37), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n436), .B1(new_n447), .B2(KEYINPUT87), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT87), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n439), .B1(new_n399), .B2(new_n407), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n449), .B1(new_n450), .B2(new_n403), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n442), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n446), .B1(new_n452), .B2(KEYINPUT88), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT88), .ZN(new_n454));
  AOI211_X1 g253(.A(new_n454), .B(new_n442), .C1(new_n448), .C2(new_n451), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n419), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT86), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n272), .A2(new_n275), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT81), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n430), .A2(new_n459), .A3(new_n336), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n459), .B1(new_n430), .B2(new_n336), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n434), .B(new_n422), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  AND2_X1   g261(.A1(new_n413), .A2(new_n417), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n458), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(G71gat), .B(G99gat), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT69), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n465), .B(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(G15gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n465), .B(KEYINPUT69), .ZN(new_n469));
  INV_X1    g268(.A(G15gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AND3_X1   g270(.A1(new_n468), .A2(new_n471), .A3(G43gat), .ZN(new_n472));
  AOI21_X1  g271(.A(G43gat), .B1(new_n468), .B2(new_n471), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n394), .A2(new_n306), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n371), .B(new_n309), .C1(new_n392), .C2(new_n393), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(G227gat), .A2(G233gat), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT33), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n475), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n479), .B1(new_n476), .B2(new_n477), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT32), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  AOI221_X4 g287(.A(new_n485), .B1(new_n474), .B2(KEYINPUT33), .C1(new_n478), .C2(new_n480), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  XOR2_X1   g289(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n491));
  OAI21_X1  g290(.A(new_n491), .B1(new_n478), .B2(new_n480), .ZN(new_n492));
  INV_X1    g291(.A(new_n491), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n476), .A2(new_n479), .A3(new_n477), .A4(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n488), .A2(new_n490), .A3(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n474), .B1(new_n484), .B2(KEYINPUT33), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n498), .A2(new_n486), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n495), .B1(new_n499), .B2(new_n489), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n497), .A2(new_n500), .A3(KEYINPUT36), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT36), .B1(new_n497), .B2(new_n500), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n457), .B1(new_n464), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT36), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n496), .B1(new_n488), .B2(new_n490), .ZN(new_n506));
  NOR3_X1   g305(.A1(new_n499), .A2(new_n489), .A3(new_n495), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n497), .A2(new_n500), .A3(KEYINPUT36), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n431), .A2(KEYINPUT81), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n430), .A2(new_n336), .A3(new_n459), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n422), .A2(new_n434), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n418), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n510), .B(KEYINPUT86), .C1(new_n515), .C2(new_n458), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n456), .A2(new_n504), .A3(new_n516), .ZN(new_n517));
  NOR2_X1   g316(.A1(KEYINPUT89), .A2(KEYINPUT35), .ZN(new_n518));
  AND2_X1   g317(.A1(KEYINPUT89), .A2(KEYINPUT35), .ZN(new_n519));
  NOR3_X1   g318(.A1(new_n418), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n506), .A2(new_n507), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n520), .A2(new_n435), .A3(new_n458), .A4(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n462), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n458), .ZN(new_n524));
  NOR3_X1   g323(.A1(new_n523), .A2(new_n524), .A3(new_n418), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT35), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n522), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n517), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT90), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT90), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n517), .A2(new_n530), .A3(new_n527), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(G229gat), .A2(G233gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(G15gat), .B(G22gat), .ZN(new_n534));
  INV_X1    g333(.A(G1gat), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n534), .A2(KEYINPUT16), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT94), .ZN(new_n537));
  INV_X1    g336(.A(G8gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n536), .B(new_n539), .C1(new_n535), .C2(new_n534), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n537), .A2(new_n538), .ZN(new_n541));
  OR2_X1    g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n540), .A2(new_n541), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NOR3_X1   g344(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT91), .ZN(new_n547));
  OAI21_X1  g346(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n549), .B1(new_n547), .B2(new_n548), .ZN(new_n550));
  NAND2_X1  g349(.A1(G29gat), .A2(G36gat), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AND2_X1   g351(.A1(G43gat), .A2(G50gat), .ZN(new_n553));
  NOR2_X1   g352(.A1(G43gat), .A2(G50gat), .ZN(new_n554));
  OAI21_X1  g353(.A(KEYINPUT15), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT92), .B(G43gat), .ZN(new_n556));
  INV_X1    g355(.A(G50gat), .ZN(new_n557));
  AOI211_X1 g356(.A(KEYINPUT15), .B(new_n553), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n548), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n555), .B(new_n551), .C1(new_n559), .C2(new_n546), .ZN(new_n560));
  OAI22_X1  g359(.A1(new_n552), .A2(new_n555), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT93), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n561), .A2(new_n563), .A3(KEYINPUT17), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT17), .B1(new_n561), .B2(new_n563), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n544), .B(KEYINPUT95), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n533), .B(new_n562), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(KEYINPUT96), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n533), .B(KEYINPUT13), .Z(new_n571));
  INV_X1    g370(.A(KEYINPUT97), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n572), .B1(new_n545), .B2(new_n561), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(new_n562), .ZN(new_n574));
  AOI22_X1  g373(.A1(new_n570), .A2(KEYINPUT18), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT18), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n569), .A2(KEYINPUT96), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G113gat), .B(G141gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(G197gat), .ZN(new_n580));
  XOR2_X1   g379(.A(KEYINPUT11), .B(G169gat), .Z(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n582), .B(KEYINPUT12), .Z(new_n583));
  NAND2_X1  g382(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n583), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n575), .A2(new_n577), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G134gat), .B(G162gat), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT103), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G85gat), .A2(G92gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT7), .ZN(new_n594));
  NAND2_X1  g393(.A1(G99gat), .A2(G106gat), .ZN(new_n595));
  INV_X1    g394(.A(G85gat), .ZN(new_n596));
  INV_X1    g395(.A(G92gat), .ZN(new_n597));
  AOI22_X1  g396(.A1(KEYINPUT8), .A2(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G99gat), .B(G106gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT100), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n604), .B1(new_n565), .B2(new_n566), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n561), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT101), .ZN(new_n607));
  NAND3_X1  g406(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n608));
  AND3_X1   g407(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n607), .B1(new_n606), .B2(new_n608), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n605), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT102), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT102), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n613), .B(new_n605), .C1(new_n609), .C2(new_n610), .ZN(new_n614));
  XNOR2_X1  g413(.A(G190gat), .B(G218gat), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n612), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n616), .B1(new_n612), .B2(new_n614), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n592), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n612), .A2(new_n614), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(new_n615), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n612), .A2(new_n614), .A3(new_n616), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n590), .B(new_n591), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  OR2_X1    g424(.A1(G57gat), .A2(G64gat), .ZN(new_n626));
  NAND2_X1  g425(.A1(G57gat), .A2(G64gat), .ZN(new_n627));
  AND2_X1   g426(.A1(G71gat), .A2(G78gat), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n626), .B(new_n627), .C1(new_n628), .C2(KEYINPUT9), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT98), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(G71gat), .A2(G78gat), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n631), .B(new_n633), .Z(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(new_n601), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT10), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n631), .B(new_n633), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n603), .A2(KEYINPUT10), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(G230gat), .ZN(new_n641));
  INV_X1    g440(.A(G233gat), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  OR2_X1    g444(.A1(new_n635), .A2(new_n644), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(G120gat), .B(G148gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(G176gat), .B(G204gat), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n648), .B(new_n649), .Z(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n645), .A2(new_n646), .A3(new_n650), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n638), .A2(KEYINPUT21), .ZN(new_n655));
  XNOR2_X1  g454(.A(G127gat), .B(G155gat), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n655), .B(new_n656), .Z(new_n657));
  AOI21_X1  g456(.A(new_n545), .B1(KEYINPUT21), .B2(new_n638), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(G231gat), .A2(G233gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT99), .ZN(new_n661));
  XOR2_X1   g460(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(G183gat), .B(G211gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n659), .B(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n625), .A2(new_n654), .A3(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n532), .A2(new_n587), .A3(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n669), .A2(new_n462), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(new_n535), .ZN(G1324gat));
  AND2_X1   g470(.A1(new_n532), .A2(new_n587), .ZN(new_n672));
  XOR2_X1   g471(.A(KEYINPUT16), .B(G8gat), .Z(new_n673));
  NAND4_X1  g472(.A1(new_n672), .A2(new_n418), .A3(new_n668), .A4(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(G8gat), .B1(new_n669), .B2(new_n463), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  MUX2_X1   g475(.A(new_n674), .B(new_n676), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g476(.A(G15gat), .B1(new_n669), .B2(new_n510), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n521), .A2(new_n470), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n678), .B1(new_n669), .B2(new_n679), .ZN(G1326gat));
  NOR2_X1   g479(.A1(new_n669), .A2(new_n458), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT43), .B(G22gat), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n681), .B(new_n682), .Z(G1327gat));
  AND2_X1   g482(.A1(new_n619), .A2(new_n624), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n529), .A2(new_n531), .A3(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n464), .A2(new_n503), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n456), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n527), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(new_n625), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n685), .ZN(new_n692));
  INV_X1    g491(.A(new_n587), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n666), .A2(new_n654), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n687), .A2(new_n692), .A3(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT106), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n687), .A2(KEYINPUT106), .A3(new_n692), .A4(new_n696), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n699), .A2(new_n523), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(KEYINPUT107), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT107), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n699), .A2(new_n703), .A3(new_n523), .A4(new_n700), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n702), .A2(G29gat), .A3(new_n704), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n532), .A2(new_n587), .A3(new_n625), .A4(new_n694), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n462), .A2(G29gat), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT105), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n708), .B(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n705), .A2(new_n712), .ZN(G1328gat));
  INV_X1    g512(.A(G36gat), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n418), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(KEYINPUT46), .B1(new_n706), .B2(new_n715), .ZN(new_n716));
  OR3_X1    g515(.A1(new_n706), .A2(KEYINPUT46), .A3(new_n715), .ZN(new_n717));
  AND3_X1   g516(.A1(new_n699), .A2(new_n418), .A3(new_n700), .ZN(new_n718));
  OAI211_X1 g517(.A(new_n716), .B(new_n717), .C1(new_n718), .C2(new_n714), .ZN(G1329gat));
  INV_X1    g518(.A(new_n556), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n720), .B1(new_n697), .B2(new_n510), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n521), .A2(new_n556), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n721), .B(KEYINPUT47), .C1(new_n706), .C2(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n706), .A2(new_n722), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n699), .A2(new_n503), .A3(new_n700), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n724), .B1(new_n725), .B2(new_n720), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n723), .B1(new_n726), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g526(.A(G50gat), .B1(new_n697), .B2(new_n458), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n276), .A2(new_n557), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n728), .B(KEYINPUT48), .C1(new_n706), .C2(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n706), .A2(new_n729), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n699), .A2(new_n276), .A3(new_n700), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n731), .B1(new_n732), .B2(G50gat), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n730), .B1(new_n733), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g533(.A(new_n654), .ZN(new_n735));
  NOR4_X1   g534(.A1(new_n625), .A2(new_n587), .A3(new_n735), .A4(new_n667), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT108), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n737), .A2(new_n690), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n523), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g539(.A(new_n463), .B(KEYINPUT109), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n742), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n738), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT110), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT110), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n738), .A2(new_n746), .A3(new_n743), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  OR2_X1    g547(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1333gat));
  INV_X1    g549(.A(G71gat), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n738), .A2(new_n751), .A3(new_n521), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n738), .A2(new_n503), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n753), .B2(new_n751), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(G1334gat));
  NAND2_X1  g555(.A1(new_n738), .A2(new_n276), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(G78gat), .ZN(G1335gat));
  AND2_X1   g557(.A1(new_n687), .A2(new_n692), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n587), .A2(new_n735), .A3(new_n666), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(G85gat), .B1(new_n761), .B2(new_n462), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n587), .A2(new_n666), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n690), .A2(KEYINPUT51), .A3(new_n625), .A4(new_n763), .ZN(new_n764));
  OR2_X1    g563(.A1(new_n764), .A2(KEYINPUT111), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(KEYINPUT111), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n690), .A2(new_n625), .A3(new_n763), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT51), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n765), .A2(new_n766), .A3(new_n769), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n770), .A2(new_n596), .A3(new_n523), .A4(new_n654), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n762), .A2(new_n771), .ZN(G1336gat));
  OAI21_X1  g571(.A(G92gat), .B1(new_n761), .B2(new_n742), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n742), .A2(G92gat), .A3(new_n735), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT52), .B1(new_n770), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n759), .A2(new_n418), .A3(new_n760), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n769), .A2(new_n764), .ZN(new_n778));
  AOI22_X1  g577(.A1(new_n777), .A2(G92gat), .B1(new_n778), .B2(new_n774), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n776), .B1(new_n779), .B2(new_n780), .ZN(G1337gat));
  XOR2_X1   g580(.A(KEYINPUT112), .B(G99gat), .Z(new_n782));
  NAND4_X1  g581(.A1(new_n770), .A2(new_n521), .A3(new_n654), .A4(new_n782), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n761), .A2(new_n510), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n783), .B1(new_n784), .B2(new_n782), .ZN(G1338gat));
  NAND3_X1  g584(.A1(new_n759), .A2(new_n276), .A3(new_n760), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(G106gat), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT53), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n735), .A2(new_n458), .A3(G106gat), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n770), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n787), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n786), .A2(G106gat), .B1(new_n778), .B2(new_n789), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n791), .B1(new_n788), .B2(new_n792), .ZN(G1339gat));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n637), .A2(new_n639), .A3(new_n643), .ZN(new_n795));
  AND3_X1   g594(.A1(new_n645), .A2(KEYINPUT54), .A3(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n640), .A2(new_n797), .A3(new_n644), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n651), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n794), .B1(new_n796), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n645), .A2(KEYINPUT54), .A3(new_n795), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n801), .A2(KEYINPUT55), .A3(new_n651), .A4(new_n798), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n802), .A2(new_n653), .ZN(new_n803));
  INV_X1    g602(.A(new_n586), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n585), .B1(new_n575), .B2(new_n577), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n800), .B(new_n803), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  OR2_X1    g605(.A1(new_n567), .A2(new_n568), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n533), .B1(new_n807), .B2(new_n562), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n574), .A2(new_n571), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n582), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n586), .A2(new_n654), .A3(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n684), .A2(new_n806), .A3(new_n811), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n803), .A2(new_n586), .A3(new_n810), .A4(new_n800), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n666), .B1(new_n625), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n684), .A2(new_n693), .A3(new_n735), .A4(new_n666), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n523), .A2(new_n521), .ZN(new_n819));
  NOR4_X1   g618(.A1(new_n818), .A2(new_n276), .A3(new_n741), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n587), .A2(new_n291), .ZN(new_n821));
  XOR2_X1   g620(.A(new_n821), .B(KEYINPUT114), .Z(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n820), .A2(new_n587), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(G113gat), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n825), .A2(KEYINPUT113), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n825), .A2(KEYINPUT113), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n823), .B1(new_n826), .B2(new_n827), .ZN(G1340gat));
  NAND2_X1  g627(.A1(new_n820), .A2(new_n654), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g629(.A1(new_n820), .A2(new_n666), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n831), .B(G127gat), .ZN(G1342gat));
  NOR2_X1   g631(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n818), .A2(new_n276), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n625), .A2(new_n463), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n835), .A2(G134gat), .A3(new_n819), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n833), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n820), .A2(new_n625), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(G134gat), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n841), .A2(KEYINPUT115), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n841), .A2(KEYINPUT115), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n839), .B1(new_n842), .B2(new_n843), .ZN(G1343gat));
  NAND2_X1  g643(.A1(new_n510), .A2(new_n523), .ZN(new_n845));
  OR2_X1    g644(.A1(new_n741), .A2(new_n845), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n815), .A2(KEYINPUT117), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n816), .B1(new_n815), .B2(KEYINPUT117), .ZN(new_n848));
  OAI211_X1 g647(.A(KEYINPUT57), .B(new_n276), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n817), .A2(new_n276), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT57), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n846), .B1(new_n849), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n853), .A2(G141gat), .A3(new_n587), .ZN(new_n854));
  NAND2_X1  g653(.A1(KEYINPUT118), .A2(KEYINPUT58), .ZN(new_n855));
  NOR2_X1   g654(.A1(KEYINPUT118), .A2(KEYINPUT58), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n850), .A2(new_n846), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n587), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n856), .B1(new_n858), .B2(new_n236), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n854), .A2(new_n855), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n855), .B1(new_n854), .B2(new_n859), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n860), .A2(new_n861), .ZN(G1344gat));
  AND2_X1   g661(.A1(new_n222), .A2(new_n224), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n857), .A2(new_n863), .A3(new_n654), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT59), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n846), .A2(KEYINPUT119), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n846), .A2(KEYINPUT119), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n654), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n817), .A2(KEYINPUT57), .A3(new_n276), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n868), .B1(new_n852), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT120), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n221), .B1(new_n870), .B2(new_n871), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n865), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AOI211_X1 g673(.A(KEYINPUT59), .B(new_n863), .C1(new_n853), .C2(new_n654), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n864), .B1(new_n874), .B2(new_n875), .ZN(G1345gat));
  INV_X1    g675(.A(G155gat), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n857), .A2(new_n877), .A3(new_n666), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n853), .A2(new_n666), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n878), .B1(new_n879), .B2(new_n877), .ZN(G1346gat));
  NOR4_X1   g679(.A1(new_n850), .A2(G162gat), .A3(new_n835), .A4(new_n845), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  AOI211_X1 g681(.A(new_n684), .B(new_n846), .C1(new_n849), .C2(new_n852), .ZN(new_n883));
  INV_X1    g682(.A(G162gat), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT121), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI211_X1 g686(.A(KEYINPUT121), .B(new_n882), .C1(new_n883), .C2(new_n884), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(G1347gat));
  NOR2_X1   g688(.A1(new_n523), .A2(new_n463), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(new_n524), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n817), .A2(new_n892), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n893), .A2(new_n352), .A3(new_n693), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT122), .B1(new_n818), .B2(new_n523), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT122), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n817), .A2(new_n896), .A3(new_n462), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n742), .A2(new_n524), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n898), .A2(new_n587), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n894), .B1(new_n900), .B2(new_n352), .ZN(G1348gat));
  OAI21_X1  g700(.A(G176gat), .B1(new_n893), .B2(new_n735), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n898), .A2(new_n899), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n654), .A2(new_n353), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n902), .B1(new_n903), .B2(new_n904), .ZN(G1349gat));
  OAI21_X1  g704(.A(G183gat), .B1(new_n893), .B2(new_n667), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n666), .A2(new_n378), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n906), .B1(new_n903), .B2(new_n907), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g708(.A(new_n893), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n340), .B1(new_n910), .B2(new_n625), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT123), .ZN(new_n912));
  OR3_X1    g711(.A1(new_n911), .A2(new_n912), .A3(KEYINPUT61), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n625), .A2(new_n340), .ZN(new_n914));
  OAI21_X1  g713(.A(KEYINPUT61), .B1(new_n911), .B2(new_n912), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n911), .A2(new_n912), .ZN(new_n916));
  OAI221_X1 g715(.A(new_n913), .B1(new_n903), .B2(new_n914), .C1(new_n915), .C2(new_n916), .ZN(G1351gat));
  NAND3_X1  g716(.A1(new_n741), .A2(new_n276), .A3(new_n510), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n918), .B1(new_n895), .B2(new_n897), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT124), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n693), .A2(G197gat), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n891), .A2(new_n503), .ZN(new_n923));
  AOI21_X1  g722(.A(KEYINPUT57), .B1(new_n817), .B2(new_n276), .ZN(new_n924));
  AOI211_X1 g723(.A(new_n851), .B(new_n458), .C1(new_n815), .C2(new_n816), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n587), .B(new_n923), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(KEYINPUT124), .B1(new_n926), .B2(G197gat), .ZN(new_n927));
  INV_X1    g726(.A(new_n921), .ZN(new_n928));
  AOI211_X1 g727(.A(new_n918), .B(new_n928), .C1(new_n895), .C2(new_n897), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n922), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(KEYINPUT125), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT125), .ZN(new_n932));
  OAI211_X1 g731(.A(new_n922), .B(new_n932), .C1(new_n927), .C2(new_n929), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(G1352gat));
  INV_X1    g733(.A(G204gat), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n919), .A2(new_n935), .A3(new_n654), .ZN(new_n936));
  OR2_X1    g735(.A1(new_n936), .A2(KEYINPUT62), .ZN(new_n937));
  INV_X1    g736(.A(new_n923), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n938), .B1(new_n852), .B2(new_n869), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(new_n654), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(G204gat), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n936), .A2(KEYINPUT62), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n937), .A2(new_n941), .A3(new_n942), .ZN(G1353gat));
  NAND3_X1  g742(.A1(new_n919), .A2(new_n205), .A3(new_n666), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT126), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n939), .A2(new_n666), .ZN(new_n946));
  AND4_X1   g745(.A1(new_n945), .A2(new_n946), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT63), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n205), .B1(KEYINPUT126), .B2(new_n948), .ZN(new_n949));
  AOI22_X1  g748(.A1(new_n946), .A2(new_n949), .B1(new_n945), .B2(KEYINPUT63), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n944), .B1(new_n947), .B2(new_n950), .ZN(G1354gat));
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n919), .A2(new_n206), .A3(new_n625), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n206), .B1(new_n939), .B2(new_n625), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n952), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n939), .A2(new_n625), .ZN(new_n957));
  OAI211_X1 g756(.A(KEYINPUT127), .B(new_n953), .C1(new_n957), .C2(new_n206), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n956), .A2(new_n958), .ZN(G1355gat));
endmodule


