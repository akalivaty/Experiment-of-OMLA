

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589;

  OR2_X1 U323 ( .A1(n403), .A2(n574), .ZN(n379) );
  XNOR2_X1 U324 ( .A(n306), .B(n305), .ZN(n312) );
  XNOR2_X1 U325 ( .A(n304), .B(n294), .ZN(n305) );
  NOR2_X1 U326 ( .A1(n550), .A2(n549), .ZN(n291) );
  AND2_X1 U327 ( .A1(G230GAT), .A2(G233GAT), .ZN(n292) );
  XOR2_X1 U328 ( .A(n361), .B(n360), .Z(n293) );
  AND2_X1 U329 ( .A1(G228GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U330 ( .A(KEYINPUT47), .B(KEYINPUT106), .ZN(n454) );
  XNOR2_X1 U331 ( .A(n428), .B(n292), .ZN(n430) );
  XNOR2_X1 U332 ( .A(n455), .B(n454), .ZN(n462) );
  XNOR2_X1 U333 ( .A(n430), .B(n429), .ZN(n433) );
  XNOR2_X1 U334 ( .A(KEYINPUT48), .B(KEYINPUT108), .ZN(n463) );
  XNOR2_X1 U335 ( .A(n464), .B(n463), .ZN(n547) );
  XNOR2_X1 U336 ( .A(n296), .B(G204GAT), .ZN(n297) );
  XNOR2_X1 U337 ( .A(n298), .B(n297), .ZN(n442) );
  XNOR2_X1 U338 ( .A(n362), .B(n293), .ZN(n367) );
  XNOR2_X1 U339 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U340 ( .A(n367), .B(n366), .ZN(n372) );
  XNOR2_X1 U341 ( .A(n444), .B(n443), .ZN(n458) );
  NOR2_X1 U342 ( .A1(n514), .A2(n445), .ZN(n446) );
  XNOR2_X1 U343 ( .A(n374), .B(n373), .ZN(n553) );
  INV_X1 U344 ( .A(KEYINPUT98), .ZN(n494) );
  XNOR2_X1 U345 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U346 ( .A(n447), .B(G50GAT), .ZN(n448) );
  XNOR2_X1 U347 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U348 ( .A(n473), .B(n472), .ZN(G1343GAT) );
  XNOR2_X1 U349 ( .A(n449), .B(n448), .ZN(G1331GAT) );
  XNOR2_X1 U350 ( .A(G148GAT), .B(KEYINPUT67), .ZN(n295) );
  XNOR2_X1 U351 ( .A(n295), .B(KEYINPUT68), .ZN(n298) );
  XNOR2_X1 U352 ( .A(G78GAT), .B(G106GAT), .ZN(n296) );
  XOR2_X1 U353 ( .A(KEYINPUT82), .B(G218GAT), .Z(n300) );
  XOR2_X1 U354 ( .A(G141GAT), .B(G22GAT), .Z(n411) );
  XNOR2_X1 U355 ( .A(G50GAT), .B(G162GAT), .ZN(n313) );
  XOR2_X1 U356 ( .A(n411), .B(n313), .Z(n299) );
  XNOR2_X1 U357 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U358 ( .A(n442), .B(n301), .ZN(n306) );
  XOR2_X1 U359 ( .A(KEYINPUT23), .B(KEYINPUT81), .Z(n303) );
  XNOR2_X1 U360 ( .A(KEYINPUT22), .B(KEYINPUT24), .ZN(n302) );
  XNOR2_X1 U361 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U362 ( .A(G155GAT), .B(KEYINPUT84), .Z(n308) );
  XNOR2_X1 U363 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n307) );
  XNOR2_X1 U364 ( .A(n308), .B(n307), .ZN(n386) );
  XOR2_X1 U365 ( .A(G211GAT), .B(KEYINPUT83), .Z(n310) );
  XNOR2_X1 U366 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n309) );
  XNOR2_X1 U367 ( .A(n310), .B(n309), .ZN(n355) );
  XNOR2_X1 U368 ( .A(n386), .B(n355), .ZN(n311) );
  XNOR2_X1 U369 ( .A(n312), .B(n311), .ZN(n550) );
  XOR2_X1 U370 ( .A(n550), .B(KEYINPUT28), .Z(n520) );
  XNOR2_X1 U371 ( .A(G106GAT), .B(KEYINPUT10), .ZN(n314) );
  XNOR2_X1 U372 ( .A(n314), .B(n313), .ZN(n328) );
  XNOR2_X1 U373 ( .A(G99GAT), .B(G85GAT), .ZN(n315) );
  XNOR2_X1 U374 ( .A(n315), .B(KEYINPUT69), .ZN(n436) );
  XOR2_X1 U375 ( .A(G92GAT), .B(n436), .Z(n317) );
  NAND2_X1 U376 ( .A1(G232GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U377 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U378 ( .A(KEYINPUT71), .B(KEYINPUT11), .Z(n319) );
  XNOR2_X1 U379 ( .A(G134GAT), .B(KEYINPUT9), .ZN(n318) );
  XNOR2_X1 U380 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U381 ( .A(n321), .B(n320), .Z(n326) );
  XOR2_X1 U382 ( .A(G29GAT), .B(G43GAT), .Z(n323) );
  XNOR2_X1 U383 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n322) );
  XNOR2_X1 U384 ( .A(n323), .B(n322), .ZN(n412) );
  XNOR2_X1 U385 ( .A(G36GAT), .B(G190GAT), .ZN(n324) );
  XNOR2_X1 U386 ( .A(n324), .B(G218GAT), .ZN(n354) );
  XNOR2_X1 U387 ( .A(n412), .B(n354), .ZN(n325) );
  XNOR2_X1 U388 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U389 ( .A(n328), .B(n327), .ZN(n563) );
  XNOR2_X1 U390 ( .A(KEYINPUT36), .B(n563), .ZN(n585) );
  XOR2_X1 U391 ( .A(G57GAT), .B(KEYINPUT13), .Z(n440) );
  XOR2_X1 U392 ( .A(n440), .B(G71GAT), .Z(n330) );
  XOR2_X1 U393 ( .A(G15GAT), .B(G1GAT), .Z(n413) );
  XNOR2_X1 U394 ( .A(n413), .B(G183GAT), .ZN(n329) );
  XNOR2_X1 U395 ( .A(n330), .B(n329), .ZN(n334) );
  XOR2_X1 U396 ( .A(KEYINPUT73), .B(KEYINPUT15), .Z(n332) );
  XNOR2_X1 U397 ( .A(G8GAT), .B(KEYINPUT14), .ZN(n331) );
  XNOR2_X1 U398 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U399 ( .A(n334), .B(n333), .Z(n336) );
  XNOR2_X1 U400 ( .A(G22GAT), .B(G127GAT), .ZN(n335) );
  XNOR2_X1 U401 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U402 ( .A(KEYINPUT74), .B(G64GAT), .Z(n338) );
  NAND2_X1 U403 ( .A1(G231GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U404 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U405 ( .A(n340), .B(n339), .Z(n345) );
  XOR2_X1 U406 ( .A(KEYINPUT12), .B(G211GAT), .Z(n342) );
  XNOR2_X1 U407 ( .A(G78GAT), .B(G155GAT), .ZN(n341) );
  XNOR2_X1 U408 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U409 ( .A(n343), .B(KEYINPUT72), .ZN(n344) );
  XOR2_X1 U410 ( .A(n345), .B(n344), .Z(n476) );
  INV_X1 U411 ( .A(n476), .ZN(n582) );
  XNOR2_X1 U412 ( .A(KEYINPUT79), .B(KEYINPUT19), .ZN(n346) );
  XNOR2_X1 U413 ( .A(n346), .B(G183GAT), .ZN(n347) );
  XOR2_X1 U414 ( .A(n347), .B(KEYINPUT78), .Z(n349) );
  XNOR2_X1 U415 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n348) );
  XNOR2_X1 U416 ( .A(n349), .B(n348), .ZN(n374) );
  XOR2_X1 U417 ( .A(G169GAT), .B(G8GAT), .Z(n424) );
  XOR2_X1 U418 ( .A(G204GAT), .B(n424), .Z(n351) );
  NAND2_X1 U419 ( .A1(G226GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U420 ( .A(n351), .B(n350), .ZN(n353) );
  XNOR2_X1 U421 ( .A(G176GAT), .B(G92GAT), .ZN(n352) );
  XNOR2_X1 U422 ( .A(n352), .B(G64GAT), .ZN(n429) );
  XOR2_X1 U423 ( .A(n353), .B(n429), .Z(n357) );
  XNOR2_X1 U424 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U425 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U426 ( .A(n374), .B(n358), .ZN(n546) );
  XOR2_X1 U427 ( .A(KEYINPUT27), .B(KEYINPUT90), .Z(n359) );
  XOR2_X1 U428 ( .A(n546), .B(n359), .Z(n403) );
  XOR2_X1 U429 ( .A(G120GAT), .B(G71GAT), .Z(n428) );
  XNOR2_X1 U430 ( .A(G169GAT), .B(n428), .ZN(n362) );
  XOR2_X1 U431 ( .A(KEYINPUT77), .B(G176GAT), .Z(n361) );
  NAND2_X1 U432 ( .A1(G227GAT), .A2(G233GAT), .ZN(n360) );
  XOR2_X1 U433 ( .A(KEYINPUT20), .B(G99GAT), .Z(n364) );
  XNOR2_X1 U434 ( .A(G43GAT), .B(G15GAT), .ZN(n363) );
  XNOR2_X1 U435 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U436 ( .A(n365), .B(G190GAT), .Z(n366) );
  XOR2_X1 U437 ( .A(KEYINPUT76), .B(G134GAT), .Z(n369) );
  XNOR2_X1 U438 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n368) );
  XNOR2_X1 U439 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U440 ( .A(G113GAT), .B(n370), .Z(n390) );
  XNOR2_X1 U441 ( .A(n390), .B(KEYINPUT80), .ZN(n371) );
  XNOR2_X1 U442 ( .A(n372), .B(n371), .ZN(n373) );
  NAND2_X1 U443 ( .A1(n553), .A2(n550), .ZN(n375) );
  XNOR2_X1 U444 ( .A(KEYINPUT26), .B(n375), .ZN(n574) );
  NOR2_X1 U445 ( .A1(n553), .A2(n546), .ZN(n376) );
  NOR2_X1 U446 ( .A1(n550), .A2(n376), .ZN(n377) );
  XNOR2_X1 U447 ( .A(n377), .B(KEYINPUT25), .ZN(n378) );
  NAND2_X1 U448 ( .A1(n379), .A2(n378), .ZN(n401) );
  XOR2_X1 U449 ( .A(KEYINPUT87), .B(KEYINPUT88), .Z(n381) );
  XNOR2_X1 U450 ( .A(KEYINPUT85), .B(KEYINPUT4), .ZN(n380) );
  XNOR2_X1 U451 ( .A(n381), .B(n380), .ZN(n385) );
  XOR2_X1 U452 ( .A(KEYINPUT86), .B(KEYINPUT1), .Z(n383) );
  XNOR2_X1 U453 ( .A(G1GAT), .B(G57GAT), .ZN(n382) );
  XNOR2_X1 U454 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U455 ( .A(n385), .B(n384), .Z(n392) );
  XOR2_X1 U456 ( .A(n386), .B(KEYINPUT6), .Z(n388) );
  NAND2_X1 U457 ( .A1(G225GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U458 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U459 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U460 ( .A(n392), .B(n391), .ZN(n400) );
  XOR2_X1 U461 ( .A(KEYINPUT89), .B(KEYINPUT5), .Z(n394) );
  XNOR2_X1 U462 ( .A(G141GAT), .B(G148GAT), .ZN(n393) );
  XNOR2_X1 U463 ( .A(n394), .B(n393), .ZN(n398) );
  XOR2_X1 U464 ( .A(G85GAT), .B(G162GAT), .Z(n396) );
  XNOR2_X1 U465 ( .A(G29GAT), .B(G120GAT), .ZN(n395) );
  XNOR2_X1 U466 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U467 ( .A(n398), .B(n397), .Z(n399) );
  XNOR2_X1 U468 ( .A(n400), .B(n399), .ZN(n571) );
  NAND2_X1 U469 ( .A1(n401), .A2(n571), .ZN(n402) );
  XNOR2_X1 U470 ( .A(n402), .B(KEYINPUT91), .ZN(n407) );
  INV_X1 U471 ( .A(n520), .ZN(n405) );
  NOR2_X1 U472 ( .A1(n571), .A2(n403), .ZN(n465) );
  NAND2_X1 U473 ( .A1(n465), .A2(n553), .ZN(n404) );
  NOR2_X1 U474 ( .A1(n405), .A2(n404), .ZN(n406) );
  NOR2_X1 U475 ( .A1(n407), .A2(n406), .ZN(n408) );
  XNOR2_X1 U476 ( .A(KEYINPUT92), .B(n408), .ZN(n479) );
  NOR2_X1 U477 ( .A1(n582), .A2(n479), .ZN(n409) );
  NAND2_X1 U478 ( .A1(n585), .A2(n409), .ZN(n410) );
  XOR2_X1 U479 ( .A(KEYINPUT37), .B(n410), .Z(n514) );
  XNOR2_X1 U480 ( .A(n412), .B(n411), .ZN(n414) );
  XNOR2_X1 U481 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U482 ( .A(KEYINPUT64), .B(KEYINPUT30), .Z(n416) );
  NAND2_X1 U483 ( .A1(G229GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U484 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U485 ( .A(n418), .B(n417), .Z(n423) );
  XOR2_X1 U486 ( .A(KEYINPUT65), .B(KEYINPUT66), .Z(n420) );
  XNOR2_X1 U487 ( .A(G113GAT), .B(G197GAT), .ZN(n419) );
  XNOR2_X1 U488 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U489 ( .A(n421), .B(KEYINPUT29), .ZN(n422) );
  XNOR2_X1 U490 ( .A(n423), .B(n422), .ZN(n425) );
  XOR2_X1 U491 ( .A(n425), .B(n424), .Z(n427) );
  XNOR2_X1 U492 ( .A(G50GAT), .B(G36GAT), .ZN(n426) );
  XOR2_X1 U493 ( .A(n427), .B(n426), .Z(n501) );
  INV_X1 U494 ( .A(n433), .ZN(n431) );
  NAND2_X1 U495 ( .A1(n431), .A2(KEYINPUT32), .ZN(n435) );
  INV_X1 U496 ( .A(KEYINPUT32), .ZN(n432) );
  NAND2_X1 U497 ( .A1(n433), .A2(n432), .ZN(n434) );
  NAND2_X1 U498 ( .A1(n435), .A2(n434), .ZN(n438) );
  XNOR2_X1 U499 ( .A(n436), .B(KEYINPUT31), .ZN(n437) );
  XNOR2_X1 U500 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U501 ( .A(n439), .B(KEYINPUT33), .Z(n444) );
  XNOR2_X1 U502 ( .A(n440), .B(KEYINPUT70), .ZN(n441) );
  INV_X1 U503 ( .A(n458), .ZN(n578) );
  NOR2_X1 U504 ( .A1(n501), .A2(n578), .ZN(n481) );
  INV_X1 U505 ( .A(n481), .ZN(n445) );
  XOR2_X1 U506 ( .A(KEYINPUT38), .B(n446), .Z(n497) );
  NOR2_X1 U507 ( .A1(n520), .A2(n497), .ZN(n449) );
  INV_X1 U508 ( .A(KEYINPUT100), .ZN(n447) );
  INV_X1 U509 ( .A(n501), .ZN(n575) );
  XNOR2_X1 U510 ( .A(n458), .B(KEYINPUT41), .ZN(n556) );
  NAND2_X1 U511 ( .A1(n575), .A2(n556), .ZN(n451) );
  XOR2_X1 U512 ( .A(KEYINPUT105), .B(KEYINPUT46), .Z(n450) );
  XNOR2_X1 U513 ( .A(n451), .B(n450), .ZN(n453) );
  NOR2_X1 U514 ( .A1(n563), .A2(n582), .ZN(n452) );
  NAND2_X1 U515 ( .A1(n453), .A2(n452), .ZN(n455) );
  NAND2_X1 U516 ( .A1(n582), .A2(n585), .ZN(n457) );
  XNOR2_X1 U517 ( .A(KEYINPUT45), .B(KEYINPUT107), .ZN(n456) );
  XNOR2_X1 U518 ( .A(n457), .B(n456), .ZN(n459) );
  NAND2_X1 U519 ( .A1(n459), .A2(n458), .ZN(n460) );
  NOR2_X1 U520 ( .A1(n460), .A2(n575), .ZN(n461) );
  NOR2_X1 U521 ( .A1(n462), .A2(n461), .ZN(n464) );
  INV_X1 U522 ( .A(n547), .ZN(n466) );
  NAND2_X1 U523 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U524 ( .A(n467), .B(KEYINPUT109), .ZN(n532) );
  NAND2_X1 U525 ( .A1(n532), .A2(n520), .ZN(n468) );
  NOR2_X1 U526 ( .A1(n553), .A2(n468), .ZN(n469) );
  XNOR2_X1 U527 ( .A(KEYINPUT110), .B(n469), .ZN(n529) );
  AND2_X1 U528 ( .A1(n529), .A2(n563), .ZN(n473) );
  XNOR2_X1 U529 ( .A(KEYINPUT51), .B(KEYINPUT113), .ZN(n471) );
  INV_X1 U530 ( .A(G134GAT), .ZN(n470) );
  XOR2_X1 U531 ( .A(KEYINPUT93), .B(KEYINPUT34), .Z(n475) );
  XNOR2_X1 U532 ( .A(G1GAT), .B(KEYINPUT94), .ZN(n474) );
  XNOR2_X1 U533 ( .A(n475), .B(n474), .ZN(n483) );
  NOR2_X1 U534 ( .A1(n563), .A2(n476), .ZN(n478) );
  XNOR2_X1 U535 ( .A(KEYINPUT16), .B(KEYINPUT75), .ZN(n477) );
  XNOR2_X1 U536 ( .A(n478), .B(n477), .ZN(n480) );
  NOR2_X1 U537 ( .A1(n480), .A2(n479), .ZN(n502) );
  NAND2_X1 U538 ( .A1(n481), .A2(n502), .ZN(n489) );
  NOR2_X1 U539 ( .A1(n571), .A2(n489), .ZN(n482) );
  XOR2_X1 U540 ( .A(n483), .B(n482), .Z(G1324GAT) );
  NOR2_X1 U541 ( .A1(n546), .A2(n489), .ZN(n485) );
  XNOR2_X1 U542 ( .A(G8GAT), .B(KEYINPUT95), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n485), .B(n484), .ZN(G1325GAT) );
  NOR2_X1 U544 ( .A1(n553), .A2(n489), .ZN(n487) );
  XNOR2_X1 U545 ( .A(KEYINPUT35), .B(KEYINPUT96), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U547 ( .A(G15GAT), .B(n488), .ZN(G1326GAT) );
  NOR2_X1 U548 ( .A1(n520), .A2(n489), .ZN(n490) );
  XOR2_X1 U549 ( .A(G22GAT), .B(n490), .Z(G1327GAT) );
  NOR2_X1 U550 ( .A1(n497), .A2(n571), .ZN(n492) );
  XNOR2_X1 U551 ( .A(KEYINPUT97), .B(KEYINPUT39), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n492), .B(n491), .ZN(n493) );
  XOR2_X1 U553 ( .A(G29GAT), .B(n493), .Z(G1328GAT) );
  NOR2_X1 U554 ( .A1(n497), .A2(n546), .ZN(n495) );
  XNOR2_X1 U555 ( .A(G36GAT), .B(n496), .ZN(G1329GAT) );
  NOR2_X1 U556 ( .A1(n497), .A2(n553), .ZN(n499) );
  XNOR2_X1 U557 ( .A(KEYINPUT99), .B(KEYINPUT40), .ZN(n498) );
  XNOR2_X1 U558 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U559 ( .A(G43GAT), .B(n500), .ZN(G1330GAT) );
  NAND2_X1 U560 ( .A1(n501), .A2(n556), .ZN(n513) );
  INV_X1 U561 ( .A(n513), .ZN(n503) );
  NAND2_X1 U562 ( .A1(n503), .A2(n502), .ZN(n509) );
  NOR2_X1 U563 ( .A1(n571), .A2(n509), .ZN(n505) );
  XNOR2_X1 U564 ( .A(KEYINPUT101), .B(KEYINPUT42), .ZN(n504) );
  XNOR2_X1 U565 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(n506), .ZN(G1332GAT) );
  NOR2_X1 U567 ( .A1(n546), .A2(n509), .ZN(n507) );
  XOR2_X1 U568 ( .A(G64GAT), .B(n507), .Z(G1333GAT) );
  NOR2_X1 U569 ( .A1(n553), .A2(n509), .ZN(n508) );
  XOR2_X1 U570 ( .A(G71GAT), .B(n508), .Z(G1334GAT) );
  NOR2_X1 U571 ( .A1(n520), .A2(n509), .ZN(n511) );
  XNOR2_X1 U572 ( .A(KEYINPUT102), .B(KEYINPUT43), .ZN(n510) );
  XNOR2_X1 U573 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U574 ( .A(G78GAT), .B(n512), .ZN(G1335GAT) );
  OR2_X1 U575 ( .A1(n514), .A2(n513), .ZN(n519) );
  NOR2_X1 U576 ( .A1(n571), .A2(n519), .ZN(n515) );
  XOR2_X1 U577 ( .A(G85GAT), .B(n515), .Z(G1336GAT) );
  NOR2_X1 U578 ( .A1(n546), .A2(n519), .ZN(n516) );
  XOR2_X1 U579 ( .A(G92GAT), .B(n516), .Z(G1337GAT) );
  NOR2_X1 U580 ( .A1(n553), .A2(n519), .ZN(n518) );
  XNOR2_X1 U581 ( .A(G99GAT), .B(KEYINPUT103), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n518), .B(n517), .ZN(G1338GAT) );
  NOR2_X1 U583 ( .A1(n520), .A2(n519), .ZN(n522) );
  XNOR2_X1 U584 ( .A(KEYINPUT44), .B(KEYINPUT104), .ZN(n521) );
  XNOR2_X1 U585 ( .A(n522), .B(n521), .ZN(n523) );
  XOR2_X1 U586 ( .A(G106GAT), .B(n523), .Z(G1339GAT) );
  NAND2_X1 U587 ( .A1(n529), .A2(n575), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n524), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT49), .B(KEYINPUT112), .Z(n526) );
  NAND2_X1 U590 ( .A1(n529), .A2(n556), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n526), .B(n525), .ZN(n528) );
  XOR2_X1 U592 ( .A(G120GAT), .B(KEYINPUT111), .Z(n527) );
  XNOR2_X1 U593 ( .A(n528), .B(n527), .ZN(G1341GAT) );
  NAND2_X1 U594 ( .A1(n529), .A2(n582), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n530), .B(KEYINPUT50), .ZN(n531) );
  XNOR2_X1 U596 ( .A(G127GAT), .B(n531), .ZN(G1342GAT) );
  INV_X1 U597 ( .A(n574), .ZN(n533) );
  NAND2_X1 U598 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U599 ( .A(KEYINPUT114), .B(n534), .Z(n543) );
  NAND2_X1 U600 ( .A1(n575), .A2(n543), .ZN(n535) );
  XNOR2_X1 U601 ( .A(G141GAT), .B(n535), .ZN(G1344GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT53), .B(KEYINPUT116), .Z(n537) );
  XNOR2_X1 U603 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U605 ( .A(KEYINPUT115), .B(n538), .Z(n540) );
  NAND2_X1 U606 ( .A1(n543), .A2(n556), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(G1345GAT) );
  XOR2_X1 U608 ( .A(G155GAT), .B(KEYINPUT117), .Z(n542) );
  NAND2_X1 U609 ( .A1(n582), .A2(n543), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n542), .B(n541), .ZN(G1346GAT) );
  NAND2_X1 U611 ( .A1(n543), .A2(n563), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n544), .B(KEYINPUT118), .ZN(n545) );
  XNOR2_X1 U613 ( .A(G162GAT), .B(n545), .ZN(G1347GAT) );
  NOR2_X1 U614 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n548), .B(KEYINPUT54), .ZN(n572) );
  INV_X1 U616 ( .A(n571), .ZN(n549) );
  AND2_X1 U617 ( .A1(n572), .A2(n291), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n551), .B(KEYINPUT55), .ZN(n552) );
  NOR2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n564) );
  NAND2_X1 U620 ( .A1(n564), .A2(n575), .ZN(n554) );
  XOR2_X1 U621 ( .A(KEYINPUT119), .B(n554), .Z(n555) );
  XNOR2_X1 U622 ( .A(G169GAT), .B(n555), .ZN(G1348GAT) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n560) );
  XOR2_X1 U624 ( .A(KEYINPUT120), .B(KEYINPUT56), .Z(n558) );
  NAND2_X1 U625 ( .A1(n564), .A2(n556), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1349GAT) );
  XOR2_X1 U628 ( .A(G183GAT), .B(KEYINPUT121), .Z(n562) );
  NAND2_X1 U629 ( .A1(n564), .A2(n582), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n562), .B(n561), .ZN(G1350GAT) );
  XNOR2_X1 U631 ( .A(G190GAT), .B(KEYINPUT122), .ZN(n568) );
  XOR2_X1 U632 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n566) );
  NAND2_X1 U633 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U634 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(G1351GAT) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n569), .B(KEYINPUT60), .ZN(n570) );
  XOR2_X1 U638 ( .A(KEYINPUT124), .B(n570), .Z(n577) );
  NAND2_X1 U639 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n586) );
  NAND2_X1 U641 ( .A1(n586), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n580) );
  NAND2_X1 U644 ( .A1(n586), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XOR2_X1 U646 ( .A(G204GAT), .B(n581), .Z(G1353GAT) );
  NAND2_X1 U647 ( .A1(n586), .A2(n582), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n583), .B(KEYINPUT126), .ZN(n584) );
  XNOR2_X1 U649 ( .A(G211GAT), .B(n584), .ZN(G1354GAT) );
  XOR2_X1 U650 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n588) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

