//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0 0 0 1 0 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 1 1 0 1 0 0 1 1 1 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1281, new_n1282, new_n1283, new_n1284, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1360, new_n1361;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  XOR2_X1   g0010(.A(KEYINPUT66), .B(G244), .Z(new_n211));
  AND2_X1   g0011(.A1(new_n211), .A2(G77), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G87), .A2(G250), .ZN(new_n216));
  NAND4_X1  g0016(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n210), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT67), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n210), .A2(G13), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n221), .B(G250), .C1(G257), .C2(G264), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT0), .ZN(new_n223));
  AND3_X1   g0023(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n224));
  AOI21_X1  g0024(.A(KEYINPUT64), .B1(G1), .B2(G13), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  AND2_X1   g0027(.A1(KEYINPUT65), .A2(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(KEYINPUT65), .A2(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(G50), .B1(G58), .B2(G68), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n223), .B(new_n234), .C1(new_n218), .C2(KEYINPUT1), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n220), .A2(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT2), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G226), .ZN(new_n239));
  INV_X1    g0039(.A(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT68), .B(KEYINPUT69), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G68), .B(G77), .Z(new_n251));
  XOR2_X1   g0051(.A(G50), .B(G58), .Z(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(new_n250), .B(new_n253), .Z(G351));
  INV_X1    g0054(.A(KEYINPUT13), .ZN(new_n255));
  AND2_X1   g0055(.A1(G33), .A2(G41), .ZN(new_n256));
  NOR3_X1   g0056(.A1(new_n224), .A2(new_n225), .A3(new_n256), .ZN(new_n257));
  AND2_X1   g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1698), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT70), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT70), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G1698), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n262), .A2(new_n264), .A3(G226), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G232), .A2(G1698), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n260), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G97), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n257), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT76), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI211_X1 g0072(.A(KEYINPUT76), .B(new_n257), .C1(new_n267), .C2(new_n269), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G1), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n275), .B1(G41), .B2(G45), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  INV_X1    g0078(.A(G41), .ZN(new_n279));
  OAI211_X1 g0079(.A(G1), .B(G13), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n277), .A2(new_n280), .A3(G274), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n276), .ZN(new_n282));
  INV_X1    g0082(.A(G238), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n255), .B1(new_n274), .B2(new_n285), .ZN(new_n286));
  AOI211_X1 g0086(.A(KEYINPUT13), .B(new_n284), .C1(new_n272), .C2(new_n273), .ZN(new_n287));
  OAI21_X1  g0087(.A(G200), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT70), .B(G1698), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n289), .A2(G226), .B1(G232), .B2(G1698), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n268), .B1(new_n290), .B2(new_n260), .ZN(new_n291));
  AOI21_X1  g0091(.A(KEYINPUT76), .B1(new_n291), .B2(new_n257), .ZN(new_n292));
  INV_X1    g0092(.A(new_n273), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n285), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT13), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n274), .A2(new_n255), .A3(new_n285), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n295), .A2(G190), .A3(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(G20), .A2(G33), .ZN(new_n298));
  AOI22_X1  g0098(.A1(new_n298), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n230), .A2(G33), .ZN(new_n300));
  INV_X1    g0100(.A(G77), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n303), .B1(new_n224), .B2(new_n225), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n305), .B(KEYINPUT11), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n275), .A2(G13), .A3(G20), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n308), .A2(KEYINPUT77), .A3(new_n203), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT12), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT77), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n311), .B1(new_n307), .B2(G68), .ZN(new_n312));
  OR2_X1    g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n310), .A2(new_n312), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n307), .B(new_n303), .C1(new_n224), .C2(new_n225), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n203), .B1(new_n275), .B2(G20), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n313), .A2(new_n314), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n306), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n288), .A2(new_n297), .A3(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n286), .A2(new_n287), .ZN(new_n323));
  INV_X1    g0123(.A(G169), .ZN(new_n324));
  OAI21_X1  g0124(.A(KEYINPUT14), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n295), .A2(G179), .A3(new_n296), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT14), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n327), .B(G169), .C1(new_n286), .C2(new_n287), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n325), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n322), .B1(new_n329), .B2(new_n319), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n316), .A2(KEYINPUT72), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n275), .A2(G20), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT72), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n315), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(KEYINPUT71), .A2(G58), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT8), .ZN(new_n336));
  XNOR2_X1  g0136(.A(new_n335), .B(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n331), .A2(new_n332), .A3(new_n334), .A4(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n337), .A2(new_n308), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n289), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n343));
  INV_X1    g0143(.A(G87), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n343), .A2(new_n260), .B1(new_n278), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n257), .ZN(new_n346));
  INV_X1    g0146(.A(G190), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n281), .B1(new_n282), .B2(new_n240), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n346), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n348), .B1(new_n345), .B2(new_n257), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n350), .B1(G200), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n304), .ZN(new_n353));
  AND2_X1   g0153(.A1(G58), .A2(G68), .ZN(new_n354));
  NOR2_X1   g0154(.A1(G58), .A2(G68), .ZN(new_n355));
  OAI21_X1  g0155(.A(G20), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n298), .A2(G159), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(KEYINPUT78), .B1(new_n258), .B2(new_n259), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT3), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n278), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT78), .ZN(new_n362));
  NAND2_X1  g0162(.A1(KEYINPUT3), .A2(G33), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT7), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n359), .A2(new_n364), .A3(new_n365), .A4(new_n230), .ZN(new_n366));
  INV_X1    g0166(.A(G20), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n361), .A2(new_n367), .A3(new_n363), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n203), .B1(new_n368), .B2(KEYINPUT7), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n358), .B1(new_n366), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n353), .B1(new_n370), .B2(KEYINPUT16), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT79), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT16), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n230), .A2(new_n260), .A3(KEYINPUT7), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n368), .A2(new_n365), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n203), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n373), .B1(new_n376), .B2(new_n358), .ZN(new_n377));
  AND3_X1   g0177(.A1(new_n371), .A2(new_n372), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n372), .B1(new_n371), .B2(new_n377), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n342), .B(new_n352), .C1(new_n378), .C2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT17), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n366), .A2(new_n369), .ZN(new_n382));
  INV_X1    g0182(.A(new_n358), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n382), .A2(KEYINPUT16), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n304), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n374), .A2(new_n375), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(G68), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT16), .B1(new_n387), .B2(new_n383), .ZN(new_n388));
  OAI21_X1  g0188(.A(KEYINPUT79), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n371), .A2(new_n372), .A3(new_n377), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n341), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT17), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n391), .A2(new_n392), .A3(new_n352), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n381), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n351), .A2(G179), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n324), .B2(new_n351), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NOR3_X1   g0197(.A1(new_n391), .A2(new_n397), .A3(KEYINPUT18), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT18), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n342), .B1(new_n378), .B2(new_n379), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n399), .B1(new_n400), .B2(new_n396), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n281), .ZN(new_n403));
  INV_X1    g0203(.A(new_n282), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n403), .B1(new_n404), .B2(new_n211), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n361), .A2(new_n363), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(new_n283), .B2(new_n261), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n262), .A2(new_n264), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n408), .A2(new_n240), .ZN(new_n409));
  OAI221_X1 g0209(.A(new_n257), .B1(G107), .B2(new_n406), .C1(new_n407), .C2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n411), .A2(G179), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n412), .B1(new_n324), .B2(new_n411), .ZN(new_n413));
  XOR2_X1   g0213(.A(KEYINPUT8), .B(G58), .Z(new_n414));
  XNOR2_X1  g0214(.A(new_n414), .B(KEYINPUT73), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n298), .ZN(new_n416));
  INV_X1    g0216(.A(new_n300), .ZN(new_n417));
  XNOR2_X1  g0217(.A(KEYINPUT15), .B(G87), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  OR2_X1    g0219(.A1(KEYINPUT65), .A2(G20), .ZN(new_n420));
  NAND2_X1  g0220(.A1(KEYINPUT65), .A2(G20), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n417), .A2(new_n419), .B1(G77), .B2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n353), .B1(new_n416), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n332), .A2(G77), .ZN(new_n425));
  OAI22_X1  g0225(.A1(new_n315), .A2(new_n425), .B1(G77), .B2(new_n307), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n413), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n411), .A2(G200), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n427), .B(new_n430), .C1(new_n347), .C2(new_n411), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  AND4_X1   g0232(.A1(new_n330), .A2(new_n394), .A3(new_n402), .A4(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(G223), .ZN(new_n434));
  INV_X1    g0234(.A(G222), .ZN(new_n435));
  OAI221_X1 g0235(.A(new_n406), .B1(new_n434), .B2(new_n261), .C1(new_n408), .C2(new_n435), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n436), .B(new_n257), .C1(G77), .C2(new_n406), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n403), .B1(new_n404), .B2(G226), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OR2_X1    g0239(.A1(new_n439), .A2(G169), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n298), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(new_n300), .B2(new_n337), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n442), .A2(new_n304), .B1(new_n201), .B2(new_n308), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n331), .A2(G50), .A3(new_n332), .A4(new_n334), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(G179), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n439), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n440), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n439), .A2(G190), .ZN(new_n450));
  INV_X1    g0250(.A(G200), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n450), .B1(new_n451), .B2(new_n439), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n445), .A2(KEYINPUT74), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT74), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n443), .A2(new_n444), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT9), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n452), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT75), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n459), .B1(new_n456), .B2(new_n457), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NOR3_X1   g0261(.A1(new_n456), .A2(new_n459), .A3(new_n457), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n458), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT10), .ZN(new_n464));
  INV_X1    g0264(.A(new_n462), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n460), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT10), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n466), .A2(new_n467), .A3(new_n458), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n449), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n433), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n262), .A2(new_n264), .A3(G238), .ZN(new_n471));
  NAND2_X1  g0271(.A1(G244), .A2(G1698), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n260), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G116), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n257), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G45), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n477), .A2(G1), .ZN(new_n478));
  INV_X1    g0278(.A(G274), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(G250), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n481), .B1(new_n477), .B2(G1), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n480), .A2(new_n280), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(G169), .B1(new_n476), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n483), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n289), .A2(G238), .B1(G244), .B2(G1698), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n474), .B1(new_n486), .B2(new_n260), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n485), .B1(new_n487), .B2(new_n257), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n484), .B1(new_n446), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n420), .A2(new_n421), .A3(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT83), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n420), .A2(KEYINPUT83), .A3(new_n421), .A4(new_n490), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n344), .A2(new_n206), .A3(new_n207), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n420), .A2(G33), .A3(G97), .A4(new_n421), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT19), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n406), .A2(new_n230), .A3(G68), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n304), .B1(new_n496), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n278), .A2(G1), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n315), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n419), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n419), .A2(new_n307), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n502), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n504), .A2(G87), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n502), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n476), .A2(new_n347), .A3(new_n483), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n488), .B2(G200), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n489), .A2(new_n508), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n279), .A2(KEYINPUT5), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n275), .B(G45), .C1(new_n279), .C2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT81), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G41), .ZN(new_n519));
  AOI21_X1  g0319(.A(KEYINPUT81), .B1(new_n478), .B2(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(G257), .B(new_n280), .C1(new_n517), .C2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(G1), .A2(G13), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n256), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n523), .A2(new_n479), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n478), .A2(KEYINPUT81), .A3(new_n519), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n515), .A2(new_n516), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n524), .A2(new_n525), .A3(new_n526), .A4(new_n514), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n521), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G33), .A2(G283), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n481), .B1(new_n361), .B2(new_n363), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n530), .B1(new_n531), .B2(G1698), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT4), .ZN(new_n533));
  OAI21_X1  g0333(.A(G244), .B1(new_n258), .B2(new_n259), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n533), .B1(new_n534), .B2(new_n408), .ZN(new_n535));
  INV_X1    g0335(.A(G244), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n536), .B1(new_n361), .B2(new_n363), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n537), .A2(KEYINPUT4), .A3(new_n289), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n532), .A2(new_n535), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n257), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n528), .A2(new_n540), .A3(G190), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT82), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n307), .A2(G97), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n543), .B1(new_n504), .B2(G97), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n207), .B1(new_n374), .B2(new_n375), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n298), .A2(G77), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT6), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(KEYINPUT80), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT80), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(KEYINPUT6), .ZN(new_n552));
  NAND2_X1  g0352(.A1(G97), .A2(G107), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n550), .A2(new_n552), .B1(new_n208), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n206), .A2(G107), .ZN(new_n555));
  AND3_X1   g0355(.A1(new_n555), .A2(new_n550), .A3(new_n552), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n422), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n547), .A2(new_n548), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n545), .B1(new_n558), .B2(new_n304), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT82), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n528), .A2(new_n540), .A3(new_n560), .A4(G190), .ZN(new_n561));
  INV_X1    g0361(.A(new_n257), .ZN(new_n562));
  AOI21_X1  g0362(.A(KEYINPUT4), .B1(new_n537), .B2(new_n289), .ZN(new_n563));
  OAI211_X1 g0363(.A(G250), .B(G1698), .C1(new_n258), .C2(new_n259), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n529), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n562), .B1(new_n566), .B2(new_n538), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n521), .A2(new_n527), .ZN(new_n568));
  OAI21_X1  g0368(.A(G200), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n542), .A2(new_n559), .A3(new_n561), .A4(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n324), .B1(new_n567), .B2(new_n568), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n551), .A2(KEYINPUT6), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n549), .A2(KEYINPUT80), .ZN(new_n573));
  NOR2_X1   g0373(.A1(G97), .A2(G107), .ZN(new_n574));
  AND2_X1   g0374(.A1(G97), .A2(G107), .ZN(new_n575));
  OAI22_X1  g0375(.A1(new_n572), .A2(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n555), .A2(new_n550), .A3(new_n552), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n230), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n548), .ZN(new_n579));
  NOR3_X1   g0379(.A1(new_n546), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n544), .B1(new_n580), .B2(new_n353), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n528), .A2(new_n540), .A3(new_n446), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n571), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n504), .A2(G107), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n275), .A2(new_n207), .A3(G13), .A4(G20), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT25), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT86), .ZN(new_n588));
  XNOR2_X1  g0388(.A(new_n587), .B(new_n588), .ZN(new_n589));
  OR3_X1    g0389(.A1(new_n585), .A2(KEYINPUT85), .A3(new_n586), .ZN(new_n590));
  OAI21_X1  g0390(.A(KEYINPUT85), .B1(new_n585), .B2(new_n586), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n584), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  XNOR2_X1  g0393(.A(KEYINPUT84), .B(KEYINPUT22), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n420), .B(new_n421), .C1(new_n258), .C2(new_n259), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n595), .B1(new_n596), .B2(new_n344), .ZN(new_n597));
  OR2_X1    g0397(.A1(KEYINPUT23), .A2(G107), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n598), .B1(new_n420), .B2(new_n421), .ZN(new_n599));
  OAI21_X1  g0399(.A(KEYINPUT23), .B1(new_n367), .B2(G107), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n600), .B1(G20), .B2(new_n474), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n230), .A2(new_n406), .A3(new_n594), .A4(G87), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n597), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT24), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n353), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n597), .A2(new_n602), .A3(KEYINPUT24), .A4(new_n603), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n593), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(G250), .B1(new_n258), .B2(new_n259), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n609), .A2(new_n408), .ZN(new_n610));
  AND2_X1   g0410(.A1(G257), .A2(G1698), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(new_n258), .B2(new_n259), .ZN(new_n612));
  NAND2_X1  g0412(.A1(G33), .A2(G294), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n257), .B1(new_n610), .B2(new_n614), .ZN(new_n615));
  OAI211_X1 g0415(.A(G264), .B(new_n280), .C1(new_n517), .C2(new_n520), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(new_n616), .A3(new_n527), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n451), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n615), .A2(new_n616), .A3(new_n527), .A4(new_n347), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n608), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n513), .A2(new_n570), .A3(new_n583), .A4(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT21), .ZN(new_n623));
  INV_X1    g0423(.A(G116), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n315), .A2(new_n624), .A3(new_n503), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n307), .A2(G116), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n278), .A2(G97), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n627), .A2(new_n529), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n628), .A2(new_n230), .B1(G20), .B2(new_n624), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n629), .A2(KEYINPUT20), .A3(new_n304), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT20), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n627), .A2(new_n529), .ZN(new_n632));
  OAI22_X1  g0432(.A1(new_n422), .A2(new_n632), .B1(new_n367), .B2(G116), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n631), .B1(new_n633), .B2(new_n353), .ZN(new_n634));
  AOI211_X1 g0434(.A(new_n625), .B(new_n626), .C1(new_n630), .C2(new_n634), .ZN(new_n635));
  OAI211_X1 g0435(.A(G270), .B(new_n280), .C1(new_n517), .C2(new_n520), .ZN(new_n636));
  INV_X1    g0436(.A(G303), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n260), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(G264), .A2(G1698), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n406), .A2(new_n639), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n262), .A2(new_n264), .A3(G257), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n257), .B(new_n638), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n636), .A2(new_n642), .A3(new_n527), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(G169), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n623), .B1(new_n635), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n626), .B1(new_n630), .B2(new_n634), .ZN(new_n646));
  INV_X1    g0446(.A(new_n625), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n636), .A2(new_n642), .A3(new_n527), .A4(G179), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n645), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n617), .A2(new_n324), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n653), .B1(G179), .B2(new_n617), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n654), .A2(new_n608), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n648), .A2(KEYINPUT21), .A3(G169), .A4(new_n643), .ZN(new_n656));
  INV_X1    g0456(.A(new_n643), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(G190), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n643), .A2(G200), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(new_n635), .A3(new_n659), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n652), .A2(new_n655), .A3(new_n656), .A4(new_n660), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n470), .A2(new_n622), .A3(new_n661), .ZN(G372));
  AND2_X1   g0462(.A1(new_n381), .A2(new_n393), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n328), .A2(new_n326), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n295), .A2(new_n296), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n327), .B1(new_n665), .B2(G169), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n319), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n321), .A2(new_n428), .A3(new_n413), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n663), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(KEYINPUT18), .B1(new_n391), .B2(new_n397), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n400), .A2(new_n399), .A3(new_n396), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n468), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n467), .B1(new_n466), .B2(new_n458), .ZN(new_n674));
  OAI22_X1  g0474(.A1(new_n669), .A2(new_n672), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n675), .A2(new_n448), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n488), .A2(new_n446), .ZN(new_n677));
  INV_X1    g0477(.A(new_n484), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n508), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n680), .A2(new_n500), .A3(new_n499), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n506), .B1(new_n681), .B2(new_n304), .ZN(new_n682));
  INV_X1    g0482(.A(new_n511), .ZN(new_n683));
  AOI21_X1  g0483(.A(G200), .B1(new_n476), .B2(new_n483), .ZN(new_n684));
  OAI211_X1 g0484(.A(new_n682), .B(new_n509), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n621), .A2(new_n679), .A3(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT87), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n686), .A2(new_n687), .A3(new_n583), .A4(new_n570), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n570), .A2(new_n583), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n621), .A2(new_n679), .A3(new_n685), .ZN(new_n690));
  OAI21_X1  g0490(.A(KEYINPUT87), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n652), .A2(new_n656), .A3(new_n655), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n688), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT26), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT88), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n528), .A2(new_n540), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n557), .A2(new_n548), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n304), .B1(new_n697), .B2(new_n546), .ZN(new_n698));
  AOI22_X1  g0498(.A1(new_n696), .A2(new_n324), .B1(new_n698), .B2(new_n544), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n695), .B1(new_n699), .B2(new_n582), .ZN(new_n700));
  AND4_X1   g0500(.A1(new_n695), .A2(new_n571), .A3(new_n581), .A4(new_n582), .ZN(new_n701));
  OAI211_X1 g0501(.A(new_n694), .B(new_n513), .C1(new_n700), .C2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n679), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n699), .A2(new_n679), .A3(new_n685), .A4(new_n582), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n703), .B1(new_n704), .B2(KEYINPUT26), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n693), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n676), .B1(new_n470), .B2(new_n708), .ZN(G369));
  NAND3_X1  g0509(.A1(new_n656), .A2(new_n645), .A3(new_n651), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n230), .A2(new_n275), .A3(G13), .ZN(new_n711));
  OR2_X1    g0511(.A1(new_n711), .A2(KEYINPUT27), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(KEYINPUT27), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(G213), .A3(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(G343), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n648), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n710), .B1(new_n660), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n718), .B1(new_n710), .B2(new_n717), .ZN(new_n719));
  XOR2_X1   g0519(.A(new_n719), .B(KEYINPUT89), .Z(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(G330), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n716), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n621), .B1(new_n608), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(new_n655), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n654), .A2(new_n608), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n723), .ZN(new_n727));
  AND2_X1   g0527(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n722), .A2(new_n728), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n710), .A2(new_n723), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n729), .A2(new_n727), .A3(new_n731), .ZN(G399));
  NOR2_X1   g0532(.A1(new_n495), .A2(G116), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n221), .A2(new_n279), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n733), .A2(new_n734), .A3(G1), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n735), .B1(new_n232), .B2(new_n734), .ZN(new_n736));
  XNOR2_X1  g0536(.A(new_n736), .B(KEYINPUT90), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT28), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n513), .A2(new_n694), .A3(new_n582), .A4(new_n699), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n710), .A2(new_n726), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n679), .B(new_n739), .C1(new_n622), .C2(new_n740), .ZN(new_n741));
  OR2_X1    g0541(.A1(new_n700), .A2(new_n701), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n694), .B1(new_n742), .B2(new_n513), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n723), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(KEYINPUT29), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT29), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n707), .A2(new_n746), .A3(new_n723), .ZN(new_n747));
  AND2_X1   g0547(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(G330), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT30), .ZN(new_n750));
  AND4_X1   g0550(.A1(new_n476), .A2(new_n615), .A3(new_n483), .A4(new_n616), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n650), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n750), .B1(new_n752), .B2(new_n696), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n657), .A2(G179), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n476), .A2(new_n483), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n754), .A2(new_n696), .A3(new_n755), .A4(new_n617), .ZN(new_n756));
  INV_X1    g0556(.A(new_n696), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n757), .A2(KEYINPUT30), .A3(new_n650), .A4(new_n751), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n753), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  AND3_X1   g0559(.A1(new_n759), .A2(KEYINPUT31), .A3(new_n716), .ZN(new_n760));
  AOI21_X1  g0560(.A(KEYINPUT31), .B1(new_n759), .B2(new_n716), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n660), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n710), .A2(new_n726), .A3(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n689), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n764), .A2(new_n765), .A3(new_n686), .A4(new_n723), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n749), .B1(new_n762), .B2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n748), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n738), .B1(new_n770), .B2(G1), .ZN(G364));
  AND2_X1   g0571(.A1(new_n230), .A2(G13), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G45), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n773), .A2(G1), .A3(new_n734), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n722), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n776), .B1(G330), .B2(new_n720), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n227), .B1(G20), .B2(new_n324), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n778), .A2(KEYINPUT94), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(KEYINPUT94), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n347), .A2(G200), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n230), .B1(new_n446), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n206), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n230), .A2(new_n446), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n451), .A2(G190), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n785), .B1(G68), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT95), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n422), .A2(new_n446), .A3(new_n787), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G107), .ZN(new_n794));
  NOR2_X1   g0594(.A1(G190), .A2(G200), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n786), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n786), .A2(new_n783), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n794), .B1(new_n796), .B2(new_n301), .C1(new_n202), .C2(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n422), .A2(new_n446), .A3(new_n795), .ZN(new_n799));
  INV_X1    g0599(.A(G159), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n799), .A2(KEYINPUT32), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n347), .A2(new_n451), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n802), .A2(G20), .A3(new_n446), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n260), .B1(new_n804), .B2(G87), .ZN(new_n805));
  OAI21_X1  g0605(.A(KEYINPUT32), .B1(new_n799), .B2(new_n800), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n786), .A2(new_n802), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n805), .B(new_n806), .C1(new_n201), .C2(new_n807), .ZN(new_n808));
  OR4_X1    g0608(.A1(new_n791), .A2(new_n798), .A3(new_n801), .A4(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(G326), .ZN(new_n810));
  XOR2_X1   g0610(.A(KEYINPUT33), .B(G317), .Z(new_n811));
  OAI22_X1  g0611(.A1(new_n810), .A2(new_n807), .B1(new_n788), .B2(new_n811), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n803), .B(KEYINPUT96), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n812), .B1(G303), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n784), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n406), .B1(new_n815), .B2(G294), .ZN(new_n816));
  INV_X1    g0616(.A(new_n796), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n817), .A2(G311), .B1(G283), .B2(new_n793), .ZN(new_n818));
  INV_X1    g0618(.A(new_n797), .ZN(new_n819));
  INV_X1    g0619(.A(new_n799), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n819), .A2(G322), .B1(G329), .B2(new_n820), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n814), .A2(new_n816), .A3(new_n818), .A4(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n782), .B1(new_n809), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(G13), .A2(G33), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n825), .A2(G20), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n781), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n253), .A2(G45), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT92), .Z(new_n829));
  NAND2_X1  g0629(.A1(new_n359), .A2(new_n364), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n221), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(KEYINPUT93), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n829), .B(new_n833), .C1(G45), .C2(new_n232), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n406), .A2(new_n221), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT91), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(G355), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n834), .B(new_n837), .C1(G116), .C2(new_n221), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n774), .B(new_n823), .C1(new_n827), .C2(new_n838), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT97), .ZN(new_n840));
  INV_X1    g0640(.A(new_n826), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n840), .B1(new_n720), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n777), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(G396));
  OAI21_X1  g0644(.A(new_n431), .B1(new_n427), .B2(new_n723), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n429), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n413), .A2(new_n428), .A3(new_n723), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n708), .B2(new_n716), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n432), .A2(new_n723), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(new_n693), .B2(new_n706), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n775), .B1(new_n853), .B2(new_n768), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n768), .B2(new_n853), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n781), .A2(new_n824), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n774), .B1(new_n856), .B2(new_n301), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n792), .A2(new_n344), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(G311), .B2(new_n820), .ZN(new_n859));
  INV_X1    g0659(.A(G294), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n859), .B1(new_n624), .B2(new_n796), .C1(new_n860), .C2(new_n797), .ZN(new_n861));
  INV_X1    g0661(.A(new_n807), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n862), .A2(G303), .B1(new_n789), .B2(G283), .ZN(new_n863));
  INV_X1    g0663(.A(new_n813), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n863), .B1(new_n207), .B2(new_n864), .ZN(new_n865));
  NOR4_X1   g0665(.A1(new_n861), .A2(new_n865), .A3(new_n406), .A4(new_n785), .ZN(new_n866));
  AOI22_X1  g0666(.A1(G137), .A2(new_n862), .B1(new_n817), .B2(G159), .ZN(new_n867));
  INV_X1    g0667(.A(G143), .ZN(new_n868));
  INV_X1    g0668(.A(G150), .ZN(new_n869));
  OAI221_X1 g0669(.A(new_n867), .B1(new_n868), .B2(new_n797), .C1(new_n869), .C2(new_n788), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT34), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n830), .B1(new_n792), .B2(new_n203), .ZN(new_n872));
  OAI22_X1  g0672(.A1(new_n864), .A2(new_n201), .B1(new_n202), .B2(new_n784), .ZN(new_n873));
  AOI211_X1 g0673(.A(new_n872), .B(new_n873), .C1(G132), .C2(new_n820), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n866), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n847), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n876), .B1(new_n429), .B2(new_n845), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n857), .B1(new_n875), .B2(new_n782), .C1(new_n877), .C2(new_n825), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n855), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(G384));
  NOR2_X1   g0680(.A1(new_n370), .A2(KEYINPUT16), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n342), .B1(new_n385), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n714), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(new_n402), .B2(new_n394), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT38), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n395), .B(new_n714), .C1(new_n324), .C2(new_n351), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n400), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT37), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n888), .A2(new_n889), .A3(new_n380), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n887), .A2(new_n882), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n380), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(KEYINPUT37), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  NOR3_X1   g0694(.A1(new_n885), .A2(new_n886), .A3(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n884), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n663), .B2(new_n672), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n890), .A2(new_n893), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT38), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n895), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n319), .A2(new_n716), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n667), .A2(new_n321), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n329), .A2(new_n319), .A3(new_n716), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n851), .B2(new_n876), .ZN(new_n905));
  OAI22_X1  g0705(.A1(new_n900), .A2(new_n905), .B1(new_n402), .B2(new_n883), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n886), .B1(new_n885), .B2(new_n894), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n897), .A2(KEYINPUT38), .A3(new_n898), .ZN(new_n908));
  AND3_X1   g0708(.A1(new_n907), .A2(KEYINPUT39), .A3(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n391), .A2(new_n714), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n402), .B2(new_n394), .ZN(new_n912));
  INV_X1    g0712(.A(new_n887), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n380), .B1(new_n391), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT99), .B1(new_n400), .B2(new_n887), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n914), .B1(new_n915), .B2(new_n889), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n888), .A2(KEYINPUT99), .A3(KEYINPUT37), .A4(new_n380), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n886), .B1(new_n912), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT39), .B1(new_n919), .B2(new_n908), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n909), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT98), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n667), .B2(new_n716), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n329), .A2(KEYINPUT98), .A3(new_n319), .A4(new_n723), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n906), .B1(new_n921), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n676), .B1(new_n748), .B2(new_n470), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n926), .B(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n664), .A2(new_n666), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n929), .A2(new_n901), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n330), .B2(new_n901), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n759), .A2(new_n716), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT31), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n759), .A2(KEYINPUT31), .A3(new_n716), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR3_X1   g0736(.A1(new_n661), .A2(new_n622), .A3(new_n716), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n877), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n931), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n895), .B2(new_n899), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT40), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n919), .B2(new_n908), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n940), .A2(new_n941), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n433), .B(new_n469), .C1(new_n937), .C2(new_n936), .ZN(new_n945));
  OAI21_X1  g0745(.A(G330), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(new_n945), .B2(new_n944), .ZN(new_n947));
  OAI22_X1  g0747(.A1(new_n928), .A2(new_n947), .B1(new_n275), .B2(new_n772), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(new_n928), .B2(new_n947), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n576), .A2(new_n577), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n950), .A2(KEYINPUT35), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(KEYINPUT35), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n951), .A2(G116), .A3(new_n231), .A4(new_n952), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n953), .B(KEYINPUT36), .Z(new_n954));
  OAI211_X1 g0754(.A(new_n233), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n201), .A2(G68), .ZN(new_n956));
  AOI211_X1 g0756(.A(new_n275), .B(G13), .C1(new_n955), .C2(new_n956), .ZN(new_n957));
  OR3_X1    g0757(.A1(new_n949), .A2(new_n954), .A3(new_n957), .ZN(G367));
  OAI21_X1  g0758(.A(new_n765), .B1(new_n559), .B2(new_n723), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n699), .A2(new_n582), .A3(new_n716), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n962), .A2(new_n731), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n964), .A2(KEYINPUT42), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n959), .A2(new_n655), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n716), .B1(new_n966), .B2(new_n583), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(new_n964), .B2(KEYINPUT42), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n513), .B1(new_n510), .B2(new_n723), .ZN(new_n969));
  OR3_X1    g0769(.A1(new_n679), .A2(new_n510), .A3(new_n723), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AOI22_X1  g0771(.A1(new_n965), .A2(new_n968), .B1(KEYINPUT43), .B2(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n972), .B(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n729), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n961), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n974), .B(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n734), .B(KEYINPUT41), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n731), .A2(KEYINPUT101), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n721), .B(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n728), .A2(new_n730), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(new_n981), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n731), .A2(new_n727), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n985), .A2(new_n962), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT45), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT44), .ZN(new_n988));
  INV_X1    g0788(.A(new_n985), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n988), .B1(new_n989), .B2(new_n961), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n985), .A2(KEYINPUT44), .A3(new_n962), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n990), .A2(KEYINPUT100), .A3(new_n991), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n987), .B(new_n992), .C1(KEYINPUT100), .C2(new_n990), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n975), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n993), .A2(new_n975), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n984), .A2(new_n770), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n978), .B1(new_n996), .B2(new_n770), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n773), .A2(G1), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n977), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n827), .B1(new_n221), .B2(new_n418), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(new_n244), .B2(new_n833), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n817), .A2(G283), .B1(G317), .B2(new_n820), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1002), .B1(new_n860), .B2(new_n788), .C1(new_n637), .C2(new_n797), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n813), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1004), .B1(new_n206), .B2(new_n792), .C1(new_n207), .C2(new_n784), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n803), .A2(new_n624), .ZN(new_n1006));
  INV_X1    g0806(.A(G311), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n831), .B1(new_n1006), .B2(KEYINPUT46), .C1(new_n807), .C2(new_n1007), .ZN(new_n1008));
  NOR3_X1   g0808(.A1(new_n1003), .A2(new_n1005), .A3(new_n1008), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n868), .A2(new_n807), .B1(new_n788), .B2(new_n800), .ZN(new_n1010));
  INV_X1    g0810(.A(G137), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n784), .A2(new_n203), .B1(new_n799), .B2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n796), .A2(new_n201), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n797), .A2(new_n869), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n792), .A2(new_n301), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n406), .B1(new_n803), .B2(new_n202), .ZN(new_n1017));
  NOR4_X1   g0817(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1009), .B1(new_n1013), .B2(new_n1018), .ZN(new_n1019));
  XOR2_X1   g0819(.A(KEYINPUT102), .B(KEYINPUT47), .Z(new_n1020));
  OR2_X1    g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n782), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n774), .B(new_n1001), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n841), .B2(new_n971), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n999), .A2(new_n1024), .ZN(G387));
  NAND2_X1  g0825(.A1(new_n984), .A2(new_n770), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n734), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n982), .A2(new_n769), .A3(new_n983), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n833), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n241), .A2(G45), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT103), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n415), .A2(new_n201), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT50), .Z(new_n1034));
  INV_X1    g0834(.A(new_n733), .ZN(new_n1035));
  AOI211_X1 g0835(.A(G45), .B(new_n1035), .C1(G68), .C2(G77), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n1030), .B(new_n1032), .C1(new_n1034), .C2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n836), .A2(new_n1035), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(G107), .B2(new_n221), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n827), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n815), .A2(new_n419), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n797), .B2(new_n201), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT105), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n830), .B1(new_n803), .B2(new_n301), .C1(new_n792), .C2(new_n206), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(KEYINPUT104), .B(G150), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n817), .A2(G68), .B1(new_n820), .B2(new_n1045), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n800), .B2(new_n807), .C1(new_n337), .C2(new_n788), .ZN(new_n1047));
  NOR3_X1   g0847(.A1(new_n1043), .A2(new_n1044), .A3(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n792), .A2(new_n624), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n831), .B1(new_n810), .B2(new_n799), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G303), .A2(new_n817), .B1(new_n862), .B2(G322), .ZN(new_n1051));
  INV_X1    g0851(.A(G317), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1051), .B1(new_n1007), .B2(new_n788), .C1(new_n1052), .C2(new_n797), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT48), .ZN(new_n1054));
  OR2_X1    g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1056));
  INV_X1    g0856(.A(G283), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n784), .A2(new_n1057), .B1(new_n860), .B2(new_n803), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT106), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1055), .A2(new_n1056), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1060), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n1049), .B(new_n1050), .C1(new_n1061), .C2(KEYINPUT49), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1061), .A2(KEYINPUT49), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1048), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1040), .B(new_n775), .C1(new_n782), .C2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n728), .A2(new_n841), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n984), .B2(new_n998), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1029), .A2(new_n1068), .ZN(G393));
  NAND3_X1  g0869(.A1(new_n995), .A2(new_n998), .A3(new_n994), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n961), .A2(new_n841), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT107), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n820), .A2(G322), .B1(G283), .B2(new_n804), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT108), .Z(new_n1074));
  OAI22_X1  g0874(.A1(new_n860), .A2(new_n796), .B1(new_n788), .B2(new_n637), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(G116), .B2(new_n815), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1074), .A2(new_n260), .A3(new_n794), .A4(new_n1076), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n1007), .A2(new_n797), .B1(new_n807), .B2(new_n1052), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT52), .Z(new_n1079));
  OAI22_X1  g0879(.A1(new_n869), .A2(new_n807), .B1(new_n797), .B2(new_n800), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT51), .Z(new_n1081));
  AOI211_X1 g0881(.A(new_n831), .B(new_n858), .C1(G68), .C2(new_n804), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n415), .A2(new_n817), .B1(G143), .B2(new_n820), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n789), .A2(G50), .B1(new_n815), .B2(G77), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n1077), .A2(new_n1079), .B1(new_n1081), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n781), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n827), .B1(new_n206), .B2(new_n221), .C1(new_n1030), .C2(new_n250), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1072), .A2(new_n775), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n995), .A2(new_n994), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1026), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n996), .A2(new_n1027), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1070), .B(new_n1089), .C1(new_n1092), .C2(new_n1093), .ZN(G390));
  NAND3_X1  g0894(.A1(new_n433), .A2(new_n469), .A3(new_n767), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n676), .B(new_n1095), .C1(new_n748), .C2(new_n470), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n931), .B1(new_n768), .B2(new_n848), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n767), .A2(new_n904), .A3(new_n877), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1097), .A2(KEYINPUT111), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n850), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n876), .B1(new_n707), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT111), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1103), .B(new_n931), .C1(new_n768), .C2(new_n848), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1099), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n723), .B(new_n846), .C1(new_n741), .C2(new_n743), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n847), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n768), .A2(new_n848), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n904), .A2(KEYINPUT109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT109), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n902), .A2(new_n1111), .A3(new_n903), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1098), .B(new_n1108), .C1(new_n1109), .C2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1096), .B1(new_n1105), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT110), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT39), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n916), .A2(new_n917), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n910), .B1(new_n663), .B2(new_n672), .ZN(new_n1120));
  AOI21_X1  g0920(.A(KEYINPUT38), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1118), .B1(new_n895), .B2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n907), .A2(KEYINPUT39), .A3(new_n908), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n925), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1122), .A2(new_n1123), .B1(new_n1124), .B2(new_n905), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n1110), .A2(new_n1112), .B1(new_n847), .B2(new_n1106), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1124), .B1(new_n895), .B2(new_n1121), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1117), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1124), .B1(new_n1101), .B2(new_n931), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n909), .B2(new_n920), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1112), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1111), .B1(new_n902), .B2(new_n903), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1107), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n925), .B1(new_n919), .B2(new_n908), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1131), .A2(new_n1136), .A3(KEYINPUT110), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1098), .B1(new_n1129), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1098), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1131), .A2(new_n1136), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1139), .B1(new_n1140), .B2(new_n1117), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1116), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n1131), .A2(KEYINPUT110), .A3(new_n1136), .ZN(new_n1143));
  AOI21_X1  g0943(.A(KEYINPUT110), .B1(new_n1131), .B2(new_n1136), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1139), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1129), .A2(new_n1098), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1145), .A2(new_n1146), .A3(new_n1115), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1142), .A2(new_n1147), .A3(new_n1027), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n824), .B1(new_n909), .B2(new_n920), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n804), .A2(new_n1045), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1150), .B(KEYINPUT53), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G125), .B2(new_n820), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(KEYINPUT54), .B(G143), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n817), .A2(new_n1154), .B1(G50), .B2(new_n793), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n260), .B(new_n1156), .C1(G159), .C2(new_n815), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n862), .A2(G128), .B1(new_n789), .B2(G137), .ZN(new_n1158));
  INV_X1    g0958(.A(G132), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1157), .B(new_n1158), .C1(new_n1159), .C2(new_n797), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n624), .A2(new_n797), .B1(new_n807), .B2(new_n1057), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(G107), .B2(new_n789), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n406), .B1(new_n793), .B2(G68), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n817), .A2(G97), .B1(new_n815), .B2(G77), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n813), .A2(G87), .B1(G294), .B2(new_n820), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .A4(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n782), .B1(new_n1160), .B2(new_n1166), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n774), .B(new_n1167), .C1(new_n337), .C2(new_n856), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1149), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT112), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1129), .A2(new_n1137), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1141), .B1(new_n1171), .B2(new_n1139), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1170), .B1(new_n1172), .B2(new_n998), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n998), .ZN(new_n1174));
  NOR4_X1   g0974(.A1(new_n1138), .A2(new_n1141), .A3(KEYINPUT112), .A4(new_n1174), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1148), .B(new_n1169), .C1(new_n1173), .C2(new_n1175), .ZN(G378));
  INV_X1    g0976(.A(new_n1096), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n919), .A2(new_n908), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n939), .A2(new_n1178), .A3(KEYINPUT40), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n848), .B1(new_n762), .B2(new_n766), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n904), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(new_n908), .B2(new_n907), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1179), .B(G330), .C1(new_n1182), .C2(KEYINPUT40), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n448), .B1(new_n673), .B2(new_n674), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n456), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1187), .A2(new_n714), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1185), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n469), .A2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1186), .A2(new_n1188), .A3(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n469), .A2(new_n1189), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n449), .B(new_n1185), .C1(new_n464), .C2(new_n468), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n1192), .A2(new_n1193), .B1(new_n1187), .B2(new_n714), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n1191), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1183), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1191), .A2(new_n1194), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n941), .B1(new_n900), .B2(new_n1181), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1197), .A2(new_n1198), .A3(G330), .A4(new_n1179), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT115), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1196), .B(new_n1199), .C1(new_n926), .C2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n921), .A2(new_n925), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n906), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1200), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1199), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1197), .B1(new_n943), .B2(G330), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1204), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n1147), .A2(new_n1177), .B1(new_n1201), .B2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(KEYINPUT116), .B1(new_n1208), .B2(KEYINPUT57), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT116), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT57), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1105), .A2(new_n1114), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1096), .B1(new_n1172), .B2(new_n1212), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1207), .A2(new_n1201), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1210), .B(new_n1211), .C1(new_n1213), .C2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1147), .A2(new_n1177), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n926), .B1(new_n1196), .B2(new_n1199), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1196), .A2(new_n1199), .A3(new_n926), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1211), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n734), .B1(new_n1216), .B2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1209), .A2(new_n1215), .A3(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1207), .A2(new_n1201), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1195), .A2(new_n824), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n819), .A2(G107), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(new_n1225), .B(KEYINPUT113), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n279), .B1(new_n803), .B2(new_n301), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n830), .B(new_n1227), .C1(new_n815), .C2(G68), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n807), .A2(new_n624), .B1(new_n1057), .B2(new_n799), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n792), .A2(new_n202), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n817), .A2(new_n419), .B1(new_n789), .B2(G97), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1226), .A2(new_n1228), .A3(new_n1231), .A4(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT58), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n279), .B1(new_n831), .B2(new_n278), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n1233), .A2(new_n1234), .B1(new_n201), .B2(new_n1235), .ZN(new_n1236));
  AOI211_X1 g1036(.A(G33), .B(G41), .C1(new_n793), .C2(G159), .ZN(new_n1237));
  INV_X1    g1037(.A(G124), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1237), .B1(new_n1238), .B2(new_n799), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1239), .B(KEYINPUT114), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n862), .A2(G125), .B1(new_n789), .B2(G132), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n817), .A2(G137), .B1(new_n819), .B2(G128), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n815), .A2(G150), .B1(new_n804), .B2(new_n1154), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1241), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(KEYINPUT59), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1240), .A2(new_n1245), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1244), .A2(KEYINPUT59), .ZN(new_n1247));
  OAI221_X1 g1047(.A(new_n1236), .B1(new_n1234), .B2(new_n1233), .C1(new_n1246), .C2(new_n1247), .ZN(new_n1248));
  AND2_X1   g1048(.A1(new_n1248), .A2(new_n781), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n774), .B(new_n1249), .C1(new_n201), .C2(new_n856), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n1223), .A2(new_n998), .B1(new_n1224), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1222), .A2(new_n1251), .ZN(G375));
  NAND2_X1  g1052(.A1(new_n1212), .A2(new_n998), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n774), .B1(new_n856), .B2(new_n203), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n864), .A2(new_n800), .B1(new_n788), .B2(new_n1153), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n819), .A2(G137), .B1(G128), .B2(new_n820), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1256), .B(new_n830), .C1(new_n202), .C2(new_n792), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n1255), .B(new_n1257), .C1(G132), .C2(new_n862), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n796), .A2(new_n869), .B1(new_n784), .B2(new_n201), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1259), .B(KEYINPUT117), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n788), .A2(new_n624), .B1(new_n637), .B2(new_n799), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1261), .B1(G294), .B2(new_n862), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n864), .A2(new_n206), .B1(new_n207), .B2(new_n796), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1041), .B1(new_n797), .B2(new_n1057), .ZN(new_n1264));
  NOR4_X1   g1064(.A1(new_n1263), .A2(new_n1264), .A3(new_n406), .A4(new_n1016), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n1258), .A2(new_n1260), .B1(new_n1262), .B2(new_n1265), .ZN(new_n1266));
  OAI221_X1 g1066(.A(new_n1254), .B1(new_n782), .B2(new_n1266), .C1(new_n1113), .C2(new_n825), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1253), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n978), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1105), .A2(new_n1096), .A3(new_n1114), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1116), .A2(new_n1270), .A3(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1269), .A2(new_n1272), .ZN(G381));
  INV_X1    g1073(.A(G387), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1029), .A2(new_n843), .A3(new_n1068), .ZN(new_n1275));
  NOR3_X1   g1075(.A1(G390), .A2(G384), .A3(new_n1275), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1274), .A2(new_n1276), .A3(new_n1269), .A4(new_n1272), .ZN(new_n1277));
  XOR2_X1   g1077(.A(new_n1277), .B(KEYINPUT118), .Z(new_n1278));
  NOR2_X1   g1078(.A1(G375), .A2(G378), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(G407));
  NAND2_X1  g1080(.A1(new_n715), .A2(G213), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1279), .A2(new_n1282), .ZN(new_n1283));
  XNOR2_X1  g1083(.A(new_n1283), .B(KEYINPUT119), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(G407), .A2(G213), .A3(new_n1284), .ZN(G409));
  INV_X1    g1085(.A(KEYINPUT63), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT122), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT120), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n1196), .A2(new_n926), .A3(new_n1199), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n998), .B1(new_n1289), .B2(new_n1217), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1224), .A2(new_n1250), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1292), .B1(new_n1208), .B2(new_n1270), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1288), .B1(new_n1293), .B2(G378), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1216), .A2(new_n1270), .A3(new_n1223), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  AND2_X1   g1097(.A1(new_n1148), .A2(new_n1169), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1175), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1300));
  OAI21_X1  g1100(.A(KEYINPUT112), .B1(new_n1300), .B2(new_n1174), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1299), .A2(new_n1301), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1297), .A2(new_n1298), .A3(KEYINPUT120), .A4(new_n1302), .ZN(new_n1303));
  AND2_X1   g1103(.A1(new_n1294), .A2(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1222), .A2(G378), .A3(new_n1251), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1282), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT60), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1271), .A2(new_n1307), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1308), .A2(new_n734), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1271), .B1(new_n1115), .B2(new_n1307), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(KEYINPUT121), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT121), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1309), .A2(new_n1313), .A3(new_n1310), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1312), .A2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(new_n1269), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n879), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1315), .A2(G384), .A3(new_n1269), .ZN(new_n1318));
  AND2_X1   g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1287), .B1(new_n1306), .B2(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1305), .A2(new_n1294), .A3(new_n1303), .ZN(new_n1321));
  AND4_X1   g1121(.A1(new_n1287), .A2(new_n1321), .A3(new_n1281), .A4(new_n1319), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1286), .B1(new_n1320), .B2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(G390), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1275), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n843), .B1(new_n1029), .B2(new_n1068), .ZN(new_n1326));
  OAI21_X1  g1126(.A(KEYINPUT123), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1326), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT123), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1328), .A2(new_n1329), .A3(new_n1275), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1327), .A2(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(KEYINPUT124), .B1(new_n999), .B2(new_n1024), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  AOI22_X1  g1133(.A1(new_n1327), .A2(new_n1330), .B1(new_n999), .B2(new_n1024), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1324), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  OAI211_X1 g1135(.A(new_n1327), .B(new_n1330), .C1(new_n1274), .C2(KEYINPUT124), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1331), .A2(G387), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1336), .A2(new_n1337), .A3(G390), .ZN(new_n1338));
  AOI21_X1  g1138(.A(KEYINPUT61), .B1(new_n1335), .B2(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(G2897), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1319), .B1(new_n1340), .B2(new_n1281), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1321), .A2(new_n1281), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1343), .A2(G2897), .A3(new_n1282), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1341), .A2(new_n1342), .A3(new_n1344), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1306), .A2(KEYINPUT63), .A3(new_n1319), .ZN(new_n1346));
  NAND4_X1  g1146(.A1(new_n1323), .A2(new_n1339), .A3(new_n1345), .A4(new_n1346), .ZN(new_n1347));
  XOR2_X1   g1147(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n1348));
  NAND2_X1  g1148(.A1(new_n1345), .A2(new_n1348), .ZN(new_n1349));
  XOR2_X1   g1149(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1350));
  OAI21_X1  g1150(.A(new_n1350), .B1(new_n1320), .B2(new_n1322), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1306), .A2(KEYINPUT62), .A3(new_n1319), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1349), .B1(new_n1351), .B2(new_n1352), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1335), .A2(new_n1338), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1347), .B1(new_n1353), .B2(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1355), .A2(KEYINPUT127), .ZN(new_n1356));
  INV_X1    g1156(.A(KEYINPUT127), .ZN(new_n1357));
  OAI211_X1 g1157(.A(new_n1347), .B(new_n1357), .C1(new_n1353), .C2(new_n1354), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1356), .A2(new_n1358), .ZN(G405));
  XNOR2_X1  g1159(.A(G375), .B(G378), .ZN(new_n1360));
  XNOR2_X1  g1160(.A(new_n1360), .B(new_n1319), .ZN(new_n1361));
  XNOR2_X1  g1161(.A(new_n1361), .B(new_n1354), .ZN(G402));
endmodule


