//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0 0 1 0 0 1 1 1 0 0 0 1 0 0 0 1 1 1 0 1 1 0 0 1 1 0 1 1 0 1 1 1 0 1 0 0 0 1 0 1 0 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n566, new_n567, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n577, new_n578, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1140, new_n1141, new_n1142,
    new_n1143;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  INV_X1    g023(.A(G2106), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT67), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n453), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n458), .A2(new_n455), .B1(new_n453), .B2(new_n449), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT68), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  AOI22_X1  g036(.A1(new_n461), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT69), .B(G2105), .ZN(new_n463));
  OAI21_X1  g038(.A(KEYINPUT70), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT71), .B(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n467), .B1(new_n468), .B2(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT69), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT69), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  AND3_X1   g048(.A1(new_n471), .A2(new_n473), .A3(G137), .ZN(new_n474));
  INV_X1    g049(.A(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT71), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT71), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(G2105), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  AOI22_X1  g054(.A1(new_n469), .A2(new_n474), .B1(G101), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n475), .A2(KEYINPUT3), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n466), .A2(new_n481), .A3(G125), .ZN(new_n482));
  NAND2_X1  g057(.A1(G113), .A2(G2104), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n463), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AND3_X1   g061(.A1(new_n464), .A2(new_n480), .A3(new_n486), .ZN(G160));
  NAND3_X1  g062(.A1(new_n476), .A2(new_n478), .A3(KEYINPUT3), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(new_n466), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT72), .ZN(new_n490));
  OR3_X1    g065(.A1(new_n489), .A2(new_n490), .A3(new_n463), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n489), .B2(new_n463), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G124), .ZN(new_n494));
  XNOR2_X1  g069(.A(new_n494), .B(KEYINPUT73), .ZN(new_n495));
  OAI221_X1 g070(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n463), .C2(G112), .ZN(new_n496));
  XNOR2_X1  g071(.A(new_n496), .B(KEYINPUT74), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n469), .A2(new_n470), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n499), .A2(G136), .ZN(new_n500));
  NOR3_X1   g075(.A1(new_n495), .A2(new_n497), .A3(new_n500), .ZN(G162));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n471), .A2(new_n473), .A3(G138), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n466), .A2(new_n481), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OR2_X1    g080(.A1(G102), .A2(G2105), .ZN(new_n506));
  OAI211_X1 g081(.A(new_n506), .B(G2104), .C1(G114), .C2(new_n470), .ZN(new_n507));
  AND2_X1   g082(.A1(G126), .A2(G2105), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT4), .A2(G138), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n508), .B1(new_n463), .B2(new_n509), .ZN(new_n510));
  OAI211_X1 g085(.A(new_n505), .B(new_n507), .C1(new_n489), .C2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(G164));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  OAI21_X1  g088(.A(KEYINPUT77), .B1(new_n513), .B2(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT77), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n515), .A2(new_n516), .A3(G543), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n514), .A2(new_n517), .B1(KEYINPUT5), .B2(new_n513), .ZN(new_n518));
  AND2_X1   g093(.A1(new_n518), .A2(G62), .ZN(new_n519));
  AND2_X1   g094(.A1(G75), .A2(G543), .ZN(new_n520));
  OAI21_X1  g095(.A(G651), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT6), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT75), .ZN(new_n524));
  OR3_X1    g099(.A1(new_n522), .A2(KEYINPUT76), .A3(KEYINPUT6), .ZN(new_n525));
  OAI21_X1  g100(.A(KEYINPUT76), .B1(new_n522), .B2(KEYINPUT6), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n524), .A2(G88), .A3(new_n518), .A4(new_n527), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n524), .A2(G50), .A3(G543), .A4(new_n527), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n521), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(G166));
  OR2_X1    g106(.A1(new_n523), .A2(KEYINPUT75), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n523), .A2(KEYINPUT75), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n532), .A2(new_n533), .B1(new_n525), .B2(new_n526), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n534), .A2(G89), .A3(new_n518), .ZN(new_n535));
  XNOR2_X1  g110(.A(KEYINPUT79), .B(KEYINPUT7), .ZN(new_n536));
  AND3_X1   g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n536), .A2(new_n537), .ZN(new_n539));
  AND2_X1   g114(.A1(G63), .A2(G651), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n538), .A2(new_n539), .B1(new_n518), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n535), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n524), .A2(G543), .A3(new_n527), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT78), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT78), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n534), .A2(new_n545), .A3(G543), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n542), .B1(new_n547), .B2(G51), .ZN(G168));
  INV_X1    g123(.A(G90), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n524), .A2(new_n518), .A3(new_n527), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n551));
  OAI22_X1  g126(.A1(new_n549), .A2(new_n550), .B1(new_n551), .B2(new_n522), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  AND2_X1   g128(.A1(new_n544), .A2(new_n546), .ZN(new_n554));
  INV_X1    g129(.A(G52), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(G301));
  INV_X1    g131(.A(G301), .ZN(G171));
  INV_X1    g132(.A(G43), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n558), .B1(new_n544), .B2(new_n546), .ZN(new_n559));
  INV_X1    g134(.A(G81), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n518), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n561));
  OAI22_X1  g136(.A1(new_n560), .A2(new_n550), .B1(new_n561), .B2(new_n522), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  NAND4_X1  g143(.A1(new_n524), .A2(G53), .A3(G543), .A4(new_n527), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n569), .B(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(G91), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n518), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n573));
  OAI22_X1  g148(.A1(new_n572), .A2(new_n550), .B1(new_n573), .B2(new_n522), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G299));
  INV_X1    g151(.A(new_n542), .ZN(new_n577));
  INV_X1    g152(.A(G51), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n554), .B2(new_n578), .ZN(G286));
  INV_X1    g154(.A(KEYINPUT80), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n521), .A2(new_n580), .A3(new_n528), .A4(new_n529), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n528), .A2(new_n529), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n520), .B1(new_n518), .B2(G62), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n522), .ZN(new_n584));
  OAI21_X1  g159(.A(KEYINPUT80), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  AND2_X1   g160(.A1(new_n581), .A2(new_n585), .ZN(G303));
  AND3_X1   g161(.A1(new_n524), .A2(new_n518), .A3(new_n527), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(G87), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n534), .A2(G49), .A3(G543), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(G288));
  AOI22_X1  g166(.A1(new_n518), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n522), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n587), .A2(G86), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n534), .A2(G48), .A3(G543), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(G305));
  NAND2_X1  g172(.A1(G72), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(new_n518), .ZN(new_n599));
  INV_X1    g174(.A(G60), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT81), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n522), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(new_n602), .B2(new_n601), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n547), .A2(G47), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n587), .A2(G85), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(G290));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  NOR2_X1   g183(.A1(G301), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n587), .A2(KEYINPUT10), .A3(G92), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  INV_X1    g186(.A(G92), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n550), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(G79), .A2(G543), .ZN(new_n614));
  INV_X1    g189(.A(G66), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n599), .B2(new_n615), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n610), .A2(new_n613), .B1(G651), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n547), .A2(G54), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT82), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n609), .B1(new_n620), .B2(new_n608), .ZN(G284));
  XOR2_X1   g196(.A(G284), .B(KEYINPUT83), .Z(G321));
  NAND2_X1  g197(.A1(G286), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n575), .ZN(G297));
  OAI21_X1  g199(.A(new_n623), .B1(G868), .B2(new_n575), .ZN(G280));
  INV_X1    g200(.A(KEYINPUT82), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n619), .B(new_n626), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n627), .A2(G559), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(G860), .B2(new_n620), .ZN(G148));
  INV_X1    g204(.A(new_n563), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(new_n608), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(new_n628), .B2(new_n608), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g208(.A1(new_n479), .A2(new_n461), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT12), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2100), .Z(new_n637));
  NAND2_X1  g212(.A1(new_n493), .A2(G123), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n499), .A2(G135), .ZN(new_n639));
  OAI221_X1 g214(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n463), .C2(G111), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n641), .A2(G2096), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(G2096), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n637), .A2(new_n642), .A3(new_n643), .ZN(G156));
  XNOR2_X1  g219(.A(G2427), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(KEYINPUT14), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n650), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2451), .B(G2454), .Z(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(G14), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n654), .A2(new_n657), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(G401));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT85), .Z(new_n664));
  AOI21_X1  g239(.A(new_n662), .B1(new_n664), .B2(KEYINPUT86), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n665), .B1(KEYINPUT86), .B2(new_n664), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2084), .B(G2090), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n664), .B(KEYINPUT17), .Z(new_n668));
  INV_X1    g243(.A(new_n662), .ZN(new_n669));
  OAI211_X1 g244(.A(new_n666), .B(new_n667), .C1(new_n668), .C2(new_n669), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n669), .A2(new_n667), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n664), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT18), .Z(new_n673));
  NOR2_X1   g248(.A1(new_n662), .A2(new_n667), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n668), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n670), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2096), .B(G2100), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G227));
  XOR2_X1   g253(.A(G1971), .B(G1976), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1956), .B(G2474), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1961), .B(G1966), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n681), .A2(new_n682), .ZN(new_n684));
  NOR3_X1   g259(.A1(new_n680), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n680), .A2(new_n683), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT20), .Z(new_n687));
  AOI211_X1 g262(.A(new_n685), .B(new_n687), .C1(new_n680), .C2(new_n684), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1991), .B(G1996), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1981), .B(G1986), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(G229));
  INV_X1    g270(.A(G16), .ZN(new_n696));
  NOR2_X1   g271(.A1(G171), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(G5), .B2(new_n696), .ZN(new_n698));
  INV_X1    g273(.A(G1961), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT24), .ZN(new_n701));
  INV_X1    g276(.A(G34), .ZN(new_n702));
  AOI21_X1  g277(.A(G29), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(new_n701), .B2(new_n702), .ZN(new_n704));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n704), .B1(G160), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT26), .Z(new_n708));
  NAND2_X1  g283(.A1(new_n479), .A2(G105), .ZN(new_n709));
  INV_X1    g284(.A(G141), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n708), .B(new_n709), .C1(new_n498), .C2(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(new_n493), .B2(G129), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n712), .A2(new_n705), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(new_n705), .B2(G32), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT27), .B(G1996), .ZN(new_n715));
  OAI221_X1 g290(.A(new_n700), .B1(G2084), .B2(new_n706), .C1(new_n714), .C2(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT92), .ZN(new_n717));
  NOR2_X1   g292(.A1(G29), .A2(G33), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT90), .Z(new_n719));
  NAND3_X1  g294(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT91), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT25), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n499), .A2(G139), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n722), .B(new_n723), .C1(new_n463), .C2(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n719), .B1(new_n725), .B2(new_n705), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G2072), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n696), .A2(G21), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G168), .B2(new_n696), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n727), .B1(G1966), .B2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT31), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(G11), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(G11), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT30), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n734), .A2(G28), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n705), .B1(new_n734), .B2(G28), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n732), .B(new_n733), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(G164), .A2(G29), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G27), .B2(G29), .ZN(new_n739));
  INV_X1    g314(.A(G2078), .ZN(new_n740));
  OAI22_X1  g315(.A1(new_n641), .A2(new_n705), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AOI211_X1 g316(.A(new_n737), .B(new_n741), .C1(new_n740), .C2(new_n739), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n705), .A2(G26), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT28), .ZN(new_n744));
  OAI221_X1 g319(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n463), .C2(G116), .ZN(new_n745));
  INV_X1    g320(.A(G140), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n745), .B1(new_n498), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n493), .B2(G128), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n744), .B1(new_n748), .B2(new_n705), .ZN(new_n749));
  INV_X1    g324(.A(G2067), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n706), .A2(G2084), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n742), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n714), .A2(new_n715), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n729), .A2(G1966), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n754), .B(new_n755), .C1(new_n699), .C2(new_n698), .ZN(new_n756));
  NOR2_X1   g331(.A1(G16), .A2(G19), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n563), .B2(G16), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT89), .B(G1341), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NOR4_X1   g335(.A1(new_n730), .A2(new_n753), .A3(new_n756), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n705), .A2(G35), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G162), .B2(new_n705), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT29), .Z(new_n764));
  INV_X1    g339(.A(G2090), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(G4), .A2(G16), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n620), .B2(G16), .ZN(new_n768));
  INV_X1    g343(.A(G1348), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n717), .A2(new_n761), .A3(new_n766), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n696), .A2(G20), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT23), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n575), .B2(new_n696), .ZN(new_n774));
  INV_X1    g349(.A(G1956), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n764), .B2(new_n765), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n777), .A2(KEYINPUT93), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n777), .A2(KEYINPUT93), .ZN(new_n779));
  NOR3_X1   g354(.A1(new_n771), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n696), .A2(G22), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G166), .B2(new_n696), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1971), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n696), .A2(G23), .ZN(new_n785));
  AND3_X1   g360(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n785), .B1(new_n786), .B2(new_n696), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT33), .B(G1976), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n787), .B(new_n788), .Z(new_n789));
  MUX2_X1   g364(.A(G6), .B(G305), .S(G16), .Z(new_n790));
  XOR2_X1   g365(.A(KEYINPUT32), .B(G1981), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT87), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n790), .A2(new_n792), .ZN(new_n794));
  AOI211_X1 g369(.A(new_n784), .B(new_n789), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT34), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n696), .A2(G24), .ZN(new_n798));
  INV_X1    g373(.A(G290), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(new_n696), .ZN(new_n800));
  INV_X1    g375(.A(G1986), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n705), .A2(G25), .ZN(new_n803));
  OAI221_X1 g378(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n463), .C2(G107), .ZN(new_n804));
  INV_X1    g379(.A(G131), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n498), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n493), .B2(G119), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n803), .B1(new_n807), .B2(new_n705), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT35), .B(G1991), .Z(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n797), .A2(new_n802), .A3(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT88), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n795), .A2(new_n796), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(KEYINPUT36), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT36), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n812), .A2(new_n817), .A3(new_n814), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n781), .B1(new_n816), .B2(new_n818), .ZN(G311));
  NAND2_X1  g394(.A1(new_n816), .A2(new_n818), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(new_n780), .ZN(G150));
  NAND2_X1  g396(.A1(new_n620), .A2(G559), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT38), .ZN(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT94), .B(G55), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(new_n544), .B2(new_n546), .ZN(new_n826));
  INV_X1    g401(.A(G93), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n828));
  OAI22_X1  g403(.A1(new_n827), .A2(new_n550), .B1(new_n828), .B2(new_n522), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n563), .A2(new_n830), .ZN(new_n831));
  OAI22_X1  g406(.A1(new_n559), .A2(new_n562), .B1(new_n826), .B2(new_n829), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n823), .B(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT39), .ZN(new_n835));
  AOI21_X1  g410(.A(G860), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(new_n835), .B2(new_n834), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT95), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(G860), .B1(new_n826), .B2(new_n829), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT96), .B(KEYINPUT37), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n839), .A2(new_n842), .ZN(G145));
  INV_X1    g418(.A(G37), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n748), .B(G164), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(new_n712), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n725), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n807), .B(new_n635), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n463), .A2(G118), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT98), .ZN(new_n850));
  OAI21_X1  g425(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n850), .B2(new_n851), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT97), .ZN(new_n854));
  AND3_X1   g429(.A1(new_n499), .A2(new_n854), .A3(G142), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n854), .B1(new_n499), .B2(G142), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n853), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n857), .B1(G130), .B2(new_n493), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n848), .B(new_n858), .Z(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(KEYINPUT100), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n847), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n847), .A2(new_n860), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n641), .B(G160), .ZN(new_n863));
  XNOR2_X1  g438(.A(G162), .B(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n847), .A2(new_n859), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT99), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n865), .B1(new_n847), .B2(new_n859), .ZN(new_n869));
  AND3_X1   g444(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n868), .B1(new_n867), .B2(new_n869), .ZN(new_n871));
  OAI221_X1 g446(.A(new_n844), .B1(new_n861), .B2(new_n866), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g448(.A(new_n628), .B(new_n833), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n619), .A2(new_n575), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT41), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n617), .B(new_n618), .C1(new_n571), .C2(new_n574), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n875), .A2(KEYINPUT101), .A3(new_n877), .ZN(new_n880));
  OR3_X1    g455(.A1(new_n619), .A2(new_n575), .A3(KEYINPUT101), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n879), .B1(new_n882), .B2(KEYINPUT41), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n874), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n885), .B1(new_n874), .B2(new_n882), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n886), .A2(KEYINPUT42), .ZN(new_n887));
  XNOR2_X1  g462(.A(G290), .B(G305), .ZN(new_n888));
  XNOR2_X1  g463(.A(G288), .B(new_n530), .ZN(new_n889));
  XOR2_X1   g464(.A(new_n888), .B(new_n889), .Z(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n891), .A2(KEYINPUT102), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n886), .A2(KEYINPUT42), .ZN(new_n893));
  AND3_X1   g468(.A1(new_n887), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n892), .B1(new_n887), .B2(new_n893), .ZN(new_n895));
  OAI21_X1  g470(.A(G868), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n896), .B1(G868), .B2(new_n830), .ZN(G295));
  OAI21_X1  g472(.A(new_n896), .B1(G868), .B2(new_n830), .ZN(G331));
  INV_X1    g473(.A(KEYINPUT103), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n553), .B(new_n899), .C1(new_n554), .C2(new_n555), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n555), .B1(new_n544), .B2(new_n546), .ZN(new_n901));
  OAI21_X1  g476(.A(KEYINPUT103), .B1(new_n901), .B2(new_n552), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n900), .A2(G168), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(G301), .A2(G286), .A3(KEYINPUT103), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(KEYINPUT104), .B1(new_n905), .B2(new_n833), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n831), .A2(new_n832), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT104), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n907), .A2(new_n908), .A3(new_n904), .A4(new_n903), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n905), .A2(new_n833), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n906), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT105), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n880), .A2(new_n881), .A3(new_n876), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n875), .A2(KEYINPUT41), .A3(new_n877), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n911), .A2(new_n912), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n912), .B1(new_n911), .B2(new_n915), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n882), .A2(new_n910), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n905), .A2(new_n833), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR3_X1   g495(.A1(new_n916), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(KEYINPUT106), .B1(new_n921), .B2(new_n891), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n911), .A2(new_n915), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT105), .ZN(new_n925));
  INV_X1    g500(.A(new_n920), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n923), .B(new_n890), .C1(new_n927), .C2(new_n916), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n905), .B(new_n833), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n883), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n882), .A2(new_n906), .A3(new_n910), .A4(new_n909), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n844), .B1(new_n932), .B2(new_n890), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n922), .A2(new_n928), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT43), .ZN(new_n936));
  INV_X1    g511(.A(new_n932), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n934), .B1(new_n891), .B2(new_n937), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n936), .B(KEYINPUT44), .C1(KEYINPUT43), .C2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n922), .A2(new_n928), .A3(new_n941), .A4(new_n934), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n937), .A2(new_n891), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT43), .B1(new_n943), .B2(new_n933), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n940), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AOI211_X1 g522(.A(KEYINPUT107), .B(KEYINPUT44), .C1(new_n942), .C2(new_n944), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n939), .B1(new_n947), .B2(new_n948), .ZN(G397));
  XOR2_X1   g524(.A(KEYINPUT108), .B(G40), .Z(new_n950));
  NAND4_X1  g525(.A1(new_n464), .A2(new_n480), .A3(new_n486), .A4(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G1384), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n511), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(G8), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(G86), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n596), .B1(new_n958), .B2(new_n550), .ZN(new_n959));
  OAI21_X1  g534(.A(G1981), .B1(new_n959), .B2(new_n593), .ZN(new_n960));
  INV_X1    g535(.A(G1981), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n594), .A2(new_n595), .A3(new_n961), .A4(new_n596), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT49), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n963), .A2(new_n956), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n960), .A2(new_n962), .A3(KEYINPUT49), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT114), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n965), .A2(new_n966), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n964), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(G1976), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n969), .A2(new_n970), .A3(new_n786), .ZN(new_n971));
  INV_X1    g546(.A(new_n962), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n957), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n974));
  NOR2_X1   g549(.A1(G288), .A2(new_n970), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n974), .B1(new_n956), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n786), .A2(G1976), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n977), .A2(KEYINPUT112), .A3(G8), .A4(new_n955), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n976), .A2(KEYINPUT52), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT52), .B1(G288), .B2(new_n970), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT113), .ZN(new_n981));
  OR2_X1    g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n981), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n982), .A2(new_n957), .A3(new_n977), .A4(new_n983), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n969), .A2(new_n979), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n953), .A2(KEYINPUT50), .ZN(new_n986));
  AND4_X1   g561(.A1(new_n486), .A2(new_n464), .A3(new_n480), .A4(new_n950), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT50), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n511), .A2(new_n988), .A3(new_n952), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n986), .A2(new_n987), .A3(new_n765), .A4(new_n989), .ZN(new_n990));
  AND3_X1   g565(.A1(new_n511), .A2(KEYINPUT45), .A3(new_n952), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT45), .B1(new_n511), .B2(new_n952), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n991), .A2(new_n992), .A3(new_n951), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n990), .B1(new_n993), .B2(G1971), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT110), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n581), .A2(new_n585), .A3(G8), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n581), .A2(new_n585), .A3(KEYINPUT55), .A4(G8), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT110), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n990), .B(new_n1001), .C1(new_n993), .C2(G1971), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n995), .A2(G8), .A3(new_n1000), .A4(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT111), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G8), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1006), .B1(new_n994), .B2(KEYINPUT110), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1007), .A2(KEYINPUT111), .A3(new_n1000), .A4(new_n1002), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n985), .A2(new_n1005), .A3(new_n1008), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n973), .A2(new_n1009), .A3(KEYINPUT115), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT115), .B1(new_n973), .B2(new_n1009), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n994), .A2(G8), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1014), .A2(new_n998), .A3(new_n999), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n986), .A2(new_n987), .A3(new_n989), .ZN(new_n1016));
  OAI22_X1  g591(.A1(new_n993), .A2(G1966), .B1(new_n1016), .B2(G2084), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1017), .A2(G8), .A3(G168), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1013), .A2(new_n1015), .A3(new_n985), .A4(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT63), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1020), .A2(KEYINPUT116), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1000), .B1(new_n1007), .B2(new_n1002), .ZN(new_n1023));
  NOR3_X1   g598(.A1(new_n1023), .A2(new_n1021), .A3(new_n1018), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1024), .A2(new_n1013), .A3(new_n985), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT117), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT117), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1024), .A2(new_n1013), .A3(new_n1027), .A4(new_n985), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1022), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT116), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1012), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT118), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT118), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1012), .B(new_n1033), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1034));
  AND2_X1   g609(.A1(new_n1017), .A2(G286), .ZN(new_n1035));
  OAI21_X1  g610(.A(G8), .B1(new_n1017), .B2(G286), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT51), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1037), .B1(KEYINPUT51), .B2(new_n1036), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT119), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1016), .A2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n986), .A2(new_n987), .A3(KEYINPUT119), .A4(new_n989), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(new_n699), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n993), .A2(new_n740), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n993), .A2(KEYINPUT53), .A3(new_n740), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1042), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(G171), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n1048), .B(KEYINPUT122), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1038), .B1(new_n1049), .B2(KEYINPUT62), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1013), .A2(new_n1015), .A3(new_n985), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1053));
  XNOR2_X1  g628(.A(KEYINPUT56), .B(G2072), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n993), .A2(new_n1054), .ZN(new_n1055));
  OR3_X1    g630(.A1(new_n571), .A2(KEYINPUT57), .A3(new_n574), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1016), .A2(new_n775), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n954), .A2(new_n750), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1040), .A2(new_n769), .A3(new_n1041), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n627), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1053), .A2(new_n1056), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1058), .B1(new_n1061), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  OAI211_X1 g643(.A(KEYINPUT120), .B(new_n1058), .C1(new_n1061), .C2(new_n1065), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1064), .A2(new_n1058), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT61), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT60), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n627), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n620), .A2(KEYINPUT60), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1074), .A2(new_n1075), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1060), .A2(new_n1059), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1077), .A2(KEYINPUT60), .A3(new_n620), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1064), .A2(KEYINPUT61), .A3(new_n1058), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1072), .A2(new_n1076), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G1996), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n993), .A2(new_n1081), .ZN(new_n1082));
  OR2_X1    g657(.A1(new_n1082), .A2(KEYINPUT121), .ZN(new_n1083));
  XOR2_X1   g658(.A(KEYINPUT58), .B(G1341), .Z(new_n1084));
  AOI22_X1  g659(.A1(new_n1082), .A2(KEYINPUT121), .B1(new_n955), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n630), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n1086), .B(KEYINPUT59), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1068), .B(new_n1069), .C1(new_n1080), .C2(new_n1087), .ZN(new_n1088));
  OR2_X1    g663(.A1(new_n1047), .A2(G171), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n991), .A2(new_n992), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n480), .A2(KEYINPUT123), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n480), .A2(KEYINPUT123), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n740), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1093), .A2(new_n484), .A3(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1091), .A2(new_n1092), .A3(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1042), .A2(new_n1045), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1090), .B1(new_n1097), .B2(G171), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1089), .A2(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n1099), .B(KEYINPUT124), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1097), .A2(G171), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1090), .B1(new_n1049), .B2(new_n1101), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1088), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT62), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1049), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n1038), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1052), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1032), .A2(new_n1034), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n992), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1109), .A2(new_n951), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n807), .B(new_n809), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1111), .B(KEYINPUT109), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n748), .B(G2067), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n712), .B(G1996), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  OR2_X1    g690(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g691(.A(G290), .B(G1986), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1110), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1108), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1116), .A2(new_n1110), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n799), .A2(new_n801), .A3(new_n1110), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1121), .B(KEYINPUT48), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n748), .A2(new_n750), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n807), .A2(new_n809), .ZN(new_n1124));
  XOR2_X1   g699(.A(new_n1124), .B(KEYINPUT125), .Z(new_n1125));
  OAI21_X1  g700(.A(new_n1123), .B1(new_n1125), .B2(new_n1115), .ZN(new_n1126));
  AOI22_X1  g701(.A1(new_n1120), .A2(new_n1122), .B1(new_n1110), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1081), .A2(KEYINPUT46), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1113), .A2(new_n712), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1110), .ZN(new_n1130));
  AOI21_X1  g705(.A(KEYINPUT46), .B1(new_n1110), .B2(new_n1081), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT126), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1134));
  OAI22_X1  g709(.A1(new_n1129), .A2(new_n1130), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1135), .B(KEYINPUT47), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1127), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1119), .A2(new_n1137), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g713(.A(G319), .B1(new_n659), .B2(new_n660), .ZN(new_n1140));
  OAI21_X1  g714(.A(KEYINPUT127), .B1(G227), .B2(new_n1140), .ZN(new_n1141));
  OR3_X1    g715(.A1(G227), .A2(KEYINPUT127), .A3(new_n1140), .ZN(new_n1142));
  AND3_X1   g716(.A1(new_n694), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  NAND3_X1  g717(.A1(new_n1143), .A2(new_n872), .A3(new_n945), .ZN(G225));
  INV_X1    g718(.A(G225), .ZN(G308));
endmodule


