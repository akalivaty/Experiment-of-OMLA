//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 0 1 1 0 0 1 1 0 1 1 0 1 0 0 0 1 1 1 0 0 1 1 0 0 1 1 1 0 0 0 0 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  NAND3_X1  g001(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT22), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(G137), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  XOR2_X1   g005(.A(G119), .B(G128), .Z(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT24), .B(G110), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT16), .ZN(new_n195));
  INV_X1    g009(.A(G140), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(new_n196), .A3(G125), .ZN(new_n197));
  XOR2_X1   g011(.A(G125), .B(G140), .Z(new_n198));
  OAI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(new_n195), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  OAI211_X1 g015(.A(G146), .B(new_n197), .C1(new_n198), .C2(new_n195), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n194), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT78), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n206));
  INV_X1    g020(.A(G119), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(G128), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT77), .B1(new_n207), .B2(G128), .ZN(new_n209));
  XNOR2_X1  g023(.A(new_n208), .B(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n205), .B1(new_n210), .B2(G110), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(G110), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(KEYINPUT78), .ZN(new_n213));
  NOR3_X1   g027(.A1(new_n204), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n192), .A2(new_n193), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT79), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n192), .A2(new_n193), .A3(KEYINPUT79), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n217), .B(new_n218), .C1(new_n210), .C2(G110), .ZN(new_n219));
  XNOR2_X1  g033(.A(G125), .B(G140), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(new_n200), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n219), .A2(new_n202), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n191), .B1(new_n214), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G902), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n213), .A2(new_n211), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n203), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(new_n222), .A3(new_n190), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n224), .A2(new_n225), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT25), .ZN(new_n230));
  INV_X1    g044(.A(G217), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n231), .B1(G234), .B2(new_n225), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT25), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n224), .A2(new_n233), .A3(new_n225), .A4(new_n228), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n230), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n232), .A2(G902), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n224), .A2(new_n228), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G469), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n187), .A2(G227), .ZN(new_n240));
  XNOR2_X1  g054(.A(new_n240), .B(new_n196), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n241), .B(KEYINPUT81), .ZN(new_n242));
  XOR2_X1   g056(.A(new_n242), .B(G110), .Z(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT86), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT65), .B1(new_n200), .B2(G143), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT65), .ZN(new_n247));
  INV_X1    g061(.A(G143), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(new_n248), .A3(G146), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G128), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n200), .A2(G143), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n251), .B1(new_n252), .B2(KEYINPUT1), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n250), .A2(new_n253), .A3(new_n252), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT85), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n250), .A2(new_n252), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n248), .A2(G146), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT1), .ZN(new_n258));
  OAI21_X1  g072(.A(G128), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n257), .B1(new_n246), .B2(new_n249), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT85), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n261), .A2(new_n262), .A3(new_n253), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n255), .A2(new_n260), .A3(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT83), .B(G101), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT82), .ZN(new_n266));
  INV_X1    g080(.A(G104), .ZN(new_n267));
  AOI22_X1  g081(.A1(new_n266), .A2(KEYINPUT3), .B1(new_n267), .B2(G107), .ZN(new_n268));
  OAI22_X1  g082(.A1(new_n266), .A2(KEYINPUT3), .B1(new_n267), .B2(G107), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT3), .ZN(new_n270));
  INV_X1    g084(.A(G107), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n270), .A2(new_n271), .A3(KEYINPUT82), .A4(G104), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n265), .A2(new_n268), .A3(new_n269), .A4(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n271), .A2(G104), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n267), .A2(G107), .ZN(new_n275));
  OAI21_X1  g089(.A(G101), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n264), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT10), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n245), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI211_X1 g094(.A(KEYINPUT86), .B(KEYINPUT10), .C1(new_n264), .C2(new_n277), .ZN(new_n281));
  OR2_X1    g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT11), .ZN(new_n283));
  INV_X1    g097(.A(G134), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n283), .B1(new_n284), .B2(G137), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(G137), .ZN(new_n286));
  INV_X1    g100(.A(G137), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n287), .A2(KEYINPUT11), .A3(G134), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n285), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT67), .ZN(new_n290));
  XNOR2_X1  g104(.A(KEYINPUT66), .B(G131), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n289), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n285), .A2(new_n286), .A3(new_n288), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT67), .B1(new_n294), .B2(new_n291), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n293), .A2(new_n295), .B1(G131), .B2(new_n294), .ZN(new_n296));
  NAND2_X1  g110(.A1(KEYINPUT0), .A2(G128), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT64), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n297), .B(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(KEYINPUT0), .A2(G128), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n248), .A2(G146), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n301), .B1(new_n252), .B2(new_n302), .ZN(new_n303));
  AOI22_X1  g117(.A1(new_n298), .A2(new_n261), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n268), .A2(new_n269), .A3(new_n272), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT84), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(new_n306), .A3(G101), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT4), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n305), .A2(new_n306), .A3(KEYINPUT4), .A4(G101), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n273), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n304), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n252), .A2(new_n302), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n259), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n254), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n277), .A2(KEYINPUT10), .A3(new_n316), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n282), .A2(new_n296), .A3(new_n313), .A4(new_n317), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n313), .B(new_n317), .C1(new_n280), .C2(new_n281), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n294), .A2(G131), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n290), .B1(new_n289), .B2(new_n292), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n294), .A2(KEYINPUT67), .A3(new_n291), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n244), .B1(new_n318), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT12), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n277), .A2(new_n316), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n327), .B1(new_n277), .B2(new_n264), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n326), .B1(new_n328), .B2(new_n296), .ZN(new_n329));
  INV_X1    g143(.A(new_n278), .ZN(new_n330));
  OAI211_X1 g144(.A(KEYINPUT12), .B(new_n323), .C1(new_n330), .C2(new_n327), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n332), .B(new_n244), .C1(new_n319), .C2(new_n323), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n239), .B(new_n225), .C1(new_n325), .C2(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n239), .A2(new_n225), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n318), .A2(new_n324), .A3(new_n244), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n332), .B1(new_n319), .B2(new_n323), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n243), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(new_n340), .A3(G469), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n335), .A2(new_n337), .A3(new_n341), .ZN(new_n342));
  XOR2_X1   g156(.A(KEYINPUT9), .B(G234), .Z(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n225), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n344), .A2(G221), .ZN(new_n345));
  XOR2_X1   g159(.A(new_n345), .B(KEYINPUT80), .Z(new_n346));
  OAI21_X1  g160(.A(G214), .B1(G237), .B2(G902), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  XOR2_X1   g162(.A(G110), .B(G122), .Z(new_n349));
  OAI21_X1  g163(.A(KEYINPUT68), .B1(new_n207), .B2(G116), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT68), .ZN(new_n351));
  INV_X1    g165(.A(G116), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(new_n352), .A3(G119), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n207), .A2(G116), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  XOR2_X1   g170(.A(KEYINPUT2), .B(G113), .Z(new_n357));
  XNOR2_X1  g171(.A(new_n356), .B(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n312), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n358), .B1(new_n359), .B2(new_n309), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n354), .A2(KEYINPUT5), .A3(new_n355), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n361), .B(G113), .C1(KEYINPUT5), .C2(new_n355), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n357), .A2(new_n354), .A3(new_n355), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n277), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n349), .B1(new_n360), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n358), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n368), .B1(new_n310), .B2(new_n312), .ZN(new_n369));
  AND2_X1   g183(.A1(new_n362), .A2(new_n363), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n277), .ZN(new_n371));
  INV_X1    g185(.A(new_n349), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n369), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n367), .A2(new_n373), .A3(KEYINPUT6), .ZN(new_n374));
  MUX2_X1   g188(.A(new_n316), .B(new_n304), .S(G125), .Z(new_n375));
  NAND2_X1  g189(.A1(new_n187), .A2(G224), .ZN(new_n376));
  XOR2_X1   g190(.A(new_n376), .B(KEYINPUT87), .Z(new_n377));
  XOR2_X1   g191(.A(new_n375), .B(new_n377), .Z(new_n378));
  INV_X1    g192(.A(KEYINPUT6), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n379), .B(new_n349), .C1(new_n360), .C2(new_n366), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n374), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n300), .A2(new_n303), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n382), .B1(new_n297), .B2(new_n256), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G125), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT7), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n377), .A2(new_n385), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n384), .B(new_n386), .C1(G125), .C2(new_n316), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT89), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n387), .B(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT88), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n390), .B1(new_n364), .B2(new_n365), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n371), .A2(new_n391), .ZN(new_n392));
  XOR2_X1   g206(.A(new_n349), .B(KEYINPUT8), .Z(new_n393));
  NAND3_X1  g207(.A1(new_n370), .A2(new_n390), .A3(new_n277), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  OR2_X1    g209(.A1(new_n375), .A2(new_n386), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n389), .A2(new_n395), .A3(new_n373), .A4(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n381), .A2(new_n397), .A3(new_n225), .ZN(new_n398));
  OAI21_X1  g212(.A(G210), .B1(G237), .B2(G902), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n381), .A2(new_n397), .A3(new_n225), .A4(new_n399), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n348), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G237), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(new_n187), .A3(G214), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n405), .B(new_n248), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(KEYINPUT17), .A3(new_n291), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(new_n201), .A3(new_n202), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT91), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n406), .A2(new_n291), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n405), .B(G143), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n292), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT17), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n410), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT91), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n407), .A2(new_n201), .A3(new_n415), .A4(new_n202), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n409), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(G113), .B(G122), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(new_n267), .ZN(new_n419));
  NAND2_X1  g233(.A1(KEYINPUT18), .A2(G131), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n406), .B(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n198), .A2(G146), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n221), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n417), .A2(new_n419), .A3(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n419), .B1(new_n417), .B2(new_n424), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n225), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(G475), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n352), .A2(G122), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n430), .B(KEYINPUT14), .ZN(new_n431));
  OAI21_X1  g245(.A(KEYINPUT92), .B1(new_n352), .B2(G122), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT92), .ZN(new_n433));
  INV_X1    g247(.A(G122), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(new_n434), .A3(G116), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(G107), .B1(new_n431), .B2(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(G128), .B(G143), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(new_n284), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n436), .A2(new_n271), .A3(new_n430), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n438), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n284), .B1(new_n439), .B2(KEYINPUT13), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n248), .A2(G128), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n443), .B1(KEYINPUT13), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n441), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n271), .B1(new_n436), .B2(new_n430), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n439), .A2(new_n284), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(KEYINPUT93), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n442), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n343), .A2(G217), .A3(new_n187), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(KEYINPUT94), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT93), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n449), .B(new_n455), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n456), .B(new_n445), .C1(new_n446), .C2(new_n447), .ZN(new_n457));
  XOR2_X1   g271(.A(new_n452), .B(KEYINPUT94), .Z(new_n458));
  NAND3_X1  g272(.A1(new_n457), .A2(new_n458), .A3(new_n442), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n454), .A2(new_n459), .A3(new_n225), .ZN(new_n460));
  INV_X1    g274(.A(G478), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(KEYINPUT15), .ZN(new_n462));
  OR2_X1    g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n460), .A2(new_n462), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n187), .A2(G952), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n465), .B1(G234), .B2(G237), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  XOR2_X1   g281(.A(KEYINPUT21), .B(G898), .Z(new_n468));
  NAND2_X1  g282(.A1(G234), .A2(G237), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(G902), .A3(G953), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n467), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n463), .A2(new_n464), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n410), .A2(new_n412), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n198), .A2(KEYINPUT19), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT19), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n220), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n474), .A2(new_n200), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n477), .A2(KEYINPUT90), .A3(new_n202), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT90), .B1(new_n477), .B2(new_n202), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n424), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n419), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(G475), .B1(new_n425), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT20), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n485), .A3(new_n225), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n485), .B1(new_n484), .B2(new_n225), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n429), .B(new_n472), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n342), .A2(new_n346), .A3(new_n403), .A4(new_n490), .ZN(new_n491));
  XOR2_X1   g305(.A(KEYINPUT75), .B(KEYINPUT32), .Z(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT74), .ZN(new_n494));
  NOR2_X1   g308(.A1(G472), .A2(G902), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n287), .A2(G134), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n286), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n498), .A2(G131), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n316), .B(new_n500), .C1(new_n321), .C2(new_n322), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n293), .A2(new_n295), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n383), .B1(new_n503), .B2(new_n320), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT30), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT30), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n501), .B(new_n506), .C1(new_n296), .C2(new_n383), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n358), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n501), .B(new_n358), .C1(new_n296), .C2(new_n383), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n404), .A2(new_n187), .A3(G210), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(KEYINPUT70), .ZN(new_n511));
  XOR2_X1   g325(.A(KEYINPUT26), .B(G101), .Z(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OR2_X1    g327(.A1(new_n510), .A2(KEYINPUT70), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n510), .A2(KEYINPUT70), .ZN(new_n515));
  INV_X1    g329(.A(new_n512), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n513), .A2(new_n517), .A3(new_n519), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n509), .A2(new_n523), .A3(KEYINPUT71), .ZN(new_n524));
  AOI21_X1  g338(.A(KEYINPUT71), .B1(new_n509), .B2(new_n523), .ZN(new_n525));
  NOR3_X1   g339(.A1(new_n508), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT31), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT72), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n507), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n323), .A2(new_n304), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n506), .B1(new_n530), .B2(new_n501), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n368), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n509), .A2(new_n523), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT71), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n509), .A2(new_n523), .A3(KEYINPUT71), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n532), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT72), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(new_n538), .A3(KEYINPUT31), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n528), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n509), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n541), .A2(KEYINPUT28), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n499), .B1(new_n293), .B2(new_n295), .ZN(new_n544));
  AOI22_X1  g358(.A1(new_n323), .A2(new_n304), .B1(new_n544), .B2(new_n316), .ZN(new_n545));
  OAI21_X1  g359(.A(KEYINPUT73), .B1(new_n545), .B2(new_n358), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT73), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n547), .B(new_n368), .C1(new_n502), .C2(new_n504), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n541), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT28), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n543), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n523), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n551), .A2(new_n552), .B1(new_n526), .B2(new_n527), .ZN(new_n553));
  AOI211_X1 g367(.A(new_n494), .B(new_n496), .C1(new_n540), .C2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n526), .A2(new_n527), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n551), .A2(new_n552), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n537), .A2(new_n538), .A3(KEYINPUT31), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n538), .B1(new_n537), .B2(KEYINPUT31), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n555), .B(new_n556), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(KEYINPUT74), .B1(new_n559), .B2(new_n495), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n493), .B1(new_n554), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n496), .B1(new_n540), .B2(new_n553), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n523), .B(new_n543), .C1(new_n549), .C2(new_n550), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT29), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n532), .A2(new_n509), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n552), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n368), .B1(new_n502), .B2(new_n504), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n509), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT28), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n543), .A2(new_n570), .A3(KEYINPUT29), .A4(new_n523), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT76), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n542), .B1(KEYINPUT28), .B2(new_n569), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n574), .A2(KEYINPUT76), .A3(KEYINPUT29), .A4(new_n523), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n567), .A2(new_n225), .A3(new_n573), .A4(new_n575), .ZN(new_n576));
  AOI22_X1  g390(.A1(new_n562), .A2(KEYINPUT32), .B1(new_n576), .B2(G472), .ZN(new_n577));
  AOI211_X1 g391(.A(new_n238), .B(new_n491), .C1(new_n561), .C2(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(new_n265), .ZN(G3));
  NAND2_X1  g393(.A1(new_n403), .A2(new_n471), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n559), .A2(new_n495), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n494), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n562), .A2(KEYINPUT74), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n557), .A2(new_n558), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n556), .A2(new_n555), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n225), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g400(.A1(new_n582), .A2(new_n583), .B1(G472), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n238), .ZN(new_n588));
  INV_X1    g402(.A(new_n346), .ZN(new_n589));
  INV_X1    g403(.A(new_n319), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n243), .B1(new_n590), .B2(new_n296), .ZN(new_n591));
  AOI22_X1  g405(.A1(new_n591), .A2(new_n324), .B1(new_n243), .B2(new_n339), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n336), .B1(new_n592), .B2(G469), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n589), .B1(new_n593), .B2(new_n335), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n587), .A2(new_n588), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n580), .B1(new_n595), .B2(KEYINPUT95), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n596), .B1(KEYINPUT95), .B2(new_n595), .ZN(new_n597));
  INV_X1    g411(.A(new_n488), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n598), .A2(new_n486), .B1(G475), .B2(new_n428), .ZN(new_n599));
  OAI21_X1  g413(.A(KEYINPUT33), .B1(new_n453), .B2(KEYINPUT96), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n454), .A2(new_n601), .A3(new_n459), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n601), .B1(new_n454), .B2(new_n459), .ZN(new_n604));
  OAI211_X1 g418(.A(G478), .B(new_n225), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT97), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n460), .A2(new_n461), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n454), .A2(new_n459), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n600), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n602), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n611), .A2(KEYINPUT97), .A3(G478), .A4(new_n225), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n607), .A2(new_n608), .A3(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT98), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n607), .A2(KEYINPUT98), .A3(new_n608), .A4(new_n612), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n599), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n597), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT34), .B(G104), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G6));
  NAND2_X1  g435(.A1(new_n463), .A2(new_n464), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT99), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n598), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n624), .A2(new_n486), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n487), .B1(new_n598), .B2(new_n623), .ZN(new_n626));
  OAI211_X1 g440(.A(new_n429), .B(new_n622), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n597), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(KEYINPUT35), .B(G107), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G9));
  INV_X1    g444(.A(new_n587), .ZN(new_n631));
  OAI21_X1  g445(.A(KEYINPUT100), .B1(new_n214), .B2(new_n223), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n191), .A2(KEYINPUT36), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT100), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n227), .A2(new_n634), .A3(new_n222), .ZN(new_n635));
  AND3_X1   g449(.A1(new_n632), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n633), .B1(new_n632), .B2(new_n635), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n236), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n638), .A2(KEYINPUT101), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n638), .A2(KEYINPUT101), .ZN(new_n640));
  INV_X1    g454(.A(new_n235), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n631), .A2(new_n491), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT37), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G110), .ZN(G12));
  NAND2_X1  g459(.A1(new_n561), .A2(new_n577), .ZN(new_n646));
  OR3_X1    g460(.A1(new_n470), .A2(KEYINPUT102), .A3(G900), .ZN(new_n647));
  OAI21_X1  g461(.A(KEYINPUT102), .B1(new_n470), .B2(G900), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n647), .A2(new_n467), .A3(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n627), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n594), .A2(new_n403), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n642), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n646), .A2(new_n651), .A3(new_n653), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G128), .ZN(G30));
  INV_X1    g470(.A(new_n622), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n599), .A2(new_n657), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n642), .A2(new_n347), .A3(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT103), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n523), .B1(new_n568), .B2(new_n509), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n225), .B1(new_n526), .B2(new_n662), .ZN(new_n663));
  AOI22_X1  g477(.A1(new_n562), .A2(KEYINPUT32), .B1(G472), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n561), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n665), .B1(new_n659), .B2(new_n660), .ZN(new_n666));
  XOR2_X1   g480(.A(new_n649), .B(KEYINPUT39), .Z(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n594), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT40), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n401), .A2(new_n402), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n671), .B(KEYINPUT38), .Z(new_n672));
  NOR4_X1   g486(.A1(new_n661), .A2(new_n666), .A3(new_n670), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(new_n248), .ZN(G45));
  NAND2_X1  g488(.A1(new_n617), .A2(new_n649), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n646), .A2(new_n653), .A3(new_n654), .A4(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n652), .B1(new_n561), .B2(new_n577), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n680), .A2(KEYINPUT104), .A3(new_n654), .A4(new_n676), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G146), .ZN(G48));
  AOI21_X1  g497(.A(new_n238), .B1(new_n561), .B2(new_n577), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n319), .A2(new_n323), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n319), .A2(new_n323), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n243), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n333), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(G469), .B1(new_n689), .B2(G902), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n335), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n691), .A2(new_n345), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n671), .A2(new_n347), .A3(new_n471), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n617), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n684), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT41), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G113), .ZN(G15));
  INV_X1    g512(.A(new_n345), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n690), .A2(new_n699), .A3(new_n335), .A4(new_n403), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n700), .A2(new_n627), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n646), .A2(new_n701), .A3(new_n588), .A4(new_n471), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT105), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G116), .ZN(G18));
  NOR2_X1   g518(.A1(new_n700), .A2(new_n642), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n646), .A2(new_n705), .A3(new_n490), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G119), .ZN(G21));
  NAND2_X1  g521(.A1(new_n238), .A2(KEYINPUT107), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT107), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n235), .A2(new_n709), .A3(new_n237), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT106), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n574), .B(new_n713), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n555), .B1(new_n714), .B2(new_n523), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n526), .A2(new_n527), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n495), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n586), .A2(G472), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n712), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n690), .A2(new_n658), .A3(new_n699), .A4(new_n335), .ZN(new_n720));
  OR3_X1    g534(.A1(new_n719), .A2(new_n580), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G122), .ZN(G24));
  NAND2_X1  g536(.A1(new_n717), .A2(new_n718), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n723), .A2(new_n675), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n705), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G125), .ZN(G27));
  NOR2_X1   g540(.A1(new_n671), .A2(new_n348), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n675), .A2(KEYINPUT42), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n345), .B1(new_n593), .B2(new_n335), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n684), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n675), .A2(new_n728), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT32), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n581), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n577), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(KEYINPUT108), .B1(new_n735), .B2(new_n712), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT108), .ZN(new_n737));
  AOI211_X1 g551(.A(new_n737), .B(new_n711), .C1(new_n577), .C2(new_n734), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n730), .B(new_n732), .C1(new_n736), .C2(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n731), .B1(new_n739), .B2(KEYINPUT42), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G131), .ZN(G33));
  NAND4_X1  g555(.A1(new_n684), .A2(new_n651), .A3(new_n730), .A4(new_n727), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G134), .ZN(G36));
  NAND2_X1  g557(.A1(new_n615), .A2(new_n616), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n599), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT43), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n747), .A2(new_n631), .A3(new_n654), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(KEYINPUT109), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n748), .A2(new_n749), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT46), .ZN(new_n753));
  XOR2_X1   g567(.A(new_n592), .B(KEYINPUT45), .Z(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(G469), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n753), .B1(new_n756), .B2(new_n336), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n755), .A2(KEYINPUT46), .A3(new_n337), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(new_n335), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n699), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n667), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n751), .A2(new_n727), .A3(new_n752), .A4(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G137), .ZN(G39));
  INV_X1    g577(.A(KEYINPUT47), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n759), .A2(KEYINPUT47), .A3(new_n699), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n646), .A2(new_n588), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(new_n732), .A3(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G140), .ZN(G42));
  XNOR2_X1  g584(.A(new_n691), .B(KEYINPUT49), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n771), .A2(new_n589), .A3(new_n745), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n665), .A2(new_n348), .A3(new_n711), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n672), .A3(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n655), .A2(new_n725), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n730), .A2(new_n649), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n665), .A2(new_n671), .A3(new_n659), .A4(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n682), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n776), .B1(new_n679), .B2(new_n681), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(KEYINPUT52), .A3(new_n779), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n739), .A2(KEYINPUT42), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n696), .A2(new_n721), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n702), .A2(new_n706), .ZN(new_n789));
  INV_X1    g603(.A(new_n731), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n787), .A2(new_n788), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n599), .A2(new_n622), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(KEYINPUT111), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n595), .A2(new_n580), .A3(new_n794), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n594), .B(new_n718), .C1(new_n560), .C2(new_n554), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n796), .A2(new_n238), .A3(new_n694), .ZN(new_n797));
  OAI21_X1  g611(.A(KEYINPUT110), .B1(new_n578), .B2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n491), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n646), .A2(new_n588), .A3(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n695), .A2(new_n587), .A3(new_n588), .A4(new_n594), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT110), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  AOI211_X1 g617(.A(new_n643), .B(new_n795), .C1(new_n798), .C2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n624), .B(new_n486), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n622), .A2(new_n650), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n805), .A2(new_n429), .A3(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT112), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n805), .A2(KEYINPUT112), .A3(new_n429), .A4(new_n806), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n809), .A2(new_n646), .A3(new_n594), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n724), .A2(new_n730), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n813), .A2(new_n654), .A3(new_n727), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n792), .A2(new_n742), .A3(new_n804), .A4(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n775), .B1(new_n786), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT113), .ZN(new_n817));
  AOI21_X1  g631(.A(KEYINPUT52), .B1(new_n783), .B2(new_n779), .ZN(new_n818));
  AND4_X1   g632(.A1(KEYINPUT52), .A2(new_n682), .A3(new_n777), .A4(new_n779), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT115), .ZN(new_n821));
  OAI21_X1  g635(.A(KEYINPUT53), .B1(new_n791), .B2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n782), .A2(KEYINPUT113), .A3(new_n784), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n643), .B1(new_n798), .B2(new_n803), .ZN(new_n825));
  INV_X1    g639(.A(new_n795), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n825), .A2(new_n742), .A3(new_n826), .A4(new_n814), .ZN(new_n827));
  AND4_X1   g641(.A1(new_n696), .A2(new_n702), .A3(new_n721), .A4(new_n706), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT115), .B1(new_n740), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n820), .A2(new_n823), .A3(new_n824), .A4(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n816), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n798), .A2(new_n803), .ZN(new_n834));
  INV_X1    g648(.A(new_n643), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n834), .A2(new_n835), .A3(new_n742), .A4(new_n826), .ZN(new_n836));
  INV_X1    g650(.A(new_n814), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n836), .A2(new_n791), .A3(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n820), .A2(new_n838), .A3(new_n824), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT114), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n839), .A2(new_n840), .A3(new_n775), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n840), .B1(new_n839), .B2(new_n775), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n786), .A2(new_n815), .A3(new_n775), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n833), .B1(new_n844), .B2(new_n832), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n747), .A2(new_n466), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n846), .B(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n848), .A2(new_n719), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n672), .A2(new_n348), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n849), .A2(new_n692), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT50), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n849), .A2(KEYINPUT50), .A3(new_n692), .A4(new_n850), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n691), .A2(new_n346), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n849), .B(new_n727), .C1(new_n767), .C2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n692), .A2(new_n727), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n858), .A2(new_n238), .ZN(new_n859));
  INV_X1    g673(.A(new_n665), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n859), .A2(new_n466), .A3(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n862), .A2(new_n599), .A3(new_n615), .A4(new_n616), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n848), .A2(new_n858), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n864), .A2(new_n718), .A3(new_n654), .A4(new_n717), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n855), .A2(new_n857), .A3(new_n863), .A4(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT51), .ZN(new_n867));
  OR2_X1    g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n849), .A2(new_n403), .A3(new_n692), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT48), .ZN(new_n870));
  OR2_X1    g684(.A1(new_n736), .A2(new_n738), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n864), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n870), .B1(new_n864), .B2(new_n871), .ZN(new_n873));
  OAI22_X1  g687(.A1(new_n872), .A2(new_n873), .B1(new_n618), .B2(new_n861), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n874), .B1(new_n866), .B2(new_n867), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n868), .A2(new_n869), .A3(new_n875), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n465), .B(KEYINPUT117), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n845), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(G952), .A2(G953), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n774), .B1(new_n878), .B2(new_n879), .ZN(G75));
  NAND2_X1  g694(.A1(new_n816), .A2(new_n831), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n881), .A2(G210), .A3(G902), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n882), .A2(KEYINPUT56), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n374), .A2(new_n380), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(new_n378), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT55), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n883), .B(new_n886), .C1(KEYINPUT118), .C2(new_n882), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n886), .B1(new_n882), .B2(KEYINPUT118), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n888), .B1(KEYINPUT56), .B2(new_n882), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n187), .A2(G952), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n887), .A2(new_n889), .A3(new_n891), .ZN(G51));
  XNOR2_X1  g706(.A(new_n336), .B(KEYINPUT57), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n881), .A2(KEYINPUT54), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n894), .B1(new_n895), .B2(new_n833), .ZN(new_n896));
  OAI21_X1  g710(.A(KEYINPUT119), .B1(new_n896), .B2(new_n689), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT53), .B1(new_n838), .B2(new_n785), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n782), .A2(KEYINPUT113), .A3(new_n784), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT113), .B1(new_n782), .B2(new_n784), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n822), .A2(new_n827), .A3(new_n829), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n898), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n903), .A2(new_n225), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n756), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n816), .A2(new_n831), .A3(new_n832), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n832), .B1(new_n816), .B2(new_n831), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n893), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT119), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n908), .A2(new_n909), .A3(new_n688), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n897), .A2(new_n905), .A3(new_n910), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n911), .A2(new_n891), .ZN(G54));
  NAND3_X1  g726(.A1(new_n904), .A2(KEYINPUT58), .A3(G475), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n913), .A2(new_n483), .A3(new_n425), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n913), .B1(new_n483), .B2(new_n425), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n914), .A2(new_n915), .A3(new_n890), .ZN(G60));
  NAND2_X1  g730(.A1(G478), .A2(G902), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT59), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n611), .B1(new_n845), .B2(new_n918), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n611), .B(new_n918), .C1(new_n906), .C2(new_n907), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n920), .A2(KEYINPUT120), .A3(new_n891), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT120), .B1(new_n920), .B2(new_n891), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n919), .A2(new_n921), .A3(new_n922), .ZN(G63));
  INV_X1    g737(.A(KEYINPUT122), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(KEYINPUT61), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n891), .B1(new_n924), .B2(KEYINPUT61), .ZN(new_n926));
  NAND2_X1  g740(.A1(G217), .A2(G902), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT60), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT121), .B1(new_n903), .B2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT121), .ZN(new_n930));
  INV_X1    g744(.A(new_n928), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n881), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  OR2_X1    g747(.A1(new_n636), .A2(new_n637), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n926), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n224), .A2(new_n228), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n929), .A2(new_n936), .A3(new_n932), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n925), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n930), .B1(new_n881), .B2(new_n931), .ZN(new_n939));
  AOI211_X1 g753(.A(KEYINPUT121), .B(new_n928), .C1(new_n816), .C2(new_n831), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n934), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n926), .ZN(new_n942));
  AND4_X1   g756(.A1(new_n925), .A2(new_n941), .A3(new_n937), .A4(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n938), .A2(new_n943), .ZN(G66));
  AOI21_X1  g758(.A(new_n187), .B1(new_n468), .B2(G224), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n804), .A2(new_n828), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n945), .B1(new_n946), .B2(new_n187), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n884), .B1(G898), .B2(new_n187), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT123), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n947), .B(new_n949), .ZN(G69));
  NOR2_X1   g764(.A1(new_n529), .A2(new_n531), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n474), .A2(new_n476), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT124), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n951), .B(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n761), .A2(new_n403), .A3(new_n658), .A4(new_n871), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n762), .A2(new_n740), .A3(new_n769), .A4(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n783), .A2(new_n742), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n955), .B1(new_n959), .B2(new_n187), .ZN(new_n960));
  INV_X1    g774(.A(G900), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n960), .B1(new_n961), .B2(new_n187), .ZN(new_n962));
  INV_X1    g776(.A(G227), .ZN(new_n963));
  OAI21_X1  g777(.A(G953), .B1(new_n963), .B2(new_n961), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT126), .ZN(new_n965));
  OR2_X1    g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n783), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n967), .A2(new_n673), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT62), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n794), .A2(new_n618), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n970), .A2(KEYINPUT125), .ZN(new_n971));
  NOR3_X1   g785(.A1(new_n971), .A2(new_n669), .A3(new_n728), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n970), .A2(KEYINPUT125), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n972), .A2(new_n684), .A3(new_n973), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n969), .A2(new_n762), .A3(new_n769), .A4(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n187), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n955), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n962), .A2(new_n966), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n964), .A2(new_n965), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n978), .B(new_n979), .ZN(G72));
  NAND2_X1  g794(.A1(G472), .A2(G902), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT63), .Z(new_n982));
  OAI21_X1  g796(.A(new_n982), .B1(new_n975), .B2(new_n946), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n565), .B(KEYINPUT127), .Z(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n983), .A2(new_n523), .A3(new_n985), .ZN(new_n986));
  NOR3_X1   g800(.A1(new_n957), .A2(new_n946), .A3(new_n958), .ZN(new_n987));
  INV_X1    g801(.A(new_n982), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n552), .B(new_n984), .C1(new_n987), .C2(new_n988), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n986), .A2(new_n891), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n844), .B1(new_n537), .B2(new_n566), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n990), .B1(new_n991), .B2(new_n982), .ZN(G57));
endmodule


