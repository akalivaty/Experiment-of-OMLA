//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 0 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 1 0 1 1 1 1 0 0 0 0 1 1 0 1 0 1 0 0 0 0 1 0 0 1 0 1 1 0 1 0 0 1 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:15 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027;
  NAND2_X1  g000(.A1(G234), .A2(G237), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  AND3_X1   g002(.A1(new_n187), .A2(G952), .A3(new_n188), .ZN(new_n189));
  AND3_X1   g003(.A1(new_n187), .A2(G902), .A3(G953), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT21), .B(G898), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n189), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  OAI21_X1  g006(.A(G214), .B1(G237), .B2(G902), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  OAI21_X1  g008(.A(G210), .B1(G237), .B2(G902), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(G143), .B(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(KEYINPUT0), .A2(G128), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT65), .B1(new_n201), .B2(G146), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT65), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(new_n204), .A3(G143), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n201), .A2(G146), .ZN(new_n206));
  AND3_X1   g020(.A1(new_n202), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(KEYINPUT0), .A3(G128), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT0), .ZN(new_n210));
  INV_X1    g024(.A(G128), .ZN(new_n211));
  AOI21_X1  g025(.A(KEYINPUT64), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n209), .B1(new_n212), .B2(new_n199), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n200), .B1(new_n207), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G125), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT89), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n211), .A2(KEYINPUT1), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n204), .A2(G143), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n218), .A3(new_n206), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT66), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT66), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n197), .A2(new_n221), .A3(new_n217), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n211), .B1(new_n218), .B2(KEYINPUT1), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n202), .A2(new_n205), .A3(new_n206), .ZN(new_n225));
  AOI22_X1  g039(.A1(new_n220), .A2(new_n222), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G125), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT89), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n214), .A2(new_n229), .A3(G125), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n216), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n188), .A2(G224), .ZN(new_n232));
  XNOR2_X1  g046(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(G110), .B(G122), .ZN(new_n234));
  INV_X1    g048(.A(G107), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT79), .B1(new_n235), .B2(G104), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT79), .ZN(new_n237));
  INV_X1    g051(.A(G104), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n237), .A2(new_n238), .A3(G107), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n235), .A2(KEYINPUT3), .A3(G104), .ZN(new_n240));
  AOI21_X1  g054(.A(KEYINPUT3), .B1(new_n235), .B2(G104), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n236), .B(new_n239), .C1(new_n240), .C2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G101), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT3), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n244), .B1(new_n238), .B2(G107), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n235), .A2(KEYINPUT3), .A3(G104), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G101), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n247), .A2(new_n248), .A3(new_n236), .A4(new_n239), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n243), .A2(KEYINPUT4), .A3(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT80), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n253), .B1(new_n242), .B2(G101), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(KEYINPUT80), .A3(new_n249), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT67), .ZN(new_n258));
  INV_X1    g072(.A(G119), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(KEYINPUT67), .A2(G119), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(G116), .A3(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n259), .A2(G116), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G113), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT2), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT2), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G113), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n262), .A2(new_n264), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n269), .B1(new_n262), .B2(new_n264), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n257), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n269), .ZN(new_n273));
  AND2_X1   g087(.A1(KEYINPUT67), .A2(G119), .ZN(new_n274));
  NOR2_X1   g088(.A1(KEYINPUT67), .A2(G119), .ZN(new_n275));
  INV_X1    g089(.A(G116), .ZN(new_n276));
  NOR3_X1   g090(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n273), .B1(new_n277), .B2(new_n263), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n262), .A2(new_n264), .A3(new_n269), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n278), .A2(new_n279), .A3(KEYINPUT68), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n242), .A2(new_n253), .A3(G101), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n272), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n256), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(KEYINPUT85), .B(KEYINPUT5), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n265), .B1(new_n277), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n262), .A2(new_n264), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n286), .B1(new_n287), .B2(new_n285), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n279), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT82), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT81), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n292), .B1(new_n238), .B2(G107), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n238), .A2(G107), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n235), .A2(KEYINPUT81), .A3(G104), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G101), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n249), .A2(new_n291), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n291), .B1(new_n249), .B2(new_n297), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n290), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n234), .B1(new_n284), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT6), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT88), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT88), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n302), .A2(new_n306), .A3(new_n303), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT87), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT86), .ZN(new_n309));
  INV_X1    g123(.A(new_n234), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n282), .B1(new_n252), .B2(new_n255), .ZN(new_n311));
  NOR3_X1   g125(.A1(new_n289), .A2(new_n298), .A3(new_n299), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n309), .B(new_n310), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n284), .A2(new_n301), .A3(new_n234), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(KEYINPUT6), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n284), .A2(new_n301), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n309), .B1(new_n316), .B2(new_n310), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n308), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  AOI22_X1  g132(.A1(new_n256), .A2(new_n283), .B1(new_n290), .B2(new_n300), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT86), .B1(new_n319), .B2(new_n234), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n303), .B1(new_n319), .B2(new_n234), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n320), .A2(new_n321), .A3(KEYINPUT87), .A4(new_n313), .ZN(new_n322));
  AOI221_X4 g136(.A(new_n233), .B1(new_n305), .B2(new_n307), .C1(new_n318), .C2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G902), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n231), .A2(G224), .A3(new_n188), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT7), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n231), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT90), .B(KEYINPUT8), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n234), .B(new_n328), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n249), .A2(new_n297), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT5), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n286), .B1(new_n331), .B2(new_n287), .ZN(new_n332));
  AND3_X1   g146(.A1(new_n330), .A2(new_n332), .A3(new_n279), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n330), .B1(new_n279), .B2(new_n288), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n329), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n198), .A2(KEYINPUT64), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n208), .B1(KEYINPUT0), .B2(G128), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n336), .B1(new_n198), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n225), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n227), .B1(new_n339), .B2(new_n200), .ZN(new_n340));
  AOI22_X1  g154(.A1(new_n340), .A2(new_n229), .B1(new_n226), .B2(new_n227), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n341), .A2(KEYINPUT7), .A3(new_n232), .A4(new_n216), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n325), .A2(new_n327), .A3(new_n335), .A4(new_n342), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n343), .A2(KEYINPUT91), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n314), .B1(new_n343), .B2(KEYINPUT91), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n324), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n196), .B1(new_n323), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n318), .A2(new_n322), .ZN(new_n348));
  INV_X1    g162(.A(new_n233), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n305), .A2(new_n307), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n346), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(new_n352), .A3(new_n195), .ZN(new_n353));
  AOI211_X1 g167(.A(new_n192), .B(new_n194), .C1(new_n347), .C2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT9), .B(G234), .ZN(new_n355));
  OAI21_X1  g169(.A(G221), .B1(new_n355), .B2(G902), .ZN(new_n356));
  XOR2_X1   g170(.A(new_n356), .B(KEYINPUT77), .Z(new_n357));
  INV_X1    g171(.A(G131), .ZN(new_n358));
  INV_X1    g172(.A(G237), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n359), .A2(new_n188), .A3(G214), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n201), .ZN(new_n361));
  NOR2_X1   g175(.A1(G237), .A2(G953), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(G143), .A3(G214), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n358), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT92), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n364), .B(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT96), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT17), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n361), .A2(new_n358), .A3(new_n363), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n366), .A2(new_n367), .A3(new_n368), .A4(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G140), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G125), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n227), .A2(G140), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n373), .A3(KEYINPUT16), .ZN(new_n374));
  OR3_X1    g188(.A1(new_n227), .A2(KEYINPUT16), .A3(G140), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n204), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n374), .A2(new_n375), .A3(G146), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n363), .ZN(new_n380));
  AOI21_X1  g194(.A(G143), .B1(new_n362), .B2(G214), .ZN(new_n381));
  OAI21_X1  g195(.A(G131), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n365), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n361), .A2(new_n363), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(KEYINPUT92), .A3(G131), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n379), .B1(new_n386), .B2(KEYINPUT17), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n383), .A2(new_n368), .A3(new_n385), .A4(new_n369), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(KEYINPUT96), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n370), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(G113), .B(G122), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n391), .B(new_n238), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n384), .A2(KEYINPUT18), .A3(G131), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n372), .A2(new_n373), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G146), .ZN(new_n395));
  XNOR2_X1  g209(.A(G125), .B(G140), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n204), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(KEYINPUT18), .A2(G131), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n361), .A2(new_n363), .A3(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n393), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n390), .A2(new_n392), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n401), .ZN(new_n403));
  OAI211_X1 g217(.A(KEYINPUT93), .B(KEYINPUT19), .C1(new_n394), .C2(KEYINPUT94), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT93), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT94), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n405), .B1(new_n396), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT19), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n408), .B1(new_n396), .B2(new_n405), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n404), .B(new_n204), .C1(new_n407), .C2(new_n409), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n410), .A2(new_n378), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n383), .A2(new_n385), .A3(new_n369), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n403), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT95), .ZN(new_n414));
  NOR3_X1   g228(.A1(new_n413), .A2(new_n414), .A3(new_n392), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(new_n378), .A3(new_n410), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n401), .ZN(new_n417));
  INV_X1    g231(.A(new_n392), .ZN(new_n418));
  AOI21_X1  g232(.A(KEYINPUT95), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n402), .B1(new_n415), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(G475), .A2(G902), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT97), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n414), .B1(new_n413), .B2(new_n392), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n417), .A2(KEYINPUT95), .A3(new_n418), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n423), .B1(new_n426), .B2(new_n402), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n422), .B1(new_n427), .B2(KEYINPUT20), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT20), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n420), .A2(new_n423), .A3(new_n429), .A4(new_n421), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n402), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n390), .A2(new_n401), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n418), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(KEYINPUT98), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT98), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n433), .A2(new_n436), .A3(new_n418), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n432), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(G475), .B1(new_n438), .B2(G902), .ZN(new_n439));
  XNOR2_X1  g253(.A(G128), .B(G143), .ZN(new_n440));
  INV_X1    g254(.A(G134), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n440), .B(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(G116), .B(G122), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n235), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n276), .A2(KEYINPUT14), .A3(G122), .ZN(new_n445));
  XOR2_X1   g259(.A(G116), .B(G122), .Z(new_n446));
  OAI211_X1 g260(.A(G107), .B(new_n445), .C1(new_n446), .C2(KEYINPUT14), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n442), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(G107), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n444), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n440), .A2(new_n441), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(KEYINPUT99), .B(KEYINPUT13), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n201), .A2(G128), .ZN(new_n454));
  OAI21_X1  g268(.A(G134), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n455), .B1(new_n440), .B2(new_n453), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n448), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G217), .ZN(new_n458));
  NOR3_X1   g272(.A1(new_n355), .A2(new_n458), .A3(G953), .ZN(new_n459));
  XOR2_X1   g273(.A(new_n457), .B(new_n459), .Z(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n324), .ZN(new_n461));
  INV_X1    g275(.A(G478), .ZN(new_n462));
  OR2_X1    g276(.A1(new_n462), .A2(KEYINPUT15), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n461), .B(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n431), .A2(new_n439), .A3(new_n464), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n199), .A2(new_n218), .A3(new_n206), .ZN(new_n466));
  AOI211_X1 g280(.A(KEYINPUT69), .B(new_n466), .C1(new_n338), .C2(new_n225), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT69), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n468), .B1(new_n339), .B2(new_n200), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(KEYINPUT80), .B1(new_n254), .B2(new_n249), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n254), .A2(KEYINPUT80), .A3(new_n249), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n470), .B(new_n281), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT11), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n474), .B1(new_n441), .B2(G137), .ZN(new_n475));
  INV_X1    g289(.A(G137), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n476), .A2(KEYINPUT11), .A3(G134), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n441), .A2(G137), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n475), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n479), .B(new_n358), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT10), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n226), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n219), .A2(KEYINPUT66), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n221), .B1(new_n197), .B2(new_n217), .ZN(new_n484));
  OAI22_X1  g298(.A1(new_n483), .A2(new_n484), .B1(new_n197), .B2(new_n223), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n330), .A2(new_n485), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n300), .A2(new_n482), .B1(new_n486), .B2(new_n481), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n473), .A2(new_n480), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT83), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n473), .A2(new_n487), .A3(KEYINPUT83), .A4(new_n480), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n480), .B1(new_n473), .B2(new_n487), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(G110), .B(G140), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n496), .B(KEYINPUT78), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n188), .A2(G227), .ZN(new_n498));
  XOR2_X1   g312(.A(new_n497), .B(new_n498), .Z(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n495), .A2(KEYINPUT84), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT84), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n493), .B1(new_n490), .B2(new_n491), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n502), .B1(new_n503), .B2(new_n499), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n500), .B1(new_n490), .B2(new_n491), .ZN(new_n505));
  OAI22_X1  g319(.A1(new_n483), .A2(new_n484), .B1(new_n207), .B2(new_n223), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n486), .B1(new_n506), .B2(new_n330), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n479), .B(G131), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XOR2_X1   g323(.A(new_n509), .B(KEYINPUT12), .Z(new_n510));
  NAND2_X1  g324(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n501), .A2(new_n504), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(G469), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(new_n513), .A3(new_n324), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n492), .A2(new_n510), .ZN(new_n515));
  AOI22_X1  g329(.A1(new_n515), .A2(new_n500), .B1(new_n505), .B2(new_n494), .ZN(new_n516));
  OAI21_X1  g330(.A(G469), .B1(new_n516), .B2(G902), .ZN(new_n517));
  AOI211_X1 g331(.A(new_n357), .B(new_n465), .C1(new_n514), .C2(new_n517), .ZN(new_n518));
  AND2_X1   g332(.A1(new_n354), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n378), .A2(new_n397), .ZN(new_n520));
  OAI21_X1  g334(.A(G128), .B1(new_n274), .B2(new_n275), .ZN(new_n521));
  NOR2_X1   g335(.A1(G119), .A2(G128), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n521), .A2(KEYINPUT23), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(G110), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n211), .B1(new_n274), .B2(new_n275), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT23), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n524), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT24), .B(G110), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n521), .A2(new_n523), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n520), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  XNOR2_X1  g347(.A(KEYINPUT22), .B(G137), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n534), .B(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n521), .A2(new_n523), .ZN(new_n537));
  INV_X1    g351(.A(new_n530), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n525), .B1(new_n524), .B2(new_n528), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT72), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n379), .B(new_n539), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n540), .A2(new_n541), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n533), .B(new_n536), .C1(new_n542), .C2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT25), .ZN(new_n546));
  AOI21_X1  g360(.A(G902), .B1(new_n546), .B2(KEYINPUT74), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n524), .A2(new_n528), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n541), .B1(new_n548), .B2(G110), .ZN(new_n549));
  INV_X1    g363(.A(new_n378), .ZN(new_n550));
  AOI21_X1  g364(.A(G146), .B1(new_n374), .B2(new_n375), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n539), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n532), .B1(new_n553), .B2(new_n543), .ZN(new_n554));
  XOR2_X1   g368(.A(new_n536), .B(KEYINPUT73), .Z(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n545), .B(new_n547), .C1(new_n554), .C2(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n546), .A2(KEYINPUT74), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n533), .B1(new_n542), .B2(new_n544), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n555), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n562), .A2(new_n545), .A3(new_n547), .A4(new_n558), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n458), .B1(G234), .B2(new_n324), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT75), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n564), .A2(KEYINPUT75), .A3(new_n565), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n565), .A2(G902), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n562), .A2(new_n545), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT76), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n571), .A2(new_n572), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n570), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n568), .A2(new_n569), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n214), .A2(KEYINPUT69), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n339), .A2(new_n468), .A3(new_n200), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(new_n508), .A3(new_n578), .ZN(new_n579));
  OR2_X1    g393(.A1(new_n479), .A2(G131), .ZN(new_n580));
  INV_X1    g394(.A(new_n478), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n441), .A2(G137), .ZN(new_n582));
  OAI21_X1  g396(.A(G131), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n506), .A2(new_n580), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n272), .A2(new_n280), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n579), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(KEYINPUT28), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT28), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n579), .A2(new_n588), .A3(new_n584), .A4(new_n585), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n580), .A2(new_n583), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n591), .A2(new_n226), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n480), .A2(new_n214), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n594), .A2(new_n585), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n590), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT70), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n362), .A2(G210), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(KEYINPUT27), .ZN(new_n600));
  XNOR2_X1  g414(.A(KEYINPUT26), .B(G101), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n597), .A2(new_n598), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n595), .B1(new_n587), .B2(new_n589), .ZN(new_n605));
  OAI21_X1  g419(.A(KEYINPUT70), .B1(new_n605), .B2(new_n602), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n579), .A2(KEYINPUT30), .A3(new_n584), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT30), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n608), .B1(new_n592), .B2(new_n593), .ZN(new_n609));
  INV_X1    g423(.A(new_n585), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n607), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n611), .A2(new_n586), .A3(new_n602), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(KEYINPUT31), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT31), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n611), .A2(new_n614), .A3(new_n586), .A4(new_n602), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n604), .A2(new_n606), .A3(new_n613), .A4(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(G472), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n616), .A2(new_n617), .A3(new_n324), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(KEYINPUT32), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT32), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n616), .A2(new_n620), .A3(new_n617), .A4(new_n324), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n579), .A2(new_n584), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n610), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n590), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n602), .A2(KEYINPUT29), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n611), .A2(new_n586), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n603), .ZN(new_n628));
  AOI22_X1  g442(.A1(new_n628), .A2(KEYINPUT71), .B1(new_n602), .B2(new_n605), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n605), .A2(KEYINPUT71), .A3(new_n602), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT29), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OAI221_X1 g446(.A(new_n324), .B1(new_n625), .B2(new_n626), .C1(new_n629), .C2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(G472), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n576), .B1(new_n622), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n519), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G101), .ZN(G3));
  NAND2_X1  g451(.A1(new_n514), .A2(new_n517), .ZN(new_n638));
  INV_X1    g452(.A(new_n618), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n617), .B1(new_n616), .B2(new_n324), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n639), .A2(new_n576), .A3(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n357), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n638), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n460), .A2(new_n462), .A3(new_n324), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n462), .A2(new_n324), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n460), .B(KEYINPUT33), .ZN(new_n647));
  OAI211_X1 g461(.A(new_n644), .B(new_n646), .C1(new_n647), .C2(new_n462), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n648), .B1(new_n431), .B2(new_n439), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n643), .A2(new_n354), .A3(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT34), .B(G104), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G6));
  XNOR2_X1  g466(.A(new_n422), .B(KEYINPUT20), .ZN(new_n653));
  INV_X1    g467(.A(new_n464), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n653), .A2(new_n654), .A3(new_n439), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n643), .A2(new_n354), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT35), .B(G107), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G9));
  INV_X1    g472(.A(new_n640), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n618), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n555), .A2(KEYINPUT36), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(new_n561), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n570), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n568), .A2(new_n569), .A3(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT100), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(KEYINPUT75), .B1(new_n564), .B2(new_n565), .ZN(new_n667));
  INV_X1    g481(.A(new_n565), .ZN(new_n668));
  AOI211_X1 g482(.A(new_n567), .B(new_n668), .C1(new_n560), .C2(new_n563), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n670), .A2(KEYINPUT100), .A3(new_n663), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n660), .B1(new_n666), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n519), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT37), .B(G110), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G12));
  AOI22_X1  g489(.A1(new_n622), .A2(new_n634), .B1(new_n666), .B2(new_n671), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n194), .B1(new_n347), .B2(new_n353), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n357), .B1(new_n514), .B2(new_n517), .ZN(new_n678));
  INV_X1    g492(.A(G900), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n190), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n189), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n653), .A2(new_n654), .A3(new_n439), .A4(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n676), .A2(new_n677), .A3(new_n678), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G128), .ZN(G30));
  XNOR2_X1  g500(.A(new_n682), .B(KEYINPUT39), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n678), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n688), .A2(KEYINPUT40), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(KEYINPUT40), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n347), .A2(new_n353), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT38), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n627), .A2(new_n602), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n624), .A2(new_n586), .A3(new_n603), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n693), .A2(new_n324), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(G472), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n622), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(KEYINPUT100), .B1(new_n670), .B2(new_n663), .ZN(new_n698));
  INV_X1    g512(.A(new_n663), .ZN(new_n699));
  NOR4_X1   g513(.A1(new_n667), .A2(new_n669), .A3(new_n665), .A4(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n464), .B1(new_n431), .B2(new_n439), .ZN(new_n702));
  AND4_X1   g516(.A1(new_n193), .A2(new_n697), .A3(new_n701), .A4(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n689), .A2(new_n690), .A3(new_n692), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT101), .B(G143), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G45));
  INV_X1    g520(.A(new_n682), .ZN(new_n707));
  AOI211_X1 g521(.A(new_n707), .B(new_n648), .C1(new_n431), .C2(new_n439), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n676), .A2(new_n677), .A3(new_n678), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G146), .ZN(G48));
  AND3_X1   g524(.A1(new_n512), .A2(new_n513), .A3(new_n324), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n513), .B1(new_n512), .B2(new_n324), .ZN(new_n712));
  INV_X1    g526(.A(new_n356), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n354), .A2(new_n635), .A3(new_n649), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(KEYINPUT41), .B(G113), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G15));
  NAND4_X1  g531(.A1(new_n354), .A2(new_n635), .A3(new_n655), .A4(new_n714), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G116), .ZN(G18));
  NOR2_X1   g533(.A1(new_n465), .A2(new_n192), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n714), .A2(new_n676), .A3(new_n720), .A4(new_n677), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G119), .ZN(G21));
  INV_X1    g536(.A(KEYINPUT103), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n431), .A2(new_n439), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n723), .B1(new_n724), .B2(new_n654), .ZN(new_n725));
  AOI211_X1 g539(.A(KEYINPUT103), .B(new_n464), .C1(new_n431), .C2(new_n439), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n617), .A2(new_n324), .ZN(new_n728));
  AND2_X1   g542(.A1(new_n613), .A2(new_n615), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n625), .A2(new_n603), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n616), .A2(new_n324), .ZN(new_n732));
  XOR2_X1   g546(.A(KEYINPUT102), .B(G472), .Z(new_n733));
  AOI21_X1  g547(.A(new_n731), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(new_n576), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n736), .A2(new_n192), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n714), .A2(new_n727), .A3(new_n677), .A4(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G122), .ZN(G24));
  NAND2_X1  g553(.A1(new_n512), .A2(new_n324), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(G469), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n741), .A2(new_n356), .A3(new_n514), .ZN(new_n742));
  AOI22_X1  g556(.A1(new_n318), .A2(new_n322), .B1(new_n305), .B2(new_n307), .ZN(new_n743));
  AOI211_X1 g557(.A(new_n196), .B(new_n346), .C1(new_n743), .C2(new_n349), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n195), .B1(new_n351), .B2(new_n352), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n193), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n708), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n742), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n734), .B1(new_n698), .B2(new_n700), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(KEYINPUT104), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT104), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n751), .B(new_n734), .C1(new_n698), .C2(new_n700), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n748), .A2(new_n753), .ZN(new_n754));
  XOR2_X1   g568(.A(KEYINPUT105), .B(G125), .Z(new_n755));
  XNOR2_X1  g569(.A(new_n754), .B(new_n755), .ZN(G27));
  NAND3_X1  g570(.A1(new_n347), .A2(new_n193), .A3(new_n353), .ZN(new_n757));
  AOI22_X1  g571(.A1(new_n619), .A2(new_n621), .B1(new_n633), .B2(G472), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n757), .A2(new_n758), .A3(new_n576), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT42), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(KEYINPUT106), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n638), .A2(new_n708), .A3(new_n356), .A4(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n760), .A2(KEYINPUT106), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n759), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n744), .A2(new_n745), .A3(new_n194), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n635), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n764), .B1(new_n768), .B2(new_n762), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(new_n358), .ZN(G33));
  AOI21_X1  g585(.A(new_n713), .B1(new_n514), .B2(new_n517), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n759), .A2(new_n684), .A3(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(new_n441), .ZN(G36));
  NAND2_X1  g588(.A1(new_n515), .A2(new_n500), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n505), .A2(new_n494), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT45), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n516), .A2(KEYINPUT45), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n779), .A2(G469), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(G469), .A2(G902), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n781), .A2(KEYINPUT46), .A3(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT107), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n783), .B(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT46), .B1(new_n781), .B2(new_n782), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(new_n711), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n713), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n788), .A2(new_n687), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n644), .A2(new_n646), .ZN(new_n790));
  INV_X1    g604(.A(new_n647), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n790), .B1(new_n791), .B2(G478), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n431), .A2(new_n792), .A3(new_n439), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n793), .A2(KEYINPUT108), .A3(KEYINPUT43), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT43), .B1(new_n793), .B2(KEYINPUT108), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n796), .A2(KEYINPUT109), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(KEYINPUT109), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n666), .A2(new_n671), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n799), .A2(new_n660), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n797), .A2(new_n798), .A3(KEYINPUT44), .A4(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n797), .A2(new_n798), .A3(new_n800), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT44), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n789), .A2(new_n767), .A3(new_n801), .A4(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G137), .ZN(G39));
  INV_X1    g620(.A(new_n758), .ZN(new_n807));
  NOR4_X1   g621(.A1(new_n757), .A2(new_n807), .A3(new_n747), .A4(new_n735), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n788), .A2(KEYINPUT47), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n788), .A2(KEYINPUT47), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n808), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G140), .ZN(G42));
  NAND2_X1  g626(.A1(new_n741), .A2(new_n514), .ZN(new_n813));
  XOR2_X1   g627(.A(new_n813), .B(KEYINPUT49), .Z(new_n814));
  INV_X1    g628(.A(new_n692), .ZN(new_n815));
  INV_X1    g629(.A(new_n697), .ZN(new_n816));
  NOR4_X1   g630(.A1(new_n793), .A2(new_n576), .A3(new_n194), .A4(new_n357), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n814), .A2(new_n815), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT51), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n742), .A2(new_n757), .ZN(new_n820));
  AND4_X1   g634(.A1(new_n735), .A2(new_n820), .A3(new_n189), .A4(new_n816), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n821), .A2(new_n439), .A3(new_n431), .A4(new_n648), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n794), .A2(new_n795), .A3(new_n681), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n753), .A2(new_n823), .A3(new_n820), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT115), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n826), .B1(new_n742), .B2(new_n193), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n714), .A2(KEYINPUT115), .A3(new_n194), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n815), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(KEYINPUT116), .ZN(new_n830));
  NOR4_X1   g644(.A1(new_n794), .A2(new_n795), .A3(new_n736), .A4(new_n681), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n815), .A2(new_n827), .A3(new_n828), .A4(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n830), .A2(new_n831), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT50), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n830), .A2(KEYINPUT50), .A3(new_n831), .A4(new_n833), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n825), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n642), .B1(new_n813), .B2(KEYINPUT113), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n839), .B1(KEYINPUT113), .B2(new_n813), .ZN(new_n840));
  XOR2_X1   g654(.A(new_n840), .B(KEYINPUT114), .Z(new_n841));
  NOR3_X1   g655(.A1(new_n841), .A2(new_n810), .A3(new_n809), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n831), .A2(new_n767), .ZN(new_n843));
  OAI22_X1  g657(.A1(new_n838), .A2(KEYINPUT117), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n838), .A2(KEYINPUT117), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n819), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT52), .ZN(new_n848));
  INV_X1    g662(.A(new_n752), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n751), .B1(new_n799), .B2(new_n734), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n714), .A2(new_n677), .A3(new_n708), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n685), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n670), .A2(new_n663), .A3(new_n682), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n854), .B1(new_n622), .B2(new_n696), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n727), .A2(new_n855), .A3(new_n677), .A4(new_n772), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n709), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n848), .B1(new_n853), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n638), .A2(new_n642), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n859), .A2(new_n746), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n701), .A2(new_n758), .A3(new_n683), .ZN(new_n861));
  AOI22_X1  g675(.A1(new_n748), .A2(new_n753), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n856), .A2(new_n709), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n862), .A2(new_n863), .A3(KEYINPUT52), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n858), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT53), .B1(new_n865), .B2(KEYINPUT110), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n638), .A2(new_n356), .A3(new_n708), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n867), .B1(new_n849), .B2(new_n850), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n653), .A2(new_n464), .A3(new_n439), .A4(new_n682), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n701), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n870), .A2(new_n807), .A3(new_n678), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n757), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n354), .B(new_n518), .C1(new_n635), .C2(new_n672), .ZN(new_n873));
  INV_X1    g687(.A(new_n649), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n874), .B1(new_n464), .B2(new_n724), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n643), .A2(new_n354), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n872), .A2(new_n877), .A3(new_n773), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n715), .A2(new_n718), .A3(new_n721), .A4(new_n738), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n879), .A2(new_n770), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT52), .B1(new_n862), .B2(new_n863), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n853), .A2(new_n848), .A3(new_n857), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n878), .B(new_n880), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  OR2_X1    g697(.A1(new_n866), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n866), .A2(new_n883), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n847), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n765), .B1(new_n759), .B2(new_n763), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n768), .A2(new_n764), .A3(new_n762), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT112), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n715), .A2(new_n738), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n718), .A2(new_n721), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n889), .A2(new_n890), .A3(new_n891), .A4(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT112), .B1(new_n879), .B2(new_n770), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT53), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n896), .B1(new_n858), .B2(new_n864), .ZN(new_n897));
  INV_X1    g711(.A(new_n877), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n772), .A2(new_n708), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n750), .B2(new_n752), .ZN(new_n900));
  NOR4_X1   g714(.A1(new_n859), .A2(new_n701), .A3(new_n758), .A4(new_n869), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n767), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n773), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n898), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(KEYINPUT111), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT111), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n898), .A2(new_n902), .A3(new_n903), .A4(new_n906), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n895), .A2(new_n897), .A3(new_n905), .A4(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n883), .A2(new_n896), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n908), .A2(new_n909), .A3(new_n847), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n886), .A2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(G952), .ZN(new_n912));
  AOI211_X1 g726(.A(new_n912), .B(G953), .C1(new_n821), .C2(new_n649), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n823), .A2(new_n820), .A3(new_n635), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n915), .A2(KEYINPUT119), .A3(KEYINPUT48), .ZN(new_n916));
  XOR2_X1   g730(.A(KEYINPUT119), .B(KEYINPUT48), .Z(new_n917));
  NAND2_X1  g731(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n831), .A2(new_n677), .A3(new_n714), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n913), .A2(new_n916), .A3(new_n918), .A4(new_n919), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n825), .A2(KEYINPUT118), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n825), .A2(KEYINPUT118), .ZN(new_n922));
  OAI21_X1  g736(.A(KEYINPUT51), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n809), .A2(new_n810), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n843), .B1(new_n924), .B2(new_n840), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n836), .A2(new_n837), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n920), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n846), .A2(new_n911), .A3(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(G952), .A2(G953), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n818), .B1(new_n929), .B2(new_n930), .ZN(G75));
  NOR2_X1   g745(.A1(new_n188), .A2(G952), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n324), .B1(new_n908), .B2(new_n909), .ZN(new_n934));
  AOI211_X1 g748(.A(KEYINPUT120), .B(KEYINPUT56), .C1(new_n934), .C2(G210), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n743), .A2(new_n349), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n936), .A2(new_n323), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT55), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n933), .B1(new_n935), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n939), .B1(new_n938), .B2(new_n935), .ZN(G51));
  AOI211_X1 g754(.A(new_n324), .B(new_n781), .C1(new_n908), .C2(new_n909), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n782), .B(KEYINPUT57), .Z(new_n942));
  AOI21_X1  g756(.A(new_n847), .B1(new_n908), .B2(new_n909), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n942), .B1(new_n910), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n941), .B1(new_n944), .B2(new_n512), .ZN(new_n945));
  OAI21_X1  g759(.A(KEYINPUT121), .B1(new_n945), .B2(new_n932), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT121), .ZN(new_n947));
  INV_X1    g761(.A(new_n512), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n908), .A2(new_n909), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(KEYINPUT54), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n908), .A2(new_n909), .A3(new_n847), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n948), .B1(new_n952), .B2(new_n942), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n947), .B(new_n933), .C1(new_n953), .C2(new_n941), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n946), .A2(new_n954), .ZN(G54));
  AND2_X1   g769(.A1(KEYINPUT58), .A2(G475), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n934), .A2(new_n420), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n420), .B1(new_n934), .B2(new_n956), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n957), .A2(new_n958), .A3(new_n932), .ZN(G60));
  XNOR2_X1  g773(.A(new_n645), .B(KEYINPUT59), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n961), .B1(new_n886), .B2(new_n910), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n932), .B1(new_n962), .B2(new_n791), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n791), .A2(new_n960), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n964), .B1(new_n910), .B2(new_n943), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT122), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n952), .A2(KEYINPUT122), .A3(new_n964), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n963), .A2(new_n969), .ZN(G63));
  NAND2_X1  g784(.A1(G217), .A2(G902), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT60), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n972), .B1(new_n908), .B2(new_n909), .ZN(new_n973));
  OR2_X1    g787(.A1(new_n573), .A2(new_n574), .ZN(new_n974));
  OR2_X1    g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n932), .B1(new_n973), .B2(new_n662), .ZN(new_n976));
  AOI21_X1  g790(.A(KEYINPUT123), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT61), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n977), .B(new_n978), .ZN(G66));
  INV_X1    g793(.A(G224), .ZN(new_n980));
  OAI21_X1  g794(.A(G953), .B1(new_n191), .B2(new_n980), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n879), .A2(new_n877), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n981), .B1(new_n982), .B2(G953), .ZN(new_n983));
  INV_X1    g797(.A(G898), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n743), .B1(new_n984), .B2(G953), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n983), .B(new_n985), .Z(G69));
  NAND2_X1  g800(.A1(new_n607), .A2(new_n609), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n404), .B1(new_n407), .B2(new_n409), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(G900), .A2(G953), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n811), .A2(new_n805), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n862), .A2(new_n709), .ZN(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n770), .A2(new_n773), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n789), .A2(new_n635), .A3(new_n677), .A4(new_n727), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n991), .A2(new_n993), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n989), .B(new_n990), .C1(new_n996), .C2(G953), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n875), .B(KEYINPUT124), .ZN(new_n998));
  AND4_X1   g812(.A1(new_n678), .A2(new_n998), .A3(new_n687), .A4(new_n759), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n993), .A2(KEYINPUT62), .A3(new_n704), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT62), .ZN(new_n1001));
  INV_X1    g815(.A(new_n704), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1001), .B1(new_n1002), .B2(new_n992), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n999), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(G953), .B1(new_n991), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n997), .B1(new_n1005), .B2(new_n989), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1007), .ZN(new_n1009));
  OAI211_X1 g823(.A(new_n997), .B(new_n1009), .C1(new_n1005), .C2(new_n989), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1008), .A2(new_n1010), .ZN(G72));
  XOR2_X1   g825(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n1012));
  NOR2_X1   g826(.A1(new_n617), .A2(new_n324), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n1014), .B(KEYINPUT126), .ZN(new_n1015));
  INV_X1    g829(.A(new_n982), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1015), .B1(new_n996), .B2(new_n1016), .ZN(new_n1017));
  AND2_X1   g831(.A1(new_n586), .A2(new_n603), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1017), .A2(new_n611), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n884), .A2(new_n885), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1014), .B1(new_n628), .B2(new_n612), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n932), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n991), .A2(new_n982), .A3(new_n1004), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n693), .B1(new_n1024), .B2(new_n1015), .ZN(new_n1025));
  OR2_X1    g839(.A1(new_n1025), .A2(KEYINPUT127), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1025), .A2(KEYINPUT127), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1023), .B1(new_n1026), .B2(new_n1027), .ZN(G57));
endmodule


