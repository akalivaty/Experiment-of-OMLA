//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 1 1 0 0 0 0 1 0 0 0 0 0 0 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:59 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n558,
    new_n560, new_n561, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n576, new_n577, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n616, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT66), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  XNOR2_X1  g034(.A(KEYINPUT67), .B(G2105), .ZN(new_n460));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  AND2_X1   g036(.A1(new_n461), .A2(G125), .ZN(new_n462));
  AND2_X1   g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n465), .A2(G101), .A3(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(new_n460), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G137), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n464), .A2(new_n466), .A3(new_n473), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n474), .B(KEYINPUT68), .ZN(G160));
  NAND2_X1  g050(.A1(new_n465), .A2(KEYINPUT67), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n471), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OAI221_X1 g056(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n479), .C2(G112), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n471), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n479), .A2(new_n461), .ZN(new_n488));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n468), .A2(new_n470), .A3(G126), .ZN(new_n491));
  NAND2_X1  g066(.A1(G114), .A2(G2104), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n465), .A2(G102), .A3(G2104), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n487), .A2(new_n489), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n479), .A2(new_n461), .A3(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n490), .A2(new_n494), .A3(new_n495), .A4(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT6), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT69), .B1(new_n501), .B2(G651), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n503), .A2(new_n504), .A3(KEYINPUT6), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n501), .A2(G651), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n506), .A2(G543), .A3(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G50), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n500), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n502), .A2(new_n505), .B1(new_n501), .B2(G651), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n511), .A2(KEYINPUT70), .A3(G50), .A4(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  AND2_X1   g093(.A1(new_n511), .A2(new_n518), .ZN(new_n519));
  XOR2_X1   g094(.A(KEYINPUT71), .B(G88), .Z(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(G75), .A2(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n515), .A2(new_n517), .ZN(new_n523));
  INV_X1    g098(.A(G62), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n513), .A2(new_n521), .A3(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  INV_X1    g105(.A(G89), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n511), .A2(new_n518), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n518), .A2(G63), .A3(G651), .ZN(new_n533));
  INV_X1    g108(.A(G51), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n508), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT72), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n535), .A2(new_n536), .ZN(new_n538));
  OAI221_X1 g113(.A(new_n530), .B1(new_n531), .B2(new_n532), .C1(new_n537), .C2(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  NAND2_X1  g115(.A1(new_n519), .A2(G90), .ZN(new_n541));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G64), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n523), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G651), .ZN(new_n545));
  INV_X1    g120(.A(new_n508), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G52), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n541), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(G171));
  NAND2_X1  g124(.A1(new_n519), .A2(G81), .ZN(new_n550));
  NAND2_X1  g125(.A1(G68), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G56), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n523), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G651), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n546), .A2(G43), .ZN(new_n555));
  AND3_X1   g130(.A1(new_n550), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(new_n518), .A2(KEYINPUT74), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT74), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n523), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g140(.A(KEYINPUT75), .B(G65), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n563), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n504), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AND2_X1   g144(.A1(new_n519), .A2(G91), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n511), .A2(G53), .A3(G543), .ZN(new_n572));
  AND2_X1   g147(.A1(KEYINPUT73), .A2(KEYINPUT9), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n572), .B(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n571), .A2(new_n574), .ZN(G299));
  INV_X1    g150(.A(KEYINPUT76), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n548), .B(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(G301));
  OAI21_X1  g153(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n579));
  INV_X1    g154(.A(G49), .ZN(new_n580));
  INV_X1    g155(.A(G87), .ZN(new_n581));
  OAI221_X1 g156(.A(new_n579), .B1(new_n508), .B2(new_n580), .C1(new_n532), .C2(new_n581), .ZN(G288));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n523), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(G651), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n511), .A2(G86), .A3(new_n518), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n511), .A2(G48), .A3(G543), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G305));
  AOI22_X1  g164(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n590), .A2(new_n504), .ZN(new_n591));
  XOR2_X1   g166(.A(new_n591), .B(KEYINPUT77), .Z(new_n592));
  XNOR2_X1  g167(.A(KEYINPUT78), .B(G47), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n546), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(G85), .ZN(new_n595));
  OAI211_X1 g170(.A(new_n592), .B(new_n594), .C1(new_n595), .C2(new_n532), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n563), .A2(G66), .A3(new_n565), .ZN(new_n598));
  INV_X1    g173(.A(G79), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(new_n514), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT79), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n600), .A2(new_n601), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n602), .A2(G651), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n546), .A2(G54), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n519), .A2(G92), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT10), .Z(new_n607));
  NAND3_X1  g182(.A1(new_n604), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n597), .B1(new_n609), .B2(G868), .ZN(G321));
  XNOR2_X1  g185(.A(G321), .B(KEYINPUT80), .ZN(G284));
  NAND2_X1  g186(.A1(G286), .A2(G868), .ZN(new_n612));
  INV_X1    g187(.A(G299), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(G868), .B2(new_n613), .ZN(G297));
  OAI21_X1  g189(.A(new_n612), .B1(G868), .B2(new_n613), .ZN(G280));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n609), .B1(new_n616), .B2(G860), .ZN(G148));
  NAND2_X1  g192(.A1(new_n609), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G868), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(G868), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g196(.A1(new_n465), .A2(G2104), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n471), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(KEYINPUT81), .B(KEYINPUT12), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(G2100), .Z(new_n627));
  NAND2_X1  g202(.A1(new_n480), .A2(G123), .ZN(new_n628));
  OAI221_X1 g203(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n479), .C2(G111), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n483), .A2(G135), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(G2096), .Z(new_n632));
  NAND2_X1  g207(.A1(new_n627), .A2(new_n632), .ZN(G156));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2438), .ZN(new_n635));
  XOR2_X1   g210(.A(G2427), .B(G2430), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(KEYINPUT83), .B(KEYINPUT14), .Z(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(KEYINPUT82), .B(KEYINPUT16), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2451), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2454), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n639), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n645), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(new_n649), .A3(G14), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(G401));
  XNOR2_X1  g226(.A(G2072), .B(G2078), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(KEYINPUT86), .ZN(new_n654));
  XOR2_X1   g229(.A(G2067), .B(G2678), .Z(new_n655));
  INV_X1    g230(.A(KEYINPUT86), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n654), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2084), .B(G2090), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT87), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n652), .B(KEYINPUT17), .Z(new_n662));
  OAI21_X1  g237(.A(new_n661), .B1(new_n655), .B2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n659), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n662), .A2(new_n655), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(KEYINPUT84), .B(KEYINPUT18), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT85), .ZN(new_n667));
  NOR3_X1   g242(.A1(new_n653), .A2(new_n655), .A3(new_n659), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n663), .A2(new_n665), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2096), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2100), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(G227));
  XNOR2_X1  g248(.A(KEYINPUT90), .B(G1986), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1971), .B(G1976), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT88), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  AND2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT89), .B(KEYINPUT20), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n679), .A2(new_n680), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n678), .A2(new_n685), .ZN(new_n686));
  OR3_X1    g261(.A1(new_n678), .A2(new_n681), .A3(new_n685), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n684), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n689));
  OR2_X1    g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1991), .B(G1996), .ZN(new_n691));
  INV_X1    g266(.A(G1981), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n688), .A2(new_n689), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n690), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n694), .B1(new_n690), .B2(new_n695), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n675), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n698), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n700), .A2(new_n674), .A3(new_n696), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n699), .A2(new_n701), .ZN(G229));
  XOR2_X1   g277(.A(KEYINPUT92), .B(KEYINPUT36), .Z(new_n703));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G24), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(G290), .B2(G16), .ZN(new_n707));
  INV_X1    g282(.A(G1986), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n480), .ZN(new_n710));
  INV_X1    g285(.A(G119), .ZN(new_n711));
  OR3_X1    g286(.A1(new_n710), .A2(KEYINPUT91), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(KEYINPUT91), .B1(new_n710), .B2(new_n711), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n483), .A2(G131), .ZN(new_n714));
  OAI221_X1 g289(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n479), .C2(G107), .ZN(new_n715));
  NAND4_X1  g290(.A1(new_n712), .A2(new_n713), .A3(new_n714), .A4(new_n715), .ZN(new_n716));
  MUX2_X1   g291(.A(G25), .B(new_n716), .S(G29), .Z(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT35), .B(G1991), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n717), .B(new_n718), .Z(new_n719));
  NAND2_X1  g294(.A1(new_n707), .A2(new_n708), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n709), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G288), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G16), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G16), .B2(G23), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT33), .B(G1976), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n586), .A2(new_n588), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n728), .A2(G16), .A3(new_n587), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT32), .ZN(new_n730));
  OR2_X1    g305(.A1(G6), .A2(G16), .ZN(new_n731));
  AND3_X1   g306(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n730), .B1(new_n729), .B2(new_n731), .ZN(new_n733));
  OR3_X1    g308(.A1(new_n732), .A2(new_n733), .A3(new_n692), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n692), .B1(new_n732), .B2(new_n733), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n704), .A2(G22), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G166), .B2(new_n704), .ZN(new_n738));
  INV_X1    g313(.A(G1971), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n727), .A2(new_n736), .A3(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT34), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n727), .A2(new_n736), .A3(KEYINPUT34), .A4(new_n740), .ZN(new_n744));
  AOI211_X1 g319(.A(new_n703), .B(new_n721), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n746), .A2(KEYINPUT93), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n721), .B1(new_n743), .B2(new_n744), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT36), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT93), .ZN(new_n751));
  NOR3_X1   g326(.A1(new_n750), .A2(new_n745), .A3(new_n751), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n704), .A2(KEYINPUT23), .A3(G20), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT23), .ZN(new_n754));
  INV_X1    g329(.A(G20), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n754), .B1(new_n755), .B2(G16), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n753), .B(new_n756), .C1(new_n613), .C2(new_n704), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT103), .B(G1956), .Z(new_n758));
  NOR2_X1   g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT28), .ZN(new_n760));
  INV_X1    g335(.A(G26), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n760), .B1(new_n761), .B2(G29), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n761), .A2(G29), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n480), .A2(G128), .ZN(new_n764));
  OAI221_X1 g339(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n479), .C2(G116), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n483), .A2(G140), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n763), .B1(new_n767), .B2(G29), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n762), .B1(new_n768), .B2(new_n760), .ZN(new_n769));
  NOR2_X1   g344(.A1(G27), .A2(G29), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G164), .B2(G29), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n769), .A2(G2067), .B1(new_n771), .B2(G2078), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT30), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n773), .A2(G28), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(G28), .ZN(new_n775));
  INV_X1    g350(.A(G29), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n772), .B(new_n777), .C1(G2067), .C2(new_n769), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n704), .A2(G5), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G171), .B2(new_n704), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT99), .Z(new_n781));
  INV_X1    g356(.A(G1961), .ZN(new_n782));
  OAI21_X1  g357(.A(KEYINPUT100), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n780), .B(KEYINPUT99), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT100), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n784), .A2(new_n785), .A3(G1961), .ZN(new_n786));
  AOI211_X1 g361(.A(new_n759), .B(new_n778), .C1(new_n783), .C2(new_n786), .ZN(new_n787));
  OR2_X1    g362(.A1(G4), .A2(G16), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n608), .B2(new_n704), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT94), .B(G1348), .Z(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n631), .A2(new_n776), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n704), .A2(G19), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n556), .B2(new_n704), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(G1341), .Z(new_n796));
  NAND4_X1  g371(.A1(new_n787), .A2(new_n792), .A3(new_n793), .A4(new_n796), .ZN(new_n797));
  OR2_X1    g372(.A1(KEYINPUT24), .A2(G34), .ZN(new_n798));
  NAND2_X1  g373(.A1(KEYINPUT24), .A2(G34), .ZN(new_n799));
  AOI21_X1  g374(.A(G29), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G160), .B2(G29), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT101), .ZN(new_n802));
  OR3_X1    g377(.A1(new_n801), .A2(new_n802), .A3(G2084), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n801), .B2(G2084), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n781), .A2(new_n782), .ZN(new_n806));
  INV_X1    g381(.A(G35), .ZN(new_n807));
  OAI21_X1  g382(.A(KEYINPUT102), .B1(new_n807), .B2(G29), .ZN(new_n808));
  OR3_X1    g383(.A1(new_n807), .A2(KEYINPUT102), .A3(G29), .ZN(new_n809));
  OAI211_X1 g384(.A(new_n808), .B(new_n809), .C1(G162), .C2(new_n776), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT29), .B(G2090), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT98), .B(KEYINPUT31), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G11), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n805), .A2(new_n806), .A3(new_n812), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n757), .A2(new_n758), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n801), .A2(G2084), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n816), .B(new_n817), .C1(new_n789), .C2(new_n791), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(G29), .A2(G33), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n483), .A2(G139), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n479), .A2(G103), .A3(G2104), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT25), .Z(new_n823));
  AOI22_X1  g398(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT95), .Z(new_n825));
  OAI211_X1 g400(.A(new_n821), .B(new_n823), .C1(new_n825), .C2(new_n479), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT96), .Z(new_n827));
  AOI21_X1  g402(.A(new_n820), .B1(new_n827), .B2(G29), .ZN(new_n828));
  INV_X1    g403(.A(G2072), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AOI211_X1 g405(.A(G2072), .B(new_n820), .C1(new_n827), .C2(G29), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n776), .A2(G32), .ZN(new_n833));
  AOI22_X1  g408(.A1(G129), .A2(new_n480), .B1(new_n483), .B2(G141), .ZN(new_n834));
  NAND3_X1  g409(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT26), .Z(new_n836));
  INV_X1    g411(.A(G105), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n834), .B(new_n836), .C1(new_n837), .C2(new_n622), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n833), .B1(new_n838), .B2(G29), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT97), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT27), .B(G1996), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n819), .A2(new_n832), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n797), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT104), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n771), .A2(G2078), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n704), .A2(G21), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(G168), .B2(new_n704), .ZN(new_n849));
  INV_X1    g424(.A(G1966), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n845), .A2(new_n846), .A3(new_n847), .A4(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n830), .A2(new_n831), .ZN(new_n853));
  NOR4_X1   g428(.A1(new_n853), .A2(new_n815), .A3(new_n842), .A4(new_n818), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n783), .A2(new_n786), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n759), .A2(new_n778), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n855), .A2(new_n793), .A3(new_n796), .A4(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n792), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n854), .A2(new_n859), .A3(new_n847), .A4(new_n851), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(KEYINPUT104), .ZN(new_n861));
  AOI211_X1 g436(.A(new_n747), .B(new_n752), .C1(new_n852), .C2(new_n861), .ZN(G311));
  NAND2_X1  g437(.A1(new_n852), .A2(new_n861), .ZN(new_n863));
  INV_X1    g438(.A(new_n747), .ZN(new_n864));
  INV_X1    g439(.A(new_n752), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(G150));
  NAND2_X1  g441(.A1(new_n519), .A2(G93), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n546), .A2(G55), .ZN(new_n868));
  AOI22_X1  g443(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n867), .B(new_n868), .C1(new_n504), .C2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(G860), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(KEYINPUT37), .Z(new_n872));
  OAI21_X1  g447(.A(new_n556), .B1(new_n870), .B2(KEYINPUT105), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n870), .A2(KEYINPUT105), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n873), .B(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n609), .A2(G559), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT38), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(KEYINPUT39), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n877), .A2(KEYINPUT39), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n875), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n880), .ZN(new_n882));
  INV_X1    g457(.A(new_n875), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(new_n883), .A3(new_n878), .ZN(new_n884));
  INV_X1    g459(.A(G860), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n881), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT106), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n886), .A2(new_n887), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n872), .B1(new_n888), .B2(new_n889), .ZN(G145));
  XNOR2_X1  g465(.A(G160), .B(new_n631), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(new_n485), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n838), .B(G164), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(new_n767), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT107), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(new_n826), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n827), .ZN(new_n897));
  AOI22_X1  g472(.A1(G130), .A2(new_n480), .B1(new_n483), .B2(G142), .ZN(new_n898));
  OAI221_X1 g473(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n479), .C2(G118), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(new_n625), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(new_n716), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n902), .A2(KEYINPUT108), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n896), .A2(new_n897), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n903), .B1(new_n896), .B2(new_n897), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n892), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n896), .A2(new_n897), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n902), .ZN(new_n908));
  INV_X1    g483(.A(new_n892), .ZN(new_n909));
  INV_X1    g484(.A(new_n902), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n896), .A2(new_n910), .A3(new_n897), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n908), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(G37), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n906), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT40), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT40), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n906), .A2(new_n912), .A3(new_n916), .A4(new_n913), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(G395));
  NOR2_X1   g493(.A1(new_n870), .A2(G868), .ZN(new_n919));
  XNOR2_X1  g494(.A(G288), .B(G305), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(G166), .ZN(new_n921));
  INV_X1    g496(.A(G290), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n921), .B(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(KEYINPUT42), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT109), .ZN(new_n925));
  OR2_X1    g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n925), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n618), .B(new_n875), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n608), .A2(G299), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n613), .A2(new_n604), .A3(new_n605), .A4(new_n607), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n929), .A2(KEYINPUT41), .A3(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT41), .B1(new_n929), .B2(new_n930), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n928), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n929), .A2(new_n930), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n928), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n926), .A2(new_n927), .A3(new_n935), .A4(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n935), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n924), .B(new_n925), .C1(new_n940), .C2(new_n937), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n919), .B1(new_n942), .B2(G868), .ZN(G295));
  AOI21_X1  g518(.A(new_n919), .B1(new_n942), .B2(G868), .ZN(G331));
  INV_X1    g519(.A(new_n933), .ZN(new_n945));
  NAND2_X1  g520(.A1(G286), .A2(G171), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n946), .B1(G286), .B2(new_n577), .ZN(new_n947));
  OR2_X1    g522(.A1(new_n947), .A2(new_n875), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n875), .ZN(new_n949));
  AOI22_X1  g524(.A1(new_n945), .A2(new_n931), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n948), .A2(new_n936), .A3(new_n949), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n923), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n923), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n948), .A2(new_n949), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n954), .B(new_n951), .C1(new_n955), .C2(new_n934), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n953), .A2(new_n913), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n953), .A2(new_n956), .A3(new_n960), .A4(new_n913), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n958), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT44), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n953), .A2(new_n956), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n964), .A2(KEYINPUT110), .A3(new_n960), .A4(new_n913), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n962), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n958), .A2(KEYINPUT44), .A3(new_n961), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(G397));
  INV_X1    g543(.A(G1384), .ZN(new_n969));
  INV_X1    g544(.A(new_n492), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n970), .B1(new_n461), .B2(G126), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n495), .B(new_n497), .C1(new_n971), .C2(new_n465), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT4), .B1(new_n472), .B2(G138), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n969), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(KEYINPUT111), .B(KEYINPUT45), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n464), .A2(new_n473), .A3(G40), .A4(new_n466), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n838), .B(G1996), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n767), .B(G2067), .ZN(new_n980));
  OR2_X1    g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n716), .A2(new_n718), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n716), .A2(new_n718), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n981), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n984), .B1(new_n708), .B2(new_n922), .ZN(new_n985));
  NOR2_X1   g560(.A1(G290), .A2(G1986), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n978), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT45), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n974), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n977), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n989), .B(new_n990), .C1(new_n974), .C2(new_n975), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT53), .ZN(new_n992));
  OR3_X1    g567(.A1(new_n991), .A2(new_n992), .A3(G2078), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n977), .B1(new_n974), .B2(new_n975), .ZN(new_n994));
  INV_X1    g569(.A(G2078), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n498), .A2(KEYINPUT45), .A3(new_n969), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  OAI211_X1 g572(.A(KEYINPUT50), .B(new_n969), .C1(new_n972), .C2(new_n973), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT50), .B1(new_n498), .B2(new_n969), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n990), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  XOR2_X1   g576(.A(KEYINPUT122), .B(G1961), .Z(new_n1002));
  AOI22_X1  g577(.A1(new_n992), .A2(new_n997), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n993), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n577), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT54), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT123), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n994), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n992), .A2(G2078), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n994), .A2(new_n1007), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1008), .A2(new_n996), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n1003), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1005), .B(new_n1006), .C1(new_n577), .C2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT124), .B1(new_n1004), .B2(new_n577), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1012), .A2(G171), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT124), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n993), .A2(new_n1003), .A3(new_n1016), .A4(G301), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n1014), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1013), .B1(new_n1018), .B2(new_n1006), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT114), .ZN(new_n1020));
  XNOR2_X1  g595(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n1021));
  AND3_X1   g596(.A1(G303), .A2(G8), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1024), .B1(G303), .B2(G8), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1020), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(G303), .A2(G8), .A3(new_n1021), .ZN(new_n1027));
  INV_X1    g602(.A(G8), .ZN(new_n1028));
  AOI22_X1  g603(.A1(new_n510), .A2(new_n512), .B1(G651), .B2(new_n525), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1028), .B1(new_n1029), .B2(new_n521), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1027), .B(KEYINPUT114), .C1(new_n1030), .C2(new_n1024), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1026), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n976), .A2(new_n990), .A3(new_n996), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n739), .ZN(new_n1034));
  XOR2_X1   g609(.A(KEYINPUT112), .B(G2090), .Z(new_n1035));
  OAI211_X1 g610(.A(new_n990), .B(new_n1035), .C1(new_n999), .C2(new_n1000), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1028), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1032), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT49), .ZN(new_n1039));
  NAND2_X1  g614(.A1(G305), .A2(G1981), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(G305), .A2(G1981), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1039), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n497), .A2(new_n495), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n465), .B1(new_n491), .B2(new_n492), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(G1384), .B1(new_n1046), .B2(new_n490), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1028), .B1(new_n990), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n728), .A2(new_n692), .A3(new_n587), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1049), .A2(KEYINPUT49), .A3(new_n1040), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1043), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n519), .A2(G87), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n546), .A2(G49), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1052), .A2(new_n1053), .A3(G1976), .A4(new_n579), .ZN(new_n1054));
  INV_X1    g629(.A(G1976), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT52), .B1(G288), .B2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1048), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1054), .B(G8), .C1(new_n974), .C2(new_n977), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT52), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1051), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT50), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n974), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n977), .B1(new_n1064), .B2(new_n998), .ZN(new_n1065));
  AOI22_X1  g640(.A1(new_n1065), .A2(new_n1035), .B1(new_n1033), .B2(new_n739), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1062), .B1(new_n1066), .B2(new_n1028), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n1038), .A2(new_n1061), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G2084), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n850), .A2(new_n991), .B1(new_n1065), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT51), .B1(new_n1070), .B2(G168), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1028), .B1(new_n1070), .B2(G168), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT51), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  OR2_X1    g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1019), .A2(new_n1068), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n990), .A2(new_n1047), .ZN(new_n1078));
  XOR2_X1   g653(.A(KEYINPUT58), .B(G1341), .Z(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n1033), .B2(G1996), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(new_n556), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT119), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT59), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT119), .ZN(new_n1086));
  AOI22_X1  g661(.A1(new_n1084), .A2(new_n1086), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1087));
  INV_X1    g662(.A(G1956), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1001), .A2(new_n1088), .ZN(new_n1089));
  XNOR2_X1  g664(.A(KEYINPUT56), .B(G2072), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n976), .A2(new_n990), .A3(new_n996), .A4(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT116), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n994), .A2(KEYINPUT116), .A3(new_n996), .A4(new_n1090), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1089), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n571), .A2(new_n1096), .A3(new_n574), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1096), .B1(new_n571), .B2(new_n574), .ZN(new_n1098));
  OR2_X1    g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1095), .A2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1101), .A2(new_n1089), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT120), .ZN(new_n1104));
  AOI21_X1  g679(.A(KEYINPUT61), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT61), .ZN(new_n1106));
  AOI211_X1 g681(.A(KEYINPUT120), .B(new_n1106), .C1(new_n1100), .C2(new_n1102), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1087), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT121), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  OAI211_X1 g685(.A(KEYINPUT121), .B(new_n1087), .C1(new_n1105), .C2(new_n1107), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1078), .A2(G2067), .ZN(new_n1112));
  INV_X1    g687(.A(G1348), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1112), .B1(new_n1113), .B2(new_n1001), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT60), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n1115), .B(new_n609), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1116), .B1(KEYINPUT60), .B2(new_n1114), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1110), .A2(new_n1111), .A3(new_n1117), .ZN(new_n1118));
  OR3_X1    g693(.A1(new_n1114), .A2(new_n608), .A3(KEYINPUT117), .ZN(new_n1119));
  OAI21_X1  g694(.A(KEYINPUT117), .B1(new_n1114), .B2(new_n608), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1119), .A2(new_n1120), .A3(new_n1100), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n1102), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1077), .B1(new_n1118), .B2(new_n1122), .ZN(new_n1123));
  OR3_X1    g698(.A1(new_n1073), .A2(new_n1075), .A3(KEYINPUT62), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1005), .ZN(new_n1125));
  OAI21_X1  g700(.A(KEYINPUT62), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1124), .A2(new_n1068), .A3(new_n1125), .A4(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT115), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1068), .A2(KEYINPUT63), .A3(G168), .A4(new_n1072), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1060), .B1(new_n1032), .B2(new_n1037), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1130), .A2(G168), .A3(new_n1072), .A4(new_n1067), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT63), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1129), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1051), .A2(new_n1055), .A3(new_n722), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n1049), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(new_n1048), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1137), .B1(new_n1038), .B2(new_n1060), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1128), .B1(new_n1134), .B2(new_n1139), .ZN(new_n1140));
  AOI211_X1 g715(.A(KEYINPUT115), .B(new_n1138), .C1(new_n1129), .C2(new_n1133), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1127), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n987), .B1(new_n1123), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n978), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1144), .A2(G1996), .ZN(new_n1145));
  XOR2_X1   g720(.A(new_n1145), .B(KEYINPUT46), .Z(new_n1146));
  OAI21_X1  g721(.A(new_n978), .B1(new_n838), .B2(new_n980), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1147), .B(KEYINPUT126), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n1149), .B(KEYINPUT47), .ZN(new_n1150));
  INV_X1    g725(.A(new_n983), .ZN(new_n1151));
  OAI22_X1  g726(.A1(new_n981), .A2(new_n1151), .B1(G2067), .B2(new_n767), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n978), .ZN(new_n1153));
  XOR2_X1   g728(.A(new_n1153), .B(KEYINPUT125), .Z(new_n1154));
  NAND2_X1  g729(.A1(new_n986), .A2(new_n978), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(KEYINPUT48), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1156), .B1(new_n1144), .B2(new_n984), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1150), .A2(new_n1154), .A3(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1143), .A2(new_n1159), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g735(.A1(new_n672), .A2(new_n650), .A3(G319), .ZN(new_n1162));
  INV_X1    g736(.A(KEYINPUT127), .ZN(new_n1163));
  NAND2_X1  g737(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND4_X1  g738(.A1(new_n672), .A2(new_n650), .A3(KEYINPUT127), .A4(G319), .ZN(new_n1165));
  AOI21_X1  g739(.A(G229), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NAND4_X1  g740(.A1(new_n962), .A2(new_n914), .A3(new_n965), .A4(new_n1166), .ZN(G225));
  INV_X1    g741(.A(G225), .ZN(G308));
endmodule


