//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 0 1 0 0 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 1 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n858, new_n859, new_n860, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(G8gat), .ZN(new_n206));
  INV_X1    g005(.A(G57gat), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT96), .B1(new_n207), .B2(G64gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT96), .ZN(new_n209));
  INV_X1    g008(.A(G64gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n209), .A2(new_n210), .A3(G57gat), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n208), .B(new_n211), .C1(G57gat), .C2(new_n210), .ZN(new_n212));
  NAND2_X1  g011(.A1(G71gat), .A2(G78gat), .ZN(new_n213));
  OR2_X1    g012(.A1(G71gat), .A2(G78gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT9), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n212), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT97), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n217), .B(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G57gat), .B(G64gat), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n213), .B(new_n214), .C1(new_n220), .C2(new_n215), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n222), .B(KEYINPUT98), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n206), .B1(new_n223), .B2(KEYINPUT21), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT98), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n222), .B(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT21), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G231gat), .A2(G233gat), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n229), .B(new_n231), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n232), .A2(G127gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(G127gat), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n225), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n234), .A2(new_n233), .A3(new_n225), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n238));
  INV_X1    g037(.A(G155gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(G183gat), .B(G211gat), .ZN(new_n241));
  XOR2_X1   g040(.A(new_n240), .B(new_n241), .Z(new_n242));
  NAND3_X1  g041(.A1(new_n236), .A2(new_n237), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n242), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n233), .A2(new_n225), .A3(new_n234), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n244), .B1(new_n245), .B2(new_n235), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G134gat), .B(G162gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(G232gat), .A2(G233gat), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT41), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  XOR2_X1   g050(.A(new_n248), .B(new_n251), .Z(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT99), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n255), .A2(G85gat), .A3(G92gat), .ZN(new_n256));
  MUX2_X1   g055(.A(KEYINPUT7), .B(new_n254), .S(new_n256), .Z(new_n257));
  AND3_X1   g056(.A1(KEYINPUT100), .A2(G99gat), .A3(G106gat), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT100), .B1(G99gat), .B2(G106gat), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT8), .ZN(new_n260));
  NOR3_X1   g059(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  OR2_X1    g060(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(G99gat), .B(G106gat), .Z(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT101), .ZN(new_n265));
  OR3_X1    g064(.A1(new_n257), .A2(new_n263), .A3(new_n261), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n262), .A2(KEYINPUT101), .A3(new_n263), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(G43gat), .A2(G50gat), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(G43gat), .A2(G50gat), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT15), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(G29gat), .A2(G36gat), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT14), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n276), .B1(KEYINPUT86), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(KEYINPUT86), .B(KEYINPUT14), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n278), .B1(new_n279), .B2(new_n276), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT87), .ZN(new_n281));
  XOR2_X1   g080(.A(KEYINPUT88), .B(G36gat), .Z(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(G29gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n280), .A2(KEYINPUT87), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n275), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n272), .A2(KEYINPUT15), .ZN(new_n287));
  XNOR2_X1  g086(.A(KEYINPUT89), .B(G50gat), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n287), .B1(new_n288), .B2(G43gat), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n289), .A2(new_n283), .A3(new_n280), .A4(new_n274), .ZN(new_n290));
  AND2_X1   g089(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  OAI22_X1  g090(.A1(new_n270), .A2(new_n291), .B1(new_n250), .B2(new_n249), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT103), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT103), .ZN(new_n294));
  OAI221_X1 g093(.A(new_n294), .B1(new_n250), .B2(new_n249), .C1(new_n270), .C2(new_n291), .ZN(new_n295));
  XOR2_X1   g094(.A(G190gat), .B(G218gat), .Z(new_n296));
  XNOR2_X1  g095(.A(new_n296), .B(KEYINPUT104), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  AOI22_X1  g097(.A1(new_n293), .A2(new_n295), .B1(KEYINPUT105), .B2(new_n298), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n298), .A2(KEYINPUT105), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT17), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n291), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n286), .A2(new_n290), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT17), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(new_n270), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n307), .B(KEYINPUT102), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n299), .A2(new_n301), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n301), .B1(new_n299), .B2(new_n308), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n253), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n311), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n313), .A2(new_n252), .A3(new_n309), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(G230gat), .A2(G233gat), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT10), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n264), .A2(new_n221), .A3(new_n219), .A4(new_n266), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n318), .B(new_n319), .C1(new_n223), .C2(new_n269), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n223), .A2(KEYINPUT10), .A3(new_n269), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT106), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n317), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n320), .A2(KEYINPUT106), .A3(new_n321), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n319), .B1(new_n223), .B2(new_n269), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(new_n317), .ZN(new_n328));
  XOR2_X1   g127(.A(G120gat), .B(G148gat), .Z(new_n329));
  XNOR2_X1  g128(.A(new_n329), .B(KEYINPUT107), .ZN(new_n330));
  XNOR2_X1  g129(.A(G176gat), .B(G204gat), .ZN(new_n331));
  XOR2_X1   g130(.A(new_n330), .B(new_n331), .Z(new_n332));
  NAND3_X1  g131(.A1(new_n326), .A2(new_n328), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n317), .B1(new_n320), .B2(new_n321), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(new_n328), .ZN(new_n336));
  INV_X1    g135(.A(new_n332), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n247), .A2(new_n315), .A3(new_n340), .ZN(new_n341));
  XOR2_X1   g140(.A(G15gat), .B(G43gat), .Z(new_n342));
  XNOR2_X1  g141(.A(G71gat), .B(G99gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n342), .B(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G127gat), .B(G134gat), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT66), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n346), .B1(new_n347), .B2(KEYINPUT1), .ZN(new_n348));
  XNOR2_X1  g147(.A(G113gat), .B(G120gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n349), .A2(KEYINPUT1), .ZN(new_n350));
  XOR2_X1   g149(.A(new_n348), .B(new_n350), .Z(new_n351));
  NOR3_X1   g150(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n352), .B(KEYINPUT65), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n354));
  INV_X1    g153(.A(G169gat), .ZN(new_n355));
  INV_X1    g154(.A(G176gat), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n353), .B(new_n354), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(G183gat), .A2(G190gat), .ZN(new_n358));
  XOR2_X1   g157(.A(KEYINPUT27), .B(G183gat), .Z(new_n359));
  INV_X1    g158(.A(KEYINPUT64), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(G183gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT27), .ZN(new_n363));
  AOI21_X1  g162(.A(G190gat), .B1(new_n363), .B2(KEYINPUT64), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT28), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT28), .ZN(new_n366));
  NOR3_X1   g165(.A1(new_n359), .A2(new_n366), .A3(G190gat), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n357), .B(new_n358), .C1(new_n365), .C2(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n358), .A2(KEYINPUT24), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n355), .A2(new_n356), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(G190gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n362), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n373), .A2(KEYINPUT24), .A3(new_n358), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NOR3_X1   g175(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n371), .B(new_n374), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT25), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n368), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT67), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n351), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT67), .B1(new_n368), .B2(new_n380), .ZN(new_n384));
  OR2_X1    g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(G227gat), .ZN(new_n386));
  INV_X1    g185(.A(G233gat), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n383), .A2(new_n384), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n385), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT33), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n345), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT34), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n385), .A2(new_n389), .ZN(new_n394));
  INV_X1    g193(.A(new_n388), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AOI211_X1 g195(.A(KEYINPUT34), .B(new_n388), .C1(new_n385), .C2(new_n389), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n392), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NOR3_X1   g198(.A1(new_n392), .A2(new_n396), .A3(new_n397), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n390), .A2(KEYINPUT32), .ZN(new_n401));
  NOR3_X1   g200(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n401), .ZN(new_n403));
  OR3_X1    g202(.A1(new_n392), .A2(new_n396), .A3(new_n397), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n403), .B1(new_n404), .B2(new_n398), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(G8gat), .B(G36gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(G64gat), .B(G92gat), .ZN(new_n408));
  XOR2_X1   g207(.A(new_n407), .B(new_n408), .Z(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT29), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n381), .A2(new_n411), .B1(G226gat), .B2(G233gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(G226gat), .A2(G233gat), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n413), .B1(new_n368), .B2(new_n380), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(G197gat), .B(G204gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(G211gat), .B(G218gat), .ZN(new_n417));
  INV_X1    g216(.A(G218gat), .ZN(new_n418));
  INV_X1    g217(.A(G211gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT68), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT68), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(G211gat), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n418), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n416), .B(new_n417), .C1(new_n423), .C2(KEYINPUT22), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT22), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT68), .B(G211gat), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n426), .B1(new_n427), .B2(new_n418), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n417), .B1(new_n428), .B2(new_n416), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT69), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n432), .B1(new_n425), .B2(new_n429), .ZN(new_n433));
  INV_X1    g232(.A(new_n417), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n420), .A2(new_n422), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT22), .B1(new_n435), .B2(G218gat), .ZN(new_n436));
  INV_X1    g235(.A(new_n416), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n434), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n438), .A2(KEYINPUT69), .A3(new_n424), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n433), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n440), .B1(new_n412), .B2(new_n414), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n410), .B1(new_n431), .B2(new_n441), .ZN(new_n442));
  OR3_X1    g241(.A1(new_n442), .A2(KEYINPUT70), .A3(KEYINPUT30), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n431), .A2(new_n441), .A3(new_n410), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT30), .B1(new_n442), .B2(KEYINPUT70), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT6), .ZN(new_n447));
  NAND2_X1  g246(.A1(G155gat), .A2(G162gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT2), .ZN(new_n449));
  INV_X1    g248(.A(G148gat), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n450), .A2(G141gat), .ZN(new_n451));
  INV_X1    g250(.A(G141gat), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n452), .A2(G148gat), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n449), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(G162gat), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n239), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT71), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n456), .A2(new_n457), .A3(new_n448), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n457), .B1(new_n456), .B2(new_n448), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n454), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT72), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n461), .B1(new_n450), .B2(G141gat), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT73), .B1(new_n452), .B2(G148gat), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT73), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n464), .A2(new_n450), .A3(G141gat), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n452), .A2(KEYINPUT72), .A3(G148gat), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n462), .A2(new_n463), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n448), .B1(new_n456), .B2(KEYINPUT2), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n460), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n351), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT4), .ZN(new_n472));
  NAND2_X1  g271(.A1(G225gat), .A2(G233gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n470), .A2(KEYINPUT3), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT3), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n460), .A2(new_n469), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n351), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n348), .B(new_n350), .ZN(new_n478));
  AND2_X1   g277(.A1(new_n460), .A2(new_n469), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT4), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n472), .A2(new_n473), .A3(new_n477), .A4(new_n482), .ZN(new_n483));
  OR2_X1    g282(.A1(new_n483), .A2(KEYINPUT5), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n478), .A2(new_n479), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n471), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT74), .B1(new_n486), .B2(new_n473), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT74), .ZN(new_n488));
  INV_X1    g287(.A(new_n473), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n488), .B(new_n489), .C1(new_n471), .C2(new_n485), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n487), .A2(new_n483), .A3(KEYINPUT5), .A4(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n484), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(G1gat), .B(G29gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n493), .B(KEYINPUT0), .ZN(new_n494));
  XNOR2_X1  g293(.A(G57gat), .B(G85gat), .ZN(new_n495));
  XOR2_X1   g294(.A(new_n494), .B(new_n495), .Z(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n447), .B1(new_n492), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n498), .A2(KEYINPUT75), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n492), .A2(new_n497), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n498), .A2(KEYINPUT75), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT76), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n504), .B1(new_n501), .B2(new_n447), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n492), .A2(KEYINPUT76), .A3(KEYINPUT6), .A4(new_n497), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n446), .B1(new_n503), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n476), .A2(new_n411), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n433), .A2(new_n510), .A3(new_n439), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT29), .B1(new_n438), .B2(new_n424), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n470), .B1(new_n512), .B2(KEYINPUT3), .ZN(new_n513));
  INV_X1    g312(.A(G228gat), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n514), .A2(new_n387), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n511), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT79), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n516), .B(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT77), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n513), .A2(new_n519), .B1(new_n430), .B2(new_n510), .ZN(new_n520));
  OAI211_X1 g319(.A(KEYINPUT77), .B(new_n470), .C1(new_n512), .C2(KEYINPUT3), .ZN(new_n521));
  AOI211_X1 g320(.A(KEYINPUT78), .B(new_n515), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT78), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n513), .A2(new_n519), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n510), .A2(new_n430), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(new_n521), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n515), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n523), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n518), .B1(new_n522), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT82), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n529), .A2(new_n530), .A3(G22gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(G78gat), .B(G106gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(KEYINPUT31), .B(G50gat), .ZN(new_n533));
  XOR2_X1   g332(.A(new_n532), .B(new_n533), .Z(new_n534));
  XNOR2_X1  g333(.A(new_n516), .B(KEYINPUT79), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n526), .A2(new_n527), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT78), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n526), .A2(new_n523), .A3(new_n527), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(G22gat), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n540), .A2(KEYINPUT82), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n534), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(KEYINPUT81), .B1(new_n539), .B2(new_n540), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT80), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n539), .A2(new_n545), .A3(new_n540), .ZN(new_n546));
  OAI211_X1 g345(.A(new_n540), .B(new_n518), .C1(new_n522), .C2(new_n528), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT80), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT81), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n529), .A2(new_n549), .A3(G22gat), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n544), .A2(new_n546), .A3(new_n548), .A4(new_n550), .ZN(new_n551));
  AOI221_X4 g350(.A(KEYINPUT83), .B1(new_n531), .B2(new_n543), .C1(new_n551), .C2(new_n534), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT83), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n534), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n543), .A2(new_n531), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n406), .B(new_n509), .C1(new_n552), .C2(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n401), .B1(new_n399), .B2(new_n400), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n404), .A2(new_n403), .A3(new_n398), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n534), .ZN(new_n561));
  AND3_X1   g360(.A1(new_n529), .A2(new_n549), .A3(G22gat), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n549), .B1(new_n529), .B2(G22gat), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n547), .B(new_n545), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n561), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n555), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT83), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n554), .A2(new_n553), .A3(new_n555), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n560), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT84), .B1(new_n492), .B2(new_n497), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT84), .ZN(new_n572));
  AOI211_X1 g371(.A(new_n572), .B(new_n496), .C1(new_n484), .C2(new_n491), .ZN(new_n573));
  NOR3_X1   g372(.A1(new_n498), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n574), .A2(new_n507), .ZN(new_n575));
  NOR3_X1   g374(.A1(new_n575), .A2(KEYINPUT35), .A3(new_n446), .ZN(new_n576));
  AOI22_X1  g375(.A1(KEYINPUT35), .A2(new_n557), .B1(new_n570), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n410), .A2(KEYINPUT37), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n444), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(KEYINPUT85), .B(KEYINPUT38), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n381), .A2(new_n411), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(new_n413), .ZN(new_n582));
  INV_X1    g381(.A(new_n414), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(KEYINPUT37), .B1(new_n584), .B2(new_n440), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n415), .A2(new_n430), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n580), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n431), .A2(new_n441), .ZN(new_n588));
  OAI22_X1  g387(.A1(new_n579), .A2(new_n587), .B1(new_n588), .B2(new_n410), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(KEYINPUT37), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n444), .A2(new_n578), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n580), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT39), .ZN(new_n594));
  NOR3_X1   g393(.A1(new_n471), .A2(new_n485), .A3(new_n489), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n472), .A2(new_n477), .A3(new_n482), .ZN(new_n596));
  AOI211_X1 g395(.A(new_n594), .B(new_n595), .C1(new_n596), .C2(new_n489), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n596), .A2(new_n594), .A3(new_n489), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(new_n496), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n600), .A2(KEYINPUT40), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT40), .ZN(new_n602));
  NOR3_X1   g401(.A1(new_n597), .A2(new_n599), .A3(new_n602), .ZN(new_n603));
  NOR4_X1   g402(.A1(new_n601), .A2(new_n571), .A3(new_n573), .A4(new_n603), .ZN(new_n604));
  AOI22_X1  g403(.A1(new_n575), .A2(new_n593), .B1(new_n604), .B2(new_n446), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n605), .B1(new_n552), .B2(new_n556), .ZN(new_n606));
  INV_X1    g405(.A(new_n446), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n502), .A2(new_n501), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n608), .A2(new_n499), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n607), .B1(new_n609), .B2(new_n507), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n568), .A2(new_n569), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT36), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n612), .B1(new_n402), .B2(new_n405), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n558), .A2(new_n559), .A3(KEYINPUT36), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AND3_X1   g414(.A1(new_n606), .A2(new_n611), .A3(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n577), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT18), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n206), .B1(new_n303), .B2(new_n305), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT90), .ZN(new_n620));
  AOI22_X1  g419(.A1(new_n619), .A2(new_n620), .B1(new_n206), .B2(new_n304), .ZN(new_n621));
  INV_X1    g420(.A(new_n206), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n306), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT90), .ZN(new_n624));
  NAND2_X1  g423(.A1(G229gat), .A2(G233gat), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n621), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  OR3_X1    g425(.A1(new_n304), .A2(KEYINPUT93), .A3(new_n206), .ZN(new_n627));
  OAI21_X1  g426(.A(KEYINPUT93), .B1(new_n304), .B2(new_n206), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n627), .B(new_n628), .C1(new_n622), .C2(new_n291), .ZN(new_n629));
  XNOR2_X1  g428(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(new_n625), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT94), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n629), .A2(KEYINPUT94), .A3(new_n631), .ZN(new_n635));
  AOI22_X1  g434(.A1(new_n618), .A2(new_n626), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n621), .A2(new_n624), .A3(KEYINPUT18), .A4(new_n625), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT91), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n636), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G113gat), .B(G141gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(G197gat), .ZN(new_n643));
  XOR2_X1   g442(.A(KEYINPUT11), .B(G169gat), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n645), .B(KEYINPUT12), .Z(new_n646));
  NAND2_X1  g445(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n646), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n636), .B(new_n648), .C1(new_n639), .C2(new_n640), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(KEYINPUT95), .B1(new_n617), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n557), .A2(KEYINPUT35), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n570), .A2(new_n576), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n606), .A2(new_n611), .A3(new_n615), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT95), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n657), .A2(new_n658), .A3(new_n650), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n341), .B1(new_n652), .B2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n609), .A2(new_n507), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g462(.A1(new_n660), .A2(new_n446), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT16), .B(G8gat), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(G8gat), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n667), .B1(new_n660), .B2(new_n446), .ZN(new_n668));
  OAI21_X1  g467(.A(KEYINPUT42), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT42), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n670), .B1(new_n664), .B2(new_n665), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(new_n671), .ZN(G1325gat));
  AOI21_X1  g471(.A(G15gat), .B1(new_n660), .B2(new_n406), .ZN(new_n673));
  INV_X1    g472(.A(new_n615), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(G15gat), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n675), .B(KEYINPUT108), .Z(new_n676));
  AOI21_X1  g475(.A(new_n673), .B1(new_n660), .B2(new_n676), .ZN(G1326gat));
  NOR2_X1   g476(.A1(new_n552), .A2(new_n556), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n660), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT43), .B(G22gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1327gat));
  INV_X1    g480(.A(KEYINPUT45), .ZN(new_n682));
  INV_X1    g481(.A(new_n247), .ZN(new_n683));
  INV_X1    g482(.A(new_n315), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n683), .A2(new_n684), .A3(new_n340), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n685), .B1(new_n652), .B2(new_n659), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n661), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n688), .A2(G29gat), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n682), .B1(new_n687), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n684), .B1(new_n577), .B2(new_n616), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI211_X1 g493(.A(KEYINPUT44), .B(new_n684), .C1(new_n577), .C2(new_n616), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n247), .A2(new_n651), .A3(new_n339), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n696), .A2(new_n661), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(G29gat), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n686), .A2(KEYINPUT45), .A3(new_n689), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n691), .A2(new_n699), .A3(new_n700), .ZN(G1328gat));
  NOR2_X1   g500(.A1(new_n607), .A2(new_n282), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  OR3_X1    g502(.A1(new_n687), .A2(KEYINPUT46), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n696), .A2(new_n446), .A3(new_n697), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(new_n282), .ZN(new_n706));
  OAI21_X1  g505(.A(KEYINPUT46), .B1(new_n687), .B2(new_n703), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n704), .A2(new_n706), .A3(new_n707), .ZN(G1329gat));
  NOR2_X1   g507(.A1(new_n560), .A2(G43gat), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  AOI211_X1 g509(.A(new_n685), .B(new_n710), .C1(new_n652), .C2(new_n659), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT47), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n694), .A2(new_n674), .A3(new_n695), .A4(new_n697), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(KEYINPUT111), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(G43gat), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n714), .A2(KEYINPUT111), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n713), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  AND3_X1   g517(.A1(new_n714), .A2(KEYINPUT110), .A3(G43gat), .ZN(new_n719));
  AOI21_X1  g518(.A(KEYINPUT110), .B1(new_n714), .B2(G43gat), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n719), .A2(new_n720), .A3(new_n711), .ZN(new_n721));
  XOR2_X1   g520(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n722));
  OAI21_X1  g521(.A(new_n718), .B1(new_n721), .B2(new_n722), .ZN(G1330gat));
  NAND4_X1  g522(.A1(new_n694), .A2(new_n678), .A3(new_n695), .A4(new_n697), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT48), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n724), .A2(new_n725), .A3(new_n288), .ZN(new_n726));
  INV_X1    g525(.A(new_n678), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n727), .A2(new_n288), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n686), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(KEYINPUT112), .A2(KEYINPUT48), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n726), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n686), .A2(KEYINPUT112), .A3(new_n728), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT113), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n724), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n288), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n724), .A2(new_n733), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n732), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n731), .B1(new_n737), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g537(.A1(new_n247), .A2(new_n315), .A3(new_n339), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n617), .A2(new_n650), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n661), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g541(.A(new_n446), .B(KEYINPUT114), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n743), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  XNOR2_X1  g547(.A(KEYINPUT115), .B(KEYINPUT116), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  OR3_X1    g549(.A1(new_n747), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n750), .B1(new_n747), .B2(new_n748), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(G1333gat));
  NAND2_X1  g552(.A1(new_n740), .A2(new_n674), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n560), .A2(G71gat), .ZN(new_n755));
  AOI22_X1  g554(.A1(new_n754), .A2(G71gat), .B1(new_n740), .B2(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g556(.A1(new_n740), .A2(new_n678), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g558(.A1(new_n247), .A2(new_n650), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n760), .B(new_n684), .C1(new_n577), .C2(new_n616), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n657), .A2(KEYINPUT51), .A3(new_n684), .A4(new_n760), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n340), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(G85gat), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n765), .A2(new_n766), .A3(new_n661), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n247), .A2(new_n650), .A3(new_n340), .ZN(new_n768));
  AND3_X1   g567(.A1(new_n696), .A2(new_n661), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n767), .B1(new_n769), .B2(new_n766), .ZN(G1336gat));
  NAND2_X1  g569(.A1(new_n696), .A2(new_n768), .ZN(new_n771));
  OAI21_X1  g570(.A(G92gat), .B1(new_n771), .B2(new_n743), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n743), .A2(G92gat), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT52), .B1(new_n765), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n696), .A2(new_n446), .A3(new_n768), .ZN(new_n776));
  AOI22_X1  g575(.A1(new_n776), .A2(G92gat), .B1(new_n765), .B2(new_n773), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n775), .B1(new_n777), .B2(new_n778), .ZN(G1337gat));
  OAI21_X1  g578(.A(G99gat), .B1(new_n771), .B2(new_n615), .ZN(new_n780));
  INV_X1    g579(.A(G99gat), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n765), .A2(new_n781), .A3(new_n406), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(G1338gat));
  NAND2_X1  g582(.A1(new_n763), .A2(new_n764), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT118), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n727), .A2(G106gat), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n784), .A2(new_n785), .A3(new_n339), .A4(new_n786), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n694), .A2(new_n678), .A3(new_n695), .A4(new_n768), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT117), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n788), .A2(new_n789), .A3(G106gat), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n785), .B1(new_n765), .B2(new_n786), .ZN(new_n792));
  OAI21_X1  g591(.A(KEYINPUT53), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AOI22_X1  g592(.A1(new_n788), .A2(G106gat), .B1(new_n789), .B2(KEYINPUT53), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n765), .A2(new_n786), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n794), .B1(new_n795), .B2(KEYINPUT53), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n793), .A2(new_n796), .ZN(G1339gat));
  NOR2_X1   g596(.A1(new_n341), .A2(new_n650), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n332), .B1(new_n334), .B2(new_n799), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n320), .A2(KEYINPUT106), .A3(new_n321), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT106), .B1(new_n320), .B2(new_n321), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n801), .A2(new_n802), .A3(new_n317), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n320), .A2(new_n317), .A3(new_n321), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(KEYINPUT54), .ZN(new_n805));
  OAI211_X1 g604(.A(KEYINPUT55), .B(new_n800), .C1(new_n803), .C2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n333), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n805), .B1(new_n324), .B2(new_n325), .ZN(new_n809));
  INV_X1    g608(.A(new_n800), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n808), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT119), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g612(.A(KEYINPUT119), .B(new_n808), .C1(new_n809), .C2(new_n810), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n807), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n625), .B1(new_n621), .B2(new_n624), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n629), .A2(new_n631), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n645), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n815), .A2(new_n684), .A3(new_n649), .A4(new_n818), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n339), .A2(new_n649), .A3(new_n818), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n820), .B1(new_n815), .B2(new_n650), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n819), .B1(new_n821), .B2(new_n684), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n798), .B1(new_n822), .B2(new_n683), .ZN(new_n823));
  INV_X1    g622(.A(new_n570), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n823), .A2(new_n688), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n743), .ZN(new_n826));
  OR3_X1    g625(.A1(new_n826), .A2(G113gat), .A3(new_n651), .ZN(new_n827));
  INV_X1    g626(.A(new_n798), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n806), .A2(new_n333), .ZN(new_n829));
  INV_X1    g628(.A(new_n814), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n800), .B1(new_n803), .B2(new_n805), .ZN(new_n831));
  AOI21_X1  g630(.A(KEYINPUT119), .B1(new_n831), .B2(new_n808), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n829), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n312), .A2(new_n314), .A3(new_n649), .A4(new_n818), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n820), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n836), .B1(new_n833), .B2(new_n651), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n835), .B1(new_n837), .B2(new_n315), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n828), .B1(new_n838), .B2(new_n247), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n743), .A2(new_n661), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(new_n560), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n839), .A2(new_n727), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(KEYINPUT120), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT120), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n839), .A2(new_n844), .A3(new_n727), .A4(new_n841), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n843), .A2(new_n650), .A3(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT121), .ZN(new_n847));
  AND3_X1   g646(.A1(new_n846), .A2(new_n847), .A3(G113gat), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n847), .B1(new_n846), .B2(G113gat), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n827), .B1(new_n848), .B2(new_n849), .ZN(G1340gat));
  INV_X1    g649(.A(new_n843), .ZN(new_n851));
  INV_X1    g650(.A(new_n845), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(G120gat), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n340), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n825), .A2(new_n339), .A3(new_n743), .ZN(new_n856));
  AOI22_X1  g655(.A1(new_n853), .A2(new_n855), .B1(new_n856), .B2(new_n854), .ZN(G1341gat));
  NOR3_X1   g656(.A1(new_n851), .A2(new_n683), .A3(new_n852), .ZN(new_n858));
  INV_X1    g657(.A(G127gat), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n247), .A2(new_n859), .ZN(new_n860));
  OAI22_X1  g659(.A1(new_n858), .A2(new_n859), .B1(new_n826), .B2(new_n860), .ZN(G1342gat));
  INV_X1    g660(.A(G134gat), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n315), .A2(new_n446), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n825), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  XOR2_X1   g663(.A(new_n864), .B(KEYINPUT56), .Z(new_n865));
  NOR3_X1   g664(.A1(new_n851), .A2(new_n315), .A3(new_n852), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n865), .B1(new_n866), .B2(new_n862), .ZN(G1343gat));
  INV_X1    g666(.A(KEYINPUT58), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n823), .A2(new_n688), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n674), .A2(new_n727), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n869), .A2(new_n743), .A3(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n452), .A3(new_n650), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n674), .A2(new_n840), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(KEYINPUT122), .ZN(new_n875));
  XOR2_X1   g674(.A(KEYINPUT123), .B(KEYINPUT57), .Z(new_n876));
  OAI21_X1  g675(.A(new_n876), .B1(new_n823), .B2(new_n727), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n650), .A2(new_n829), .A3(new_n811), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n684), .B1(new_n878), .B2(new_n836), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n683), .B1(new_n879), .B2(new_n835), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n828), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(KEYINPUT57), .A3(new_n678), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n875), .B1(new_n877), .B2(new_n882), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n883), .A2(new_n650), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n868), .B(new_n873), .C1(new_n884), .C2(new_n452), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n452), .B1(new_n883), .B2(new_n650), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n871), .A2(G141gat), .A3(new_n651), .ZN(new_n887));
  OAI21_X1  g686(.A(KEYINPUT58), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n885), .A2(new_n888), .ZN(G1344gat));
  NAND3_X1  g688(.A1(new_n872), .A2(new_n450), .A3(new_n339), .ZN(new_n890));
  AOI211_X1 g689(.A(KEYINPUT59), .B(new_n450), .C1(new_n883), .C2(new_n339), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n875), .A2(new_n340), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n823), .A2(new_n727), .A3(new_n876), .ZN(new_n894));
  AOI21_X1  g693(.A(KEYINPUT57), .B1(new_n881), .B2(new_n678), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n892), .B1(new_n896), .B2(G148gat), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n890), .B1(new_n891), .B2(new_n897), .ZN(G1345gat));
  NAND3_X1  g697(.A1(new_n872), .A2(new_n239), .A3(new_n247), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n883), .A2(new_n247), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n899), .B1(new_n900), .B2(new_n239), .ZN(G1346gat));
  NAND4_X1  g700(.A1(new_n869), .A2(new_n455), .A3(new_n863), .A4(new_n870), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n883), .A2(new_n684), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n902), .B1(new_n903), .B2(new_n455), .ZN(G1347gat));
  NOR2_X1   g703(.A1(new_n823), .A2(new_n661), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n824), .A2(new_n743), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(G169gat), .B1(new_n907), .B2(new_n650), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n661), .A2(new_n607), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n406), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n823), .A2(new_n678), .A3(new_n910), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n651), .A2(new_n355), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n908), .B1(new_n911), .B2(new_n912), .ZN(G1348gat));
  NAND2_X1  g712(.A1(new_n907), .A2(new_n339), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n356), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(KEYINPUT124), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n914), .A2(new_n917), .A3(new_n356), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n340), .A2(new_n356), .ZN(new_n919));
  AOI22_X1  g718(.A1(new_n916), .A2(new_n918), .B1(new_n911), .B2(new_n919), .ZN(G1349gat));
  INV_X1    g719(.A(new_n910), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n839), .A2(new_n727), .A3(new_n247), .A4(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(G183gat), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT126), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n683), .A2(new_n359), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n839), .A2(new_n688), .A3(new_n906), .A4(new_n925), .ZN(new_n926));
  AND3_X1   g725(.A1(new_n923), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n924), .B1(new_n923), .B2(new_n926), .ZN(new_n928));
  NAND2_X1  g727(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(new_n929), .ZN(new_n931));
  NOR4_X1   g730(.A1(new_n823), .A2(new_n678), .A3(new_n683), .A4(new_n910), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n926), .B1(new_n932), .B2(new_n362), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(KEYINPUT126), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n923), .A2(new_n924), .A3(new_n926), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n931), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n930), .A2(new_n936), .ZN(G1350gat));
  NAND3_X1  g736(.A1(new_n907), .A2(new_n372), .A3(new_n684), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n911), .A2(new_n684), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(G190gat), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n940), .A2(KEYINPUT61), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n940), .A2(KEYINPUT61), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n938), .B1(new_n941), .B2(new_n942), .ZN(G1351gat));
  NOR3_X1   g742(.A1(new_n674), .A2(new_n727), .A3(new_n743), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n905), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(G197gat), .B1(new_n945), .B2(new_n650), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n615), .A2(new_n909), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n881), .A2(new_n678), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT57), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(new_n876), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n839), .A2(new_n678), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n947), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n650), .A2(G197gat), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n946), .B1(new_n953), .B2(new_n954), .ZN(G1352gat));
  INV_X1    g754(.A(G204gat), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n956), .B1(new_n953), .B2(new_n339), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n340), .A2(G204gat), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n839), .A2(new_n688), .A3(new_n944), .A4(new_n958), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT62), .ZN(new_n960));
  OAI21_X1  g759(.A(KEYINPUT127), .B1(new_n957), .B2(new_n960), .ZN(new_n961));
  XOR2_X1   g760(.A(new_n959), .B(KEYINPUT62), .Z(new_n962));
  INV_X1    g761(.A(new_n947), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n963), .B1(new_n894), .B2(new_n895), .ZN(new_n964));
  OAI21_X1  g763(.A(G204gat), .B1(new_n964), .B2(new_n340), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT127), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n962), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n961), .A2(new_n967), .ZN(G1353gat));
  NAND3_X1  g767(.A1(new_n945), .A2(new_n427), .A3(new_n247), .ZN(new_n969));
  OAI211_X1 g768(.A(new_n247), .B(new_n963), .C1(new_n894), .C2(new_n895), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n970), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n971));
  AOI21_X1  g770(.A(KEYINPUT63), .B1(new_n970), .B2(G211gat), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(G1354gat));
  OAI21_X1  g772(.A(G218gat), .B1(new_n964), .B2(new_n315), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n945), .A2(new_n418), .A3(new_n684), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(G1355gat));
endmodule


