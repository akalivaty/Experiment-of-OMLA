//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 1 1 1 0 1 1 0 0 0 0 0 0 0 0 0 1 0 1 0 0 1 0 1 1 1 0 1 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n210, new_n211, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1224, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1289, new_n1290, new_n1291;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  NOR2_X1   g0009(.A1(G97), .A2(G107), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G87), .ZN(G355));
  INV_X1    g0012(.A(G1), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(G13), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n217), .B(G250), .C1(G257), .C2(G264), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT0), .Z(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  INV_X1    g0021(.A(G97), .ZN(new_n222));
  INV_X1    g0022(.A(G257), .ZN(new_n223));
  OAI22_X1  g0023(.A1(new_n220), .A2(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(G68), .B2(G238), .ZN(new_n225));
  INV_X1    g0025(.A(G107), .ZN(new_n226));
  INV_X1    g0026(.A(G264), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(G116), .B2(G270), .ZN(new_n229));
  INV_X1    g0029(.A(G226), .ZN(new_n230));
  INV_X1    g0030(.A(G77), .ZN(new_n231));
  INV_X1    g0031(.A(G244), .ZN(new_n232));
  OAI221_X1 g0032(.A(new_n229), .B1(new_n207), .B2(new_n230), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(G232), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n201), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g0035(.A(new_n216), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT1), .ZN(new_n237));
  NAND2_X1  g0037(.A1(G1), .A2(G13), .ZN(new_n238));
  NOR2_X1   g0038(.A1(new_n238), .A2(new_n214), .ZN(new_n239));
  NOR2_X1   g0039(.A1(new_n206), .A2(new_n207), .ZN(new_n240));
  AOI211_X1 g0040(.A(new_n219), .B(new_n237), .C1(new_n239), .C2(new_n240), .ZN(G361));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G232), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G238), .B(G244), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XNOR2_X1  g0045(.A(G250), .B(G257), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n227), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G270), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G358));
  XNOR2_X1  g0049(.A(G87), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G97), .B(G107), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(KEYINPUT65), .ZN(new_n253));
  XNOR2_X1  g0053(.A(G68), .B(G77), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n254), .B(new_n207), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n255), .B(G58), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n253), .B(new_n256), .ZN(G351));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(new_n220), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(KEYINPUT74), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT74), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT75), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n264), .B1(new_n258), .B2(KEYINPUT3), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT3), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(KEYINPUT75), .A3(G33), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n263), .A2(KEYINPUT3), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G1698), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n230), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n259), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n265), .A2(new_n267), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n269), .A2(G223), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT74), .B(G33), .ZN(new_n274));
  OAI211_X1 g0074(.A(new_n272), .B(new_n273), .C1(new_n266), .C2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT76), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n268), .A2(KEYINPUT76), .A3(new_n273), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n271), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G41), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n280), .A2(G1), .A3(G13), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT66), .B(G41), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n213), .B(G274), .C1(new_n285), .C2(G45), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n213), .B1(G41), .B2(G45), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n281), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G232), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n283), .A2(G179), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G169), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n291), .B1(new_n279), .B2(new_n282), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(KEYINPUT7), .B1(new_n268), .B2(G20), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n272), .B1(new_n266), .B2(new_n274), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT7), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n298), .A2(new_n299), .A3(new_n214), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n297), .A2(new_n300), .A3(G68), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n203), .B(new_n205), .C1(new_n201), .C2(new_n202), .ZN(new_n302));
  NOR2_X1   g0102(.A1(G20), .A2(G33), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n302), .A2(G20), .B1(G159), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n301), .A2(KEYINPUT16), .A3(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT16), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n260), .A2(new_n262), .A3(new_n266), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n309), .A2(KEYINPUT7), .A3(new_n214), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n266), .A2(G33), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n308), .ZN(new_n312));
  AOI21_X1  g0112(.A(KEYINPUT7), .B1(new_n312), .B2(new_n214), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n202), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n304), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n306), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n238), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n305), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n213), .A2(G13), .A3(G20), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n322), .A2(new_n319), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  XOR2_X1   g0124(.A(KEYINPUT8), .B(G58), .Z(new_n325));
  NAND2_X1  g0125(.A1(new_n213), .A2(G20), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n324), .A2(new_n327), .B1(new_n321), .B2(new_n325), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n320), .A2(new_n329), .ZN(new_n330));
  AND3_X1   g0130(.A1(new_n296), .A2(new_n330), .A3(KEYINPUT18), .ZN(new_n331));
  AOI21_X1  g0131(.A(KEYINPUT18), .B1(new_n296), .B2(new_n330), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT17), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n283), .A2(G190), .A3(new_n292), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n320), .A2(new_n335), .A3(new_n329), .ZN(new_n336));
  INV_X1    g0136(.A(G200), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n295), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n334), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n338), .ZN(new_n340));
  INV_X1    g0140(.A(new_n319), .ZN(new_n341));
  AOI21_X1  g0141(.A(G20), .B1(new_n307), .B2(new_n308), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n313), .B1(new_n342), .B2(KEYINPUT7), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n304), .B1(new_n343), .B2(new_n202), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n341), .B1(new_n344), .B2(new_n306), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n328), .B1(new_n345), .B2(new_n305), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n340), .A2(new_n346), .A3(KEYINPUT17), .A4(new_n335), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n339), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n333), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT77), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n349), .A2(new_n350), .ZN(new_n352));
  AND2_X1   g0152(.A1(new_n311), .A2(new_n308), .ZN(new_n353));
  NOR2_X1   g0153(.A1(G226), .A2(G1698), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n354), .B1(new_n234), .B2(G1698), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n353), .A2(new_n355), .B1(G33), .B2(G97), .ZN(new_n356));
  OR2_X1    g0156(.A1(new_n356), .A2(new_n281), .ZN(new_n357));
  XOR2_X1   g0157(.A(KEYINPUT73), .B(KEYINPUT13), .Z(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n289), .A2(G238), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n357), .A2(new_n286), .A3(new_n359), .A4(new_n360), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n286), .B(new_n360), .C1(new_n356), .C2(new_n281), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n358), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(G169), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(KEYINPUT14), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n362), .A2(KEYINPUT13), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n361), .A2(G179), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT14), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n364), .A2(new_n369), .A3(G169), .ZN(new_n370));
  AND3_X1   g0170(.A1(new_n366), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT69), .ZN(new_n372));
  XNOR2_X1  g0172(.A(new_n321), .B(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n373), .A2(new_n341), .A3(new_n326), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n202), .B1(new_n374), .B2(KEYINPUT12), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT12), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n375), .B1(new_n376), .B2(new_n321), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n322), .A2(new_n372), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n321), .A2(KEYINPUT69), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n380), .A2(KEYINPUT12), .A3(new_n202), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n214), .A2(G33), .ZN(new_n382));
  XNOR2_X1  g0182(.A(new_n382), .B(KEYINPUT67), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G77), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n303), .A2(G50), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n384), .B(new_n385), .C1(new_n214), .C2(G68), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT11), .ZN(new_n387));
  AND3_X1   g0187(.A1(new_n386), .A2(new_n387), .A3(new_n319), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n387), .B1(new_n386), .B2(new_n319), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n377), .B(new_n381), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n371), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  AND3_X1   g0193(.A1(new_n361), .A2(G190), .A3(new_n367), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n337), .B1(new_n361), .B2(new_n363), .ZN(new_n395));
  NOR3_X1   g0195(.A1(new_n390), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n352), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n269), .A2(G222), .ZN(new_n400));
  NAND2_X1  g0200(.A1(G223), .A2(G1698), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n353), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n402), .B(new_n282), .C1(G77), .C2(new_n353), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n403), .B(new_n286), .C1(new_n230), .C2(new_n288), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n404), .A2(G179), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n208), .A2(G20), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT68), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n383), .A2(new_n325), .B1(G150), .B2(new_n303), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n208), .A2(KEYINPUT68), .A3(G20), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n319), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n322), .A2(new_n207), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n323), .A2(G50), .A3(new_n326), .ZN(new_n414));
  AND3_X1   g0214(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  AOI211_X1 g0215(.A(new_n405), .B(new_n415), .C1(new_n294), .C2(new_n404), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n404), .A2(G200), .ZN(new_n417));
  INV_X1    g0217(.A(G190), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n404), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n419), .B1(new_n415), .B2(KEYINPUT9), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT9), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n421), .A2(KEYINPUT71), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(KEYINPUT71), .B1(new_n421), .B2(new_n422), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n417), .B(new_n420), .C1(new_n424), .C2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT10), .ZN(new_n427));
  INV_X1    g0227(.A(new_n425), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n423), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT10), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n429), .A2(new_n430), .A3(new_n417), .A4(new_n420), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n416), .B1(new_n427), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT72), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n282), .B1(new_n353), .B2(G107), .ZN(new_n434));
  NAND2_X1  g0234(.A1(G238), .A2(G1698), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(new_n234), .B2(G1698), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n312), .A2(new_n436), .ZN(new_n437));
  OAI221_X1 g0237(.A(new_n286), .B1(new_n232), .B2(new_n288), .C1(new_n434), .C2(new_n437), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n438), .A2(new_n294), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n438), .A2(G179), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT70), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  OR2_X1    g0241(.A1(new_n440), .A2(KEYINPUT70), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n325), .A2(new_n303), .B1(G20), .B2(G77), .ZN(new_n443));
  XNOR2_X1  g0243(.A(KEYINPUT15), .B(G87), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n443), .B1(new_n382), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n319), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n380), .A2(new_n231), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n446), .B(new_n447), .C1(new_n231), .C2(new_n374), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n441), .A2(new_n442), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n438), .A2(G200), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(new_n418), .B2(new_n438), .ZN(new_n451));
  OR2_X1    g0251(.A1(new_n451), .A2(new_n448), .ZN(new_n452));
  AND2_X1   g0252(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n432), .A2(new_n433), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n433), .B1(new_n432), .B2(new_n453), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n351), .B(new_n399), .C1(new_n455), .C2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n213), .A2(G33), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n321), .A2(new_n458), .A3(new_n238), .A4(new_n318), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n459), .A2(new_n444), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n380), .A2(new_n444), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n261), .A2(G33), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n258), .A2(KEYINPUT74), .ZN(new_n463));
  OAI21_X1  g0263(.A(KEYINPUT3), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n464), .A2(new_n214), .A3(G68), .A4(new_n272), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT19), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n466), .A2(new_n258), .A3(new_n222), .ZN(new_n467));
  XNOR2_X1  g0267(.A(KEYINPUT80), .B(G87), .ZN(new_n468));
  OAI22_X1  g0268(.A1(new_n467), .A2(G20), .B1(new_n468), .B2(new_n211), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n466), .B1(new_n382), .B2(new_n222), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n465), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AOI211_X1 g0271(.A(new_n460), .B(new_n461), .C1(new_n471), .C2(new_n319), .ZN(new_n472));
  NOR2_X1   g0272(.A1(G238), .A2(G1698), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n473), .B1(new_n232), .B2(G1698), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n464), .A2(new_n272), .A3(new_n474), .ZN(new_n475));
  AND3_X1   g0275(.A1(new_n260), .A2(new_n262), .A3(G116), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n281), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(G45), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n221), .B1(new_n479), .B2(G1), .ZN(new_n480));
  INV_X1    g0280(.A(G274), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n213), .A2(new_n481), .A3(G45), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n281), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT79), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n281), .A2(new_n480), .A3(new_n482), .A4(KEYINPUT79), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n294), .B1(new_n478), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G179), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n485), .A2(new_n486), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n476), .B1(new_n268), .B2(new_n474), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n489), .B(new_n490), .C1(new_n491), .C2(new_n281), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n472), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n220), .A2(G20), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n496), .A2(new_n311), .A3(new_n308), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT22), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n476), .A2(new_n214), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n464), .A2(KEYINPUT22), .A3(new_n272), .A4(new_n496), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT23), .ZN(new_n501));
  OAI211_X1 g0301(.A(G20), .B(new_n226), .C1(new_n501), .C2(KEYINPUT84), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n501), .A2(KEYINPUT84), .ZN(new_n503));
  XNOR2_X1  g0303(.A(new_n502), .B(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n499), .A2(new_n500), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(KEYINPUT24), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT24), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n499), .A2(new_n500), .A3(new_n504), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n319), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n221), .A2(new_n269), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n223), .A2(G1698), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n464), .A2(new_n272), .A3(new_n511), .A4(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n274), .A2(G294), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n282), .ZN(new_n516));
  AND2_X1   g0316(.A1(KEYINPUT66), .A2(G41), .ZN(new_n517));
  NOR2_X1   g0317(.A1(KEYINPUT66), .A2(G41), .ZN(new_n518));
  OR3_X1    g0318(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT5), .ZN(new_n519));
  INV_X1    g0319(.A(G41), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(KEYINPUT5), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n479), .A2(G1), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n519), .A2(G274), .A3(new_n521), .A4(new_n522), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n521), .B(new_n522), .C1(new_n284), .C2(KEYINPUT5), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n524), .A2(G264), .A3(new_n281), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n516), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G200), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n281), .B1(new_n513), .B2(new_n514), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n524), .A2(G264), .A3(new_n281), .ZN(new_n529));
  INV_X1    g0329(.A(new_n523), .ZN(new_n530));
  NOR3_X1   g0330(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(G190), .ZN(new_n532));
  AOI21_X1  g0332(.A(KEYINPUT25), .B1(new_n322), .B2(new_n226), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n322), .A2(KEYINPUT25), .A3(new_n226), .ZN(new_n535));
  INV_X1    g0335(.A(new_n459), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n534), .A2(new_n535), .B1(G107), .B2(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n510), .A2(new_n527), .A3(new_n532), .A4(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT4), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n539), .A2(G1698), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n540), .A2(new_n311), .A3(new_n308), .A4(G244), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G283), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n464), .A2(G244), .A3(new_n272), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n543), .B1(new_n544), .B2(new_n539), .ZN(new_n545));
  OAI21_X1  g0345(.A(KEYINPUT4), .B1(new_n312), .B2(new_n221), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(G1698), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n282), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n524), .A2(new_n281), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n523), .B1(new_n550), .B2(new_n223), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n549), .A2(G190), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n226), .A2(KEYINPUT6), .A3(G97), .ZN(new_n554));
  XOR2_X1   g0354(.A(G97), .B(G107), .Z(new_n555));
  OAI21_X1  g0355(.A(new_n554), .B1(new_n555), .B2(KEYINPUT6), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(G20), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n303), .A2(G77), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n557), .B(new_n558), .C1(new_n343), .C2(new_n226), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n321), .A2(new_n222), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n536), .B2(new_n222), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT78), .ZN(new_n562));
  OR2_X1    g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n562), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n559), .A2(new_n319), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n281), .B1(new_n545), .B2(new_n547), .ZN(new_n566));
  OAI21_X1  g0366(.A(G200), .B1(new_n566), .B2(new_n551), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n553), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(G200), .B1(new_n478), .B2(new_n487), .ZN(new_n569));
  OAI211_X1 g0369(.A(G190), .B(new_n490), .C1(new_n491), .C2(new_n281), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n471), .A2(new_n319), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n536), .A2(G87), .ZN(new_n573));
  INV_X1    g0373(.A(new_n461), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  OR2_X1    g0375(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n495), .A2(new_n538), .A3(new_n568), .A4(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n542), .B(new_n214), .C1(G33), .C2(new_n222), .ZN(new_n578));
  INV_X1    g0378(.A(G116), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(G20), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n319), .A2(KEYINPUT82), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(KEYINPUT82), .B1(new_n319), .B2(new_n580), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n578), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT20), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(KEYINPUT20), .B(new_n578), .C1(new_n581), .C2(new_n582), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n373), .A2(G116), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n579), .B1(new_n213), .B2(G33), .ZN(new_n590));
  AND4_X1   g0390(.A1(new_n341), .A2(new_n378), .A3(new_n379), .A4(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n587), .A2(new_n589), .A3(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n524), .A2(G270), .A3(new_n281), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n594), .A2(new_n523), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n223), .A2(new_n269), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n227), .A2(G1698), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n464), .A2(new_n272), .A3(new_n596), .A4(new_n597), .ZN(new_n598));
  XNOR2_X1  g0398(.A(KEYINPUT81), .B(G303), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n312), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n282), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n294), .B1(new_n595), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n593), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g0404(.A(KEYINPUT83), .B(KEYINPUT21), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n594), .A2(new_n523), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n281), .B1(new_n598), .B2(new_n600), .ZN(new_n607));
  OAI211_X1 g0407(.A(KEYINPUT21), .B(G169), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n595), .A2(new_n602), .A3(G179), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n604), .A2(new_n605), .B1(new_n610), .B2(new_n593), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n516), .A2(new_n489), .A3(new_n523), .A4(new_n525), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n341), .B1(new_n506), .B2(new_n508), .ZN(new_n613));
  INV_X1    g0413(.A(new_n537), .ZN(new_n614));
  OAI221_X1 g0414(.A(new_n612), .B1(new_n531), .B2(G169), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n559), .A2(new_n319), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n563), .A2(new_n564), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n549), .A2(new_n489), .A3(new_n552), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n294), .B1(new_n566), .B2(new_n551), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  AOI211_X1 g0421(.A(new_n588), .B(new_n591), .C1(new_n585), .C2(new_n586), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n606), .A2(new_n607), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(G190), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n622), .B(new_n624), .C1(new_n337), .C2(new_n623), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n611), .A2(new_n615), .A3(new_n621), .A4(new_n625), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n457), .A2(new_n577), .A3(new_n626), .ZN(G372));
  INV_X1    g0427(.A(new_n333), .ZN(new_n628));
  INV_X1    g0428(.A(new_n449), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n397), .B1(new_n392), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n628), .B1(new_n630), .B2(new_n348), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n427), .A2(new_n431), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n416), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT26), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n621), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n576), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT85), .ZN(new_n638));
  XNOR2_X1  g0438(.A(new_n575), .B(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n571), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n538), .A2(new_n568), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n642), .B1(new_n611), .B2(new_n615), .ZN(new_n643));
  INV_X1    g0443(.A(new_n621), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n637), .B1(new_n645), .B2(new_n634), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n646), .A2(new_n494), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n633), .B1(new_n457), .B2(new_n647), .ZN(G369));
  NAND3_X1  g0448(.A1(new_n213), .A2(new_n214), .A3(G13), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(G213), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(G343), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n611), .B(new_n625), .C1(new_n622), .C2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n610), .A2(new_n593), .ZN(new_n657));
  OAI21_X1  g0457(.A(G169), .B1(new_n606), .B2(new_n607), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n605), .B1(new_n622), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n660), .A2(new_n593), .A3(new_n654), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT86), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n662), .B(new_n663), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n664), .A2(G330), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n615), .A2(new_n654), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n613), .A2(new_n614), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n538), .B1(new_n667), .B2(new_n655), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n666), .B1(new_n615), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n611), .A2(new_n654), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(new_n666), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n670), .A2(new_n673), .ZN(G399));
  NAND2_X1  g0474(.A1(new_n217), .A2(new_n284), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G1), .ZN(new_n676));
  OR3_X1    g0476(.A1(new_n468), .A2(G116), .A3(new_n211), .ZN(new_n677));
  INV_X1    g0477(.A(new_n240), .ZN(new_n678));
  OAI22_X1  g0478(.A1(new_n676), .A2(new_n677), .B1(new_n678), .B2(new_n675), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n679), .B(KEYINPUT28), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT29), .ZN(new_n681));
  OAI22_X1  g0481(.A1(new_n472), .A2(new_n493), .B1(new_n571), .B2(new_n575), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n634), .B1(new_n621), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(KEYINPUT89), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n635), .A2(new_n641), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT89), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n686), .B(new_n634), .C1(new_n621), .C2(new_n682), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n684), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n495), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT90), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n688), .A2(KEYINPUT90), .A3(new_n495), .ZN(new_n692));
  INV_X1    g0492(.A(new_n641), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(new_n494), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n694), .A2(new_n643), .A3(new_n621), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n691), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n681), .B1(new_n696), .B2(new_n655), .ZN(new_n697));
  INV_X1    g0497(.A(G330), .ZN(new_n698));
  AND3_X1   g0498(.A1(new_n611), .A2(new_n615), .A3(new_n621), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n642), .A2(new_n682), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n699), .A2(new_n700), .A3(new_n625), .A4(new_n655), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT88), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n626), .A2(new_n577), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n704), .A2(KEYINPUT88), .A3(new_n655), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n528), .A2(new_n529), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n549), .A2(new_n707), .A3(new_n552), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n478), .A2(new_n487), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n623), .A2(new_n709), .A3(G179), .ZN(new_n710));
  NOR2_X1   g0510(.A1(KEYINPUT87), .A2(KEYINPUT30), .ZN(new_n711));
  OR3_X1    g0511(.A1(new_n708), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n566), .A2(new_n551), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n489), .B1(new_n478), .B2(new_n487), .ZN(new_n714));
  OR4_X1    g0514(.A1(new_n713), .A2(new_n531), .A3(new_n623), .A4(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n711), .B1(new_n708), .B2(new_n710), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n712), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n654), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(KEYINPUT31), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT31), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n717), .A2(new_n720), .A3(new_n654), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n698), .B1(new_n706), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n612), .B1(new_n531), .B2(G169), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n667), .A2(new_n724), .ZN(new_n725));
  OAI211_X1 g0525(.A(new_n568), .B(new_n538), .C1(new_n660), .C2(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n693), .B1(new_n726), .B2(new_n621), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n636), .B1(new_n727), .B2(KEYINPUT26), .ZN(new_n728));
  AOI211_X1 g0528(.A(KEYINPUT29), .B(new_n654), .C1(new_n728), .C2(new_n495), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n697), .A2(new_n723), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n680), .B1(new_n730), .B2(G1), .ZN(G364));
  INV_X1    g0531(.A(G13), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(G20), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n676), .B1(G45), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n665), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n735), .B1(G330), .B2(new_n664), .ZN(new_n736));
  XNOR2_X1  g0536(.A(new_n734), .B(KEYINPUT91), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n217), .A2(G355), .A3(new_n353), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n298), .A2(new_n217), .ZN(new_n740));
  XNOR2_X1  g0540(.A(new_n740), .B(KEYINPUT92), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n741), .B1(G45), .B2(new_n678), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n256), .A2(new_n479), .ZN(new_n743));
  OAI221_X1 g0543(.A(new_n739), .B1(G116), .B2(new_n217), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n214), .B1(KEYINPUT93), .B2(new_n294), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n294), .A2(KEYINPUT93), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n238), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G13), .A2(G33), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G20), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  AND2_X1   g0551(.A1(new_n744), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n489), .A2(new_n337), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n214), .A2(G190), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(G317), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(KEYINPUT33), .ZN(new_n758));
  OR2_X1    g0558(.A1(new_n757), .A2(KEYINPUT33), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n756), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G283), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n337), .A2(G179), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(new_n754), .ZN(new_n763));
  INV_X1    g0563(.A(G294), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G179), .A2(G200), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n214), .B1(new_n765), .B2(G190), .ZN(new_n766));
  OAI221_X1 g0566(.A(new_n760), .B1(new_n761), .B2(new_n763), .C1(new_n764), .C2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n489), .A2(G200), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n754), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n767), .B1(G311), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n214), .A2(new_n418), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(new_n753), .ZN(new_n773));
  INV_X1    g0573(.A(G326), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n312), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n754), .A2(new_n765), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n775), .B1(G329), .B2(new_n777), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n771), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G303), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n772), .A2(new_n762), .ZN(new_n781));
  INV_X1    g0581(.A(G322), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n772), .A2(new_n768), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n779), .B1(new_n780), .B2(new_n781), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n763), .A2(new_n226), .ZN(new_n785));
  INV_X1    g0585(.A(new_n781), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n312), .B(new_n785), .C1(new_n468), .C2(new_n786), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n787), .B(KEYINPUT95), .Z(new_n788));
  INV_X1    g0588(.A(new_n766), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n788), .B1(G97), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n756), .A2(G68), .ZN(new_n791));
  XOR2_X1   g0591(.A(KEYINPUT94), .B(G159), .Z(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n776), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT32), .ZN(new_n795));
  INV_X1    g0595(.A(new_n783), .ZN(new_n796));
  AOI22_X1  g0596(.A1(G58), .A2(new_n796), .B1(new_n770), .B2(G77), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n790), .A2(new_n791), .A3(new_n795), .A4(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n773), .A2(new_n207), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n784), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n752), .B1(new_n800), .B2(new_n747), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n750), .B(KEYINPUT96), .Z(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n738), .B(new_n801), .C1(new_n664), .C2(new_n803), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n736), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(G396));
  INV_X1    g0606(.A(G132), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n268), .B1(new_n807), .B2(new_n776), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G143), .A2(new_n796), .B1(new_n770), .B2(new_n792), .ZN(new_n809));
  INV_X1    g0609(.A(G137), .ZN(new_n810));
  INV_X1    g0610(.A(G150), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n809), .B1(new_n810), .B2(new_n773), .C1(new_n811), .C2(new_n755), .ZN(new_n812));
  XOR2_X1   g0612(.A(new_n812), .B(KEYINPUT34), .Z(new_n813));
  AOI211_X1 g0613(.A(new_n808), .B(new_n813), .C1(G50), .C2(new_n786), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n814), .B1(new_n201), .B2(new_n766), .C1(new_n202), .C2(new_n763), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n312), .B1(new_n769), .B2(new_n579), .C1(new_n220), .C2(new_n763), .ZN(new_n816));
  AOI22_X1  g0616(.A1(G311), .A2(new_n777), .B1(new_n789), .B2(G97), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n761), .B2(new_n755), .ZN(new_n818));
  INV_X1    g0618(.A(new_n773), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n816), .B(new_n818), .C1(G303), .C2(new_n819), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n820), .B1(new_n226), .B2(new_n781), .C1(new_n764), .C2(new_n783), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n815), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n737), .B1(new_n822), .B2(new_n747), .ZN(new_n823));
  INV_X1    g0623(.A(new_n747), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n749), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT97), .ZN(new_n826));
  OR3_X1    g0626(.A1(new_n449), .A2(KEYINPUT99), .A3(new_n655), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n448), .A2(new_n654), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT98), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n830), .A2(new_n449), .A3(new_n452), .ZN(new_n831));
  OAI21_X1  g0631(.A(KEYINPUT99), .B1(new_n449), .B2(new_n655), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n827), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n823), .B1(G77), .B2(new_n826), .C1(new_n749), .C2(new_n833), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n655), .B(new_n833), .C1(new_n646), .C2(new_n494), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n647), .A2(new_n654), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n833), .B(KEYINPUT100), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(new_n723), .Z(new_n839));
  OAI21_X1  g0639(.A(new_n834), .B1(new_n839), .B2(new_n734), .ZN(G384));
  INV_X1    g0640(.A(new_n457), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n697), .B2(new_n729), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n633), .ZN(new_n843));
  INV_X1    g0643(.A(new_n652), .ZN(new_n844));
  AOI21_X1  g0644(.A(KEYINPUT16), .B1(new_n301), .B2(new_n304), .ZN(new_n845));
  OAI21_X1  g0645(.A(KEYINPUT102), .B1(new_n845), .B2(new_n341), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT102), .ZN(new_n847));
  INV_X1    g0647(.A(new_n272), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n266), .B1(new_n260), .B2(new_n262), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n214), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n202), .B1(new_n850), .B2(KEYINPUT7), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n316), .B1(new_n851), .B2(new_n300), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n847), .B(new_n319), .C1(new_n852), .C2(KEYINPUT16), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n846), .A2(new_n853), .A3(new_n305), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n329), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n844), .B(new_n855), .C1(new_n333), .C2(new_n348), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n340), .A2(new_n346), .A3(new_n335), .ZN(new_n857));
  XNOR2_X1  g0657(.A(KEYINPUT103), .B(KEYINPUT37), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n296), .A2(new_n844), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n857), .B(new_n859), .C1(new_n860), .C2(new_n346), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n336), .A2(new_n338), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n294), .B1(new_n283), .B2(new_n292), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n489), .B(new_n291), .C1(new_n279), .C2(new_n282), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n652), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n862), .B1(new_n855), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT37), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n861), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n856), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT38), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n856), .A2(new_n869), .A3(KEYINPUT38), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n390), .A2(new_n654), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n397), .B(new_n875), .C1(new_n371), .C2(new_n391), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n366), .A2(new_n368), .A3(new_n370), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n390), .B(new_n654), .C1(new_n877), .C2(new_n396), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n827), .A2(new_n831), .A3(new_n832), .ZN(new_n880));
  AOI211_X1 g0680(.A(new_n654), .B(new_n880), .C1(new_n728), .C2(new_n495), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n449), .A2(new_n654), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n874), .B(new_n879), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n628), .A2(new_n844), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n330), .B(new_n844), .C1(new_n333), .C2(new_n348), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n346), .B1(new_n865), .B2(new_n652), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n858), .B1(new_n888), .B2(new_n862), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n889), .A2(new_n861), .A3(KEYINPUT104), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n888), .A2(new_n862), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT104), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n891), .A2(new_n892), .A3(new_n859), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n887), .A2(new_n890), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n871), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT39), .B1(new_n895), .B2(new_n873), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n856), .A2(new_n869), .A3(KEYINPUT38), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT38), .B1(new_n856), .B2(new_n869), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT39), .ZN(new_n899));
  NOR3_X1   g0699(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n393), .A2(new_n654), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n896), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n886), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n843), .B(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT88), .B1(new_n704), .B2(new_n655), .ZN(new_n906));
  NOR4_X1   g0706(.A1(new_n626), .A2(new_n577), .A3(new_n702), .A4(new_n654), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n722), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n841), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n879), .A2(new_n833), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(new_n706), .B2(new_n722), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT40), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n895), .B2(new_n873), .ZN(new_n913));
  INV_X1    g0713(.A(new_n910), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n908), .B(new_n914), .C1(new_n897), .C2(new_n898), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n911), .A2(new_n913), .B1(new_n915), .B2(new_n912), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n909), .B(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(G330), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n905), .B(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n213), .B2(new_n733), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n556), .B(KEYINPUT101), .Z(new_n921));
  AOI21_X1  g0721(.A(new_n579), .B1(new_n921), .B2(KEYINPUT35), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n922), .B(new_n239), .C1(KEYINPUT35), .C2(new_n921), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT36), .ZN(new_n924));
  OAI21_X1  g0724(.A(G77), .B1(new_n201), .B2(new_n202), .ZN(new_n925));
  OAI22_X1  g0725(.A1(new_n678), .A2(new_n925), .B1(G50), .B2(new_n202), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n926), .A2(G1), .A3(new_n732), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n920), .A2(new_n924), .A3(new_n927), .ZN(G367));
  OR2_X1    g0728(.A1(new_n639), .A2(new_n655), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n694), .A2(new_n929), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n929), .A2(new_n495), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(KEYINPUT43), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n621), .B(new_n568), .C1(new_n565), .C2(new_n655), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n934), .A2(KEYINPUT105), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(KEYINPUT105), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n935), .B(new_n936), .C1(new_n621), .C2(new_n655), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT106), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n725), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n654), .B1(new_n939), .B2(new_n621), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n937), .A2(new_n672), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT42), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n933), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n938), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n670), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n943), .B(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n932), .A2(KEYINPUT43), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n946), .B(new_n947), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n675), .B(KEYINPUT41), .Z(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n669), .B(new_n671), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n665), .B(new_n951), .ZN(new_n952));
  AND3_X1   g0752(.A1(new_n730), .A2(new_n952), .A3(KEYINPUT108), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT108), .B1(new_n730), .B2(new_n952), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT107), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n673), .A2(new_n937), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT44), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n673), .A2(new_n937), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT45), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n959), .B(new_n960), .ZN(new_n961));
  AND3_X1   g0761(.A1(new_n958), .A2(new_n670), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n670), .B1(new_n958), .B2(new_n961), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n956), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n955), .B(new_n964), .C1(new_n956), .C2(new_n963), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n950), .B1(new_n965), .B2(new_n730), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n733), .A2(G45), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(G1), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n948), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  AOI22_X1  g0769(.A1(G150), .A2(new_n796), .B1(new_n777), .B2(G137), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n970), .B1(new_n207), .B2(new_n769), .C1(new_n231), .C2(new_n763), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n766), .A2(new_n202), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n793), .A2(new_n755), .ZN(new_n973));
  INV_X1    g0773(.A(G143), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n353), .B1(new_n781), .B2(new_n201), .C1(new_n974), .C2(new_n773), .ZN(new_n975));
  NOR4_X1   g0775(.A1(new_n971), .A2(new_n972), .A3(new_n973), .A4(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n786), .A2(KEYINPUT46), .A3(G116), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT46), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n781), .B2(new_n579), .ZN(new_n979));
  INV_X1    g0779(.A(G311), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n977), .B(new_n979), .C1(new_n980), .C2(new_n773), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n763), .A2(new_n222), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n982), .B(new_n268), .C1(G294), .C2(new_n756), .ZN(new_n983));
  INV_X1    g0783(.A(new_n599), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n983), .B1(new_n761), .B2(new_n769), .C1(new_n984), .C2(new_n783), .ZN(new_n985));
  AOI211_X1 g0785(.A(new_n981), .B(new_n985), .C1(G317), .C2(new_n777), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n789), .A2(G107), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n976), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT47), .Z(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n747), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n930), .A2(new_n802), .A3(new_n931), .ZN(new_n991));
  INV_X1    g0791(.A(new_n741), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n751), .B1(new_n217), .B2(new_n444), .C1(new_n992), .C2(new_n248), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n990), .A2(new_n738), .A3(new_n991), .A4(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n969), .A2(new_n994), .ZN(G387));
  INV_X1    g0795(.A(new_n675), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n996), .B1(new_n730), .B2(new_n952), .C1(new_n953), .C2(new_n954), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n952), .A2(new_n968), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT109), .Z(new_n999));
  NOR2_X1   g0799(.A1(new_n766), .A2(new_n444), .ZN(new_n1000));
  INV_X1    g0800(.A(G159), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n773), .A2(new_n1001), .B1(new_n769), .B2(new_n202), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n1000), .B(new_n1002), .C1(G77), .C2(new_n786), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n777), .A2(G150), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n298), .B1(G50), .B2(new_n796), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n982), .B1(new_n325), .B2(new_n756), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n786), .A2(G294), .B1(new_n789), .B2(G283), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G322), .A2(new_n819), .B1(new_n756), .B2(G311), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n757), .B2(new_n783), .C1(new_n984), .C2(new_n769), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT48), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1008), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT111), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT49), .Z(new_n1016));
  OAI221_X1 g0816(.A(new_n298), .B1(new_n579), .B2(new_n763), .C1(new_n774), .C2(new_n776), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1007), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT112), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n747), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n325), .A2(new_n207), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1021), .B(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n479), .B1(new_n202), .B2(new_n231), .ZN(new_n1024));
  NOR3_X1   g0824(.A1(new_n1023), .A2(new_n677), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n245), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n741), .B1(new_n1026), .B2(new_n479), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n677), .A2(new_n217), .A3(new_n353), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1025), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n217), .A2(G107), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n751), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n669), .A2(new_n803), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1020), .A2(new_n738), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n997), .A2(new_n999), .A3(new_n1033), .ZN(G393));
  OAI22_X1  g0834(.A1(new_n953), .A2(new_n954), .B1(new_n962), .B2(new_n963), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n965), .A2(new_n1035), .A3(new_n996), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n962), .A2(new_n963), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n773), .A2(new_n811), .B1(new_n783), .B2(new_n1001), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT51), .Z(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(G143), .B2(new_n777), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n202), .B2(new_n781), .C1(new_n231), .C2(new_n766), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n756), .A2(G50), .B1(new_n770), .B2(new_n325), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT113), .Z(new_n1043));
  OAI211_X1 g0843(.A(new_n1043), .B(new_n268), .C1(new_n220), .C2(new_n763), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n769), .A2(new_n764), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n984), .A2(new_n755), .B1(new_n776), .B2(new_n782), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n1045), .B(new_n1046), .C1(G283), .C2(new_n786), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n773), .A2(new_n757), .B1(new_n783), .B2(new_n980), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT52), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n789), .A2(G116), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1047), .A2(new_n312), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n1041), .A2(new_n1044), .B1(new_n785), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n747), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n741), .A2(new_n252), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1054), .B(new_n751), .C1(new_n222), .C2(new_n217), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n738), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n944), .B2(new_n750), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n1037), .A2(new_n968), .B1(new_n1053), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1036), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT114), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1036), .A2(KEYINPUT114), .A3(new_n1058), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(G390));
  INV_X1    g0863(.A(new_n879), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n882), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1064), .B1(new_n835), .B2(new_n1065), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n1066), .A2(new_n901), .B1(new_n896), .B2(new_n900), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n908), .A2(G330), .A3(new_n833), .A4(new_n879), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n696), .A2(new_n655), .A3(new_n833), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1064), .B1(new_n1069), .B2(new_n1065), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n890), .A2(new_n893), .ZN(new_n1071));
  AOI21_X1  g0871(.A(KEYINPUT38), .B1(new_n1071), .B2(new_n887), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n902), .B1(new_n1072), .B2(new_n897), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1067), .B(new_n1068), .C1(new_n1070), .C2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n723), .A2(KEYINPUT115), .A3(new_n833), .A4(new_n879), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT115), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1068), .A2(new_n1076), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n879), .B1(new_n881), .B2(new_n882), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n899), .B1(new_n1072), .B2(new_n897), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n872), .A2(KEYINPUT39), .A3(new_n873), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n1079), .A2(new_n902), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1069), .A2(new_n1065), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1073), .B1(new_n1083), .B2(new_n879), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1078), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n352), .A2(new_n398), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n456), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1086), .B1(new_n1087), .B2(new_n454), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1088), .A2(G330), .A3(new_n351), .A4(new_n908), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n697), .A2(new_n729), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1089), .B(new_n633), .C1(new_n1090), .C2(new_n457), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n879), .B1(new_n723), .B2(new_n833), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n1078), .A2(new_n1092), .B1(new_n881), .B2(new_n882), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n723), .A2(new_n837), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n1064), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1095), .A2(new_n1065), .A3(new_n1069), .A4(new_n1068), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1091), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT116), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1074), .B(new_n1085), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1091), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1092), .B1(new_n1077), .B2(new_n1075), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n881), .A2(new_n882), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1096), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1085), .A2(new_n1074), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1104), .A2(new_n1105), .A3(KEYINPUT116), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1099), .A2(new_n996), .A3(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1085), .A2(new_n1074), .A3(new_n968), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n773), .A2(new_n761), .B1(new_n763), .B2(new_n202), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n764), .A2(new_n776), .B1(new_n766), .B2(new_n231), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n312), .B1(new_n783), .B2(new_n579), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n769), .A2(new_n222), .ZN(new_n1112));
  NOR4_X1   g0912(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .A4(new_n1112), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1113), .B1(new_n220), .B2(new_n781), .C1(new_n226), .C2(new_n755), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n781), .A2(new_n811), .ZN(new_n1115));
  XOR2_X1   g0915(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n1116));
  XNOR2_X1  g0916(.A(new_n1115), .B(new_n1116), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n783), .A2(new_n807), .B1(new_n763), .B2(new_n207), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(G128), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n773), .A2(new_n1120), .ZN(new_n1121));
  XOR2_X1   g0921(.A(KEYINPUT54), .B(G143), .Z(new_n1122));
  AOI211_X1 g0922(.A(new_n312), .B(new_n1121), .C1(new_n770), .C2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n777), .A2(G125), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n789), .A2(G159), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1119), .A2(new_n1123), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n755), .A2(new_n810), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1114), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n737), .B1(new_n1128), .B2(new_n747), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n896), .A2(new_n900), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1129), .B1(new_n325), .B2(new_n826), .C1(new_n1130), .C2(new_n749), .ZN(new_n1131));
  AND2_X1   g0931(.A1(new_n1108), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1107), .A2(new_n1132), .ZN(G378));
  XOR2_X1   g0933(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  OR2_X1    g0935(.A1(new_n432), .A2(new_n1135), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n415), .A2(new_n652), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n432), .A2(new_n1135), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n432), .A2(new_n1135), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n416), .B(new_n1134), .C1(new_n427), .C2(new_n431), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n1140), .A2(new_n1141), .B1(new_n415), .B2(new_n652), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1144), .A2(new_n749), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n734), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n826), .A2(G50), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n268), .A2(new_n285), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(G33), .A2(G41), .ZN(new_n1149));
  NOR3_X1   g0949(.A1(new_n1148), .A2(G50), .A3(new_n1149), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n769), .A2(new_n810), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n819), .A2(G125), .B1(new_n789), .B2(G150), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT119), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n1151), .B(new_n1153), .C1(new_n786), .C2(new_n1122), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n1154), .B1(new_n1120), .B2(new_n783), .C1(new_n807), .C2(new_n755), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1155), .B(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(G124), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n1149), .B1(new_n1158), .B2(new_n776), .C1(new_n793), .C2(new_n763), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1150), .B1(new_n1157), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n796), .A2(G107), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT118), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n781), .A2(new_n231), .B1(new_n769), .B2(new_n444), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n763), .A2(new_n201), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n776), .A2(new_n761), .ZN(new_n1166));
  NOR4_X1   g0966(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .A4(new_n972), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n1163), .A2(new_n1148), .A3(new_n1167), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n1168), .B1(new_n222), .B2(new_n755), .C1(new_n579), .C2(new_n773), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT58), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n824), .B1(new_n1161), .B2(new_n1170), .ZN(new_n1171));
  NOR4_X1   g0971(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .A4(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n915), .A2(new_n912), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n911), .B(KEYINPUT40), .C1(new_n1072), .C2(new_n897), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1173), .A2(new_n1174), .A3(G330), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(new_n1144), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n916), .A2(G330), .A3(new_n1143), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1176), .A2(new_n1177), .A3(KEYINPUT121), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(new_n904), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1130), .A2(new_n901), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1180), .A2(new_n885), .A3(new_n883), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1181), .A2(new_n1176), .A3(KEYINPUT121), .A4(new_n1177), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1172), .B1(new_n1183), .B2(new_n968), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1085), .A2(new_n1074), .A3(new_n1103), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1185), .A2(new_n1100), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1143), .B1(new_n916), .B2(G330), .ZN(new_n1187));
  AND4_X1   g0987(.A1(G330), .A2(new_n1173), .A3(new_n1174), .A4(new_n1143), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1181), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n904), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1189), .A2(new_n1190), .A3(KEYINPUT57), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n996), .B1(new_n1186), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1185), .A2(new_n1100), .ZN(new_n1193));
  AOI21_X1  g0993(.A(KEYINPUT57), .B1(new_n1183), .B2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1184), .B1(new_n1192), .B2(new_n1194), .ZN(G375));
  NAND2_X1  g0995(.A1(new_n1064), .A2(new_n748), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(G132), .A2(new_n819), .B1(new_n796), .B2(G137), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n1120), .B2(new_n776), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(G50), .B2(new_n789), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n1165), .B(new_n298), .C1(G150), .C2(new_n770), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n756), .A2(new_n1122), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n786), .A2(G159), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n773), .A2(new_n764), .B1(new_n783), .B2(new_n761), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n755), .A2(new_n579), .B1(new_n766), .B2(new_n444), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n781), .A2(new_n222), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n769), .A2(new_n226), .ZN(new_n1207));
  NOR4_X1   g1007(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n312), .B1(new_n763), .B2(new_n231), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT122), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n1208), .B(new_n1210), .C1(new_n780), .C2(new_n776), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n824), .B1(new_n1203), .B2(new_n1211), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n826), .A2(G68), .ZN(new_n1213));
  NOR3_X1   g1013(.A1(new_n1212), .A2(new_n737), .A3(new_n1213), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n1103), .A2(new_n968), .B1(new_n1196), .B2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n949), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1215), .B1(new_n1216), .B2(new_n1097), .ZN(G381));
  NAND4_X1  g1017(.A1(new_n1061), .A2(new_n969), .A3(new_n994), .A4(new_n1062), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(G393), .A2(G396), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NOR4_X1   g1020(.A1(new_n1218), .A2(G384), .A3(G381), .A4(new_n1220), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(G375), .A2(G378), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(G407));
  OAI21_X1  g1023(.A(new_n1222), .B1(new_n1221), .B2(new_n653), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(G213), .ZN(G409));
  NAND2_X1  g1025(.A1(G375), .A2(G378), .ZN(new_n1226));
  INV_X1    g1026(.A(G213), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1227), .A2(G343), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1189), .A2(new_n1190), .A3(new_n968), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n1179), .A2(new_n1182), .B1(new_n1185), .B2(new_n1100), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1231), .B1(new_n1232), .B2(new_n949), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1172), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1233), .A2(new_n1132), .A3(new_n1107), .A4(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT60), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1093), .A2(new_n1091), .A3(KEYINPUT60), .A4(new_n1096), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1237), .A2(new_n996), .A3(new_n1238), .A4(new_n1104), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1239), .A2(G384), .A3(new_n1215), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(G384), .B1(new_n1239), .B2(new_n1215), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1226), .A2(new_n1229), .A3(new_n1235), .A4(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(KEYINPUT123), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT63), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1228), .B1(G375), .B2(G378), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT123), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1247), .A2(new_n1248), .A3(new_n1235), .A4(new_n1243), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1245), .A2(new_n1246), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1239), .A2(new_n1215), .ZN(new_n1251));
  INV_X1    g1051(.A(G384), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n1240), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1228), .A2(G2897), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n1254), .B(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1247), .A2(new_n1235), .ZN(new_n1257));
  AOI21_X1  g1057(.A(KEYINPUT61), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT125), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1259), .B1(new_n1244), .B2(new_n1246), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1189), .A2(KEYINPUT57), .A3(new_n1190), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1193), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1262), .B(new_n996), .C1(new_n1232), .C2(KEYINPUT57), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n1263), .A2(new_n1184), .B1(new_n1132), .B2(new_n1107), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1183), .A2(new_n1193), .A3(new_n949), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1265), .A2(new_n1234), .A3(new_n1230), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(G378), .A2(new_n1266), .ZN(new_n1267));
  NOR3_X1   g1067(.A1(new_n1264), .A2(new_n1267), .A3(new_n1228), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1268), .A2(KEYINPUT125), .A3(KEYINPUT63), .A4(new_n1243), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1250), .A2(new_n1258), .A3(new_n1260), .A4(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(G390), .A2(G387), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT124), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(G393), .B(new_n805), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n1271), .A2(new_n1218), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1271), .A2(new_n1218), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(new_n1273), .B(new_n1272), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1274), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1270), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT62), .ZN(new_n1281));
  AND3_X1   g1081(.A1(new_n1245), .A2(new_n1281), .A3(new_n1249), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1268), .A2(KEYINPUT126), .A3(KEYINPUT62), .A4(new_n1243), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT126), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1284), .B1(new_n1244), .B2(new_n1281), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1283), .A2(new_n1285), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1278), .B(new_n1258), .C1(new_n1282), .C2(new_n1286), .ZN(new_n1287));
  AND2_X1   g1087(.A1(new_n1280), .A2(new_n1287), .ZN(G405));
  XNOR2_X1  g1088(.A(new_n1254), .B(KEYINPUT127), .ZN(new_n1289));
  OR2_X1    g1089(.A1(new_n1222), .A2(new_n1264), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(new_n1289), .B(new_n1290), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(new_n1291), .B(new_n1278), .ZN(G402));
endmodule


