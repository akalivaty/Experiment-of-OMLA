//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 1 0 0 0 0 0 0 1 0 1 1 0 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996;
  INV_X1    g000(.A(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G125), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G140), .ZN(new_n190));
  AND3_X1   g004(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT16), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT74), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT74), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n193), .B1(new_n188), .B2(KEYINPUT16), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n192), .B1(new_n191), .B2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n195), .B(G146), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n197));
  INV_X1    g011(.A(G119), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(G128), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(KEYINPUT23), .A3(G119), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n199), .B(new_n201), .C1(G119), .C2(new_n200), .ZN(new_n202));
  XNOR2_X1  g016(.A(G119), .B(G128), .ZN(new_n203));
  XOR2_X1   g017(.A(KEYINPUT24), .B(G110), .Z(new_n204));
  AOI22_X1  g018(.A1(new_n202), .A2(G110), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n196), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n195), .A2(G146), .ZN(new_n207));
  OAI22_X1  g021(.A1(new_n202), .A2(G110), .B1(new_n203), .B2(new_n204), .ZN(new_n208));
  AND2_X1   g022(.A1(new_n188), .A2(new_n190), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n207), .A2(new_n208), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n206), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G953), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(G221), .A3(G234), .ZN(new_n215));
  XNOR2_X1  g029(.A(new_n215), .B(KEYINPUT75), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT22), .B(G137), .ZN(new_n217));
  XNOR2_X1  g031(.A(new_n216), .B(new_n217), .ZN(new_n218));
  XOR2_X1   g032(.A(new_n218), .B(KEYINPUT76), .Z(new_n219));
  NAND2_X1  g033(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n206), .A2(new_n212), .A3(new_n218), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(G217), .A2(G902), .ZN(new_n223));
  INV_X1    g037(.A(G217), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n223), .B1(new_n224), .B2(G234), .ZN(new_n225));
  XOR2_X1   g039(.A(new_n225), .B(KEYINPUT73), .Z(new_n226));
  OR2_X1    g040(.A1(new_n226), .A2(G902), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT78), .B(KEYINPUT79), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n227), .B(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n222), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n231), .B1(new_n222), .B2(G902), .ZN(new_n232));
  INV_X1    g046(.A(G902), .ZN(new_n233));
  INV_X1    g047(.A(new_n231), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n220), .A2(new_n233), .A3(new_n221), .A4(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n230), .B1(new_n236), .B2(new_n226), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT31), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT71), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT0), .B(G128), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT65), .B1(new_n210), .B2(G143), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT65), .ZN(new_n244));
  INV_X1    g058(.A(G143), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n245), .A3(G146), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT64), .B1(new_n245), .B2(G146), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT64), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n249), .A2(new_n210), .A3(G143), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n242), .B1(new_n247), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n210), .A2(G143), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n245), .A2(G146), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n253), .A2(new_n254), .A3(KEYINPUT0), .A4(G128), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n241), .B1(new_n252), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT11), .ZN(new_n258));
  INV_X1    g072(.A(G134), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n258), .B1(new_n259), .B2(G137), .ZN(new_n260));
  INV_X1    g074(.A(G137), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n261), .A2(KEYINPUT11), .A3(G134), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n259), .A2(G137), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n260), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G131), .ZN(new_n265));
  INV_X1    g079(.A(G131), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n260), .A2(new_n262), .A3(new_n266), .A4(new_n263), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n242), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n248), .A2(new_n250), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n243), .A2(new_n246), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n272), .A2(KEYINPUT68), .A3(new_n255), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n257), .A2(new_n268), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT69), .ZN(new_n275));
  XOR2_X1   g089(.A(KEYINPUT2), .B(G113), .Z(new_n276));
  XNOR2_X1  g090(.A(G116), .B(G119), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n276), .B1(KEYINPUT67), .B2(new_n277), .ZN(new_n278));
  XOR2_X1   g092(.A(G116), .B(G119), .Z(new_n279));
  INV_X1    g093(.A(KEYINPUT67), .ZN(new_n280));
  XNOR2_X1  g094(.A(KEYINPUT2), .B(G113), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n253), .A2(KEYINPUT1), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G128), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n285), .B1(new_n270), .B2(new_n271), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n200), .A2(KEYINPUT1), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n287), .A2(new_n253), .A3(new_n254), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT66), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n287), .A2(new_n253), .A3(new_n254), .A4(KEYINPUT66), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n286), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n263), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n259), .A2(G137), .ZN(new_n295));
  OAI21_X1  g109(.A(G131), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(new_n267), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n283), .B1(new_n293), .B2(new_n298), .ZN(new_n299));
  AND3_X1   g113(.A1(new_n274), .A2(new_n275), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n275), .B1(new_n274), .B2(new_n299), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G237), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT70), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT70), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G237), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n307), .A2(G210), .A3(new_n214), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n308), .B(KEYINPUT27), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT26), .B(G101), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n309), .B(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n240), .B1(new_n302), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n274), .A2(new_n299), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT69), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n274), .A2(new_n275), .A3(new_n299), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n314), .A2(new_n240), .A3(new_n315), .A4(new_n311), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n251), .A2(new_n243), .A3(new_n246), .ZN(new_n317));
  AOI22_X1  g131(.A1(new_n317), .A2(new_n285), .B1(new_n290), .B2(new_n291), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n318), .A2(new_n297), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(new_n274), .A3(KEYINPUT30), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT30), .ZN(new_n322));
  INV_X1    g136(.A(new_n268), .ZN(new_n323));
  NOR3_X1   g137(.A1(new_n323), .A2(new_n252), .A3(new_n256), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n322), .B1(new_n324), .B2(new_n319), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n321), .A2(new_n325), .A3(new_n283), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n316), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n239), .B1(new_n312), .B2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n314), .A2(new_n315), .A3(new_n311), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT71), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n330), .A2(KEYINPUT31), .A3(new_n326), .A4(new_n316), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n283), .B1(new_n324), .B2(new_n319), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n314), .A2(new_n333), .A3(new_n315), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT28), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT72), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT28), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n336), .B1(new_n313), .B2(new_n337), .ZN(new_n338));
  AOI211_X1 g152(.A(KEYINPUT72), .B(KEYINPUT28), .C1(new_n274), .C2(new_n299), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n311), .B1(new_n335), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n332), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(G472), .A2(G902), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT32), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n302), .A2(new_n326), .ZN(new_n348));
  INV_X1    g162(.A(new_n311), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT29), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n335), .A2(new_n340), .A3(new_n311), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n320), .A2(new_n274), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n283), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n302), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT28), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n311), .A2(KEYINPUT29), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n340), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n352), .A2(new_n233), .A3(new_n358), .ZN(new_n359));
  AOI22_X1  g173(.A1(new_n343), .A2(new_n347), .B1(new_n359), .B2(G472), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n341), .B1(new_n328), .B2(new_n331), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n346), .B1(new_n361), .B2(new_n345), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n238), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G952), .ZN(new_n364));
  AOI211_X1 g178(.A(G953), .B(new_n364), .C1(G234), .C2(G237), .ZN(new_n365));
  AOI211_X1 g179(.A(new_n233), .B(new_n214), .C1(G234), .C2(G237), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT21), .B(G898), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(G210), .B1(G237), .B2(G902), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G104), .ZN(new_n371));
  OAI21_X1  g185(.A(KEYINPUT3), .B1(new_n371), .B2(G107), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT3), .ZN(new_n373));
  INV_X1    g187(.A(G107), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n374), .A3(G104), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n371), .A2(G107), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n372), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n377), .A2(G101), .ZN(new_n378));
  XNOR2_X1  g192(.A(KEYINPUT81), .B(KEYINPUT4), .ZN(new_n379));
  AOI22_X1  g193(.A1(new_n378), .A2(new_n379), .B1(new_n278), .B2(new_n282), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT80), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n377), .A2(G101), .ZN(new_n382));
  INV_X1    g196(.A(G101), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n372), .A2(new_n375), .A3(new_n383), .A4(new_n376), .ZN(new_n384));
  AND4_X1   g198(.A1(new_n381), .A2(new_n382), .A3(KEYINPUT4), .A4(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT4), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n386), .B1(new_n377), .B2(G101), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n381), .B1(new_n387), .B2(new_n384), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n380), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n376), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n371), .A2(G107), .ZN(new_n391));
  OAI21_X1  g205(.A(G101), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n384), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n276), .A2(new_n277), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT5), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(new_n198), .A3(G116), .ZN(new_n397));
  OAI211_X1 g211(.A(G113), .B(new_n397), .C1(new_n279), .C2(new_n396), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n394), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(G110), .B(G122), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n389), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT6), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n402), .A2(KEYINPUT85), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n400), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n377), .A2(G101), .A3(new_n379), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n283), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n382), .A2(KEYINPUT4), .A3(new_n384), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT80), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n387), .A2(new_n381), .A3(new_n384), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n407), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n394), .A2(new_n395), .A3(new_n398), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n405), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n404), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n400), .B1(new_n389), .B2(new_n399), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n403), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n286), .A2(new_n292), .A3(new_n189), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(KEYINPUT86), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT86), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n318), .A2(new_n419), .A3(new_n189), .ZN(new_n420));
  INV_X1    g234(.A(G224), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n421), .A2(G953), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(G125), .B1(new_n252), .B2(new_n256), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n418), .A2(new_n420), .A3(new_n423), .A4(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n424), .B1(new_n417), .B2(KEYINPUT86), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n419), .B1(new_n318), .B2(new_n189), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n422), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n414), .A2(new_n416), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT7), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n430), .B1(new_n426), .B2(new_n427), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n400), .B(KEYINPUT8), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n394), .B1(new_n395), .B2(new_n398), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n432), .B1(new_n412), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n428), .A2(new_n431), .A3(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n401), .B1(new_n425), .B2(new_n430), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n233), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n370), .B1(new_n429), .B2(new_n437), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n428), .A2(new_n431), .A3(new_n434), .ZN(new_n439));
  NOR3_X1   g253(.A1(new_n426), .A2(new_n427), .A3(new_n422), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n409), .A2(new_n410), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n412), .B1(new_n441), .B2(new_n380), .ZN(new_n442));
  AOI22_X1  g256(.A1(new_n440), .A2(KEYINPUT7), .B1(new_n442), .B2(new_n400), .ZN(new_n443));
  AOI21_X1  g257(.A(G902), .B1(new_n439), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n428), .A2(new_n425), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n415), .B1(new_n403), .B2(new_n401), .ZN(new_n446));
  INV_X1    g260(.A(new_n403), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n413), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n445), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n444), .A2(new_n449), .A3(new_n369), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n438), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(G214), .B1(G237), .B2(G902), .ZN(new_n452));
  AOI21_X1  g266(.A(KEYINPUT87), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT87), .ZN(new_n455));
  INV_X1    g269(.A(new_n452), .ZN(new_n456));
  AOI211_X1 g270(.A(new_n455), .B(new_n456), .C1(new_n438), .C2(new_n450), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n368), .B1(new_n454), .B2(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(G110), .B(G140), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n214), .A2(G227), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n460), .B(new_n461), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n441), .A2(new_n257), .A3(new_n273), .A4(new_n406), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n253), .A2(new_n254), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n285), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n393), .B1(new_n292), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT10), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n468), .B1(new_n286), .B2(new_n292), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n467), .A2(new_n468), .B1(new_n469), .B2(new_n394), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n463), .A2(new_n323), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n323), .B1(new_n463), .B2(new_n470), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n462), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n463), .A2(new_n470), .A3(new_n323), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT12), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n323), .B1(KEYINPUT82), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n293), .A2(new_n394), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n476), .B1(new_n477), .B2(new_n466), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n475), .A2(KEYINPUT82), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI221_X1 g294(.A(new_n476), .B1(KEYINPUT82), .B2(new_n475), .C1(new_n477), .C2(new_n466), .ZN(new_n481));
  INV_X1    g295(.A(new_n462), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n474), .A2(new_n480), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n473), .A2(KEYINPUT84), .A3(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(G469), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT84), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n486), .B(new_n462), .C1(new_n471), .C2(new_n472), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n484), .A2(new_n485), .A3(new_n233), .A4(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n474), .A2(new_n480), .A3(new_n481), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT83), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT83), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n474), .A2(new_n480), .A3(new_n481), .A4(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n490), .A2(new_n462), .A3(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n471), .A2(new_n472), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n482), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n493), .A2(new_n495), .A3(G469), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n485), .A2(new_n233), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n488), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  XNOR2_X1  g313(.A(KEYINPUT9), .B(G234), .ZN(new_n500));
  OAI21_X1  g314(.A(G221), .B1(new_n500), .B2(G902), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT20), .ZN(new_n503));
  XNOR2_X1  g317(.A(G113), .B(G122), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(new_n371), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n305), .A2(G237), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n303), .A2(KEYINPUT70), .ZN(new_n508));
  OAI211_X1 g322(.A(G214), .B(new_n214), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT88), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n307), .A2(KEYINPUT88), .A3(G214), .A4(new_n214), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n511), .A2(KEYINPUT89), .A3(new_n245), .A4(new_n512), .ZN(new_n513));
  OR2_X1    g327(.A1(new_n509), .A2(new_n245), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(G143), .B1(new_n509), .B2(new_n510), .ZN(new_n516));
  AOI21_X1  g330(.A(KEYINPUT89), .B1(new_n516), .B2(new_n512), .ZN(new_n517));
  OAI211_X1 g331(.A(KEYINPUT18), .B(G131), .C1(new_n515), .C2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n511), .A2(new_n245), .A3(new_n512), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT89), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(KEYINPUT18), .A2(G131), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n521), .A2(new_n514), .A3(new_n513), .A4(new_n522), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n209), .B(new_n210), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n518), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  XOR2_X1   g339(.A(new_n209), .B(KEYINPUT19), .Z(new_n526));
  OAI21_X1  g340(.A(new_n207), .B1(G146), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(G131), .B1(new_n515), .B2(new_n517), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n521), .A2(new_n266), .A3(new_n514), .A4(new_n513), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n506), .B1(new_n525), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n518), .A2(new_n523), .A3(new_n524), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT17), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n528), .A2(new_n533), .A3(new_n529), .ZN(new_n534));
  INV_X1    g348(.A(new_n196), .ZN(new_n535));
  OAI211_X1 g349(.A(KEYINPUT17), .B(G131), .C1(new_n515), .C2(new_n517), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n505), .B(new_n532), .C1(new_n534), .C2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n531), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(G475), .A2(G902), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n503), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n540), .ZN(new_n542));
  AOI211_X1 g356(.A(KEYINPUT20), .B(new_n542), .C1(new_n531), .C2(new_n538), .ZN(new_n543));
  INV_X1    g357(.A(G475), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n532), .B1(new_n534), .B2(new_n537), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n506), .ZN(new_n546));
  AOI21_X1  g360(.A(G902), .B1(new_n546), .B2(new_n538), .ZN(new_n547));
  OAI22_X1  g361(.A1(new_n541), .A2(new_n543), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(G116), .B(G122), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT14), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(G122), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n552), .A2(G116), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n374), .B1(new_n553), .B2(KEYINPUT14), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n552), .A2(G116), .ZN(new_n555));
  INV_X1    g369(.A(G116), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(G122), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n555), .A2(new_n557), .A3(new_n374), .ZN(new_n558));
  AOI22_X1  g372(.A1(new_n551), .A2(new_n554), .B1(KEYINPUT94), .B2(new_n558), .ZN(new_n559));
  OR2_X1    g373(.A1(new_n558), .A2(KEYINPUT94), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT90), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n561), .B1(new_n200), .B2(G143), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n245), .A2(KEYINPUT90), .A3(G128), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT92), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n565), .B1(new_n245), .B2(G128), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n200), .A2(KEYINPUT92), .A3(G143), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n564), .A2(new_n568), .A3(new_n259), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n259), .B1(new_n564), .B2(new_n568), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n559), .B(new_n560), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n500), .A2(new_n224), .A3(G953), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n549), .B(new_n374), .ZN(new_n574));
  AOI22_X1  g388(.A1(new_n562), .A2(new_n563), .B1(new_n566), .B2(new_n567), .ZN(new_n575));
  AOI21_X1  g389(.A(KEYINPUT93), .B1(new_n575), .B2(new_n259), .ZN(new_n576));
  AND4_X1   g390(.A1(KEYINPUT93), .A2(new_n564), .A3(new_n568), .A4(new_n259), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n574), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(KEYINPUT91), .B(KEYINPUT13), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n568), .B1(new_n564), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT13), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(KEYINPUT91), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT91), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(KEYINPUT13), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n586), .B1(new_n562), .B2(new_n563), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n259), .B1(new_n581), .B2(new_n588), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n572), .B(new_n573), .C1(new_n578), .C2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT95), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT93), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n569), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n575), .A2(KEYINPUT93), .A3(new_n259), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(G134), .B1(new_n580), .B2(new_n587), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(new_n597), .A3(new_n574), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n573), .B1(new_n598), .B2(new_n572), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n592), .A2(new_n599), .ZN(new_n600));
  AOI211_X1 g414(.A(new_n591), .B(new_n573), .C1(new_n598), .C2(new_n572), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(G478), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(KEYINPUT15), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n602), .A2(new_n233), .A3(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n599), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n607), .A2(new_n591), .A3(new_n590), .ZN(new_n608));
  INV_X1    g422(.A(new_n601), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n608), .A2(new_n609), .A3(new_n233), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n604), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n502), .A2(new_n548), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n363), .A2(new_n459), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(G101), .ZN(G3));
  NAND2_X1  g429(.A1(new_n343), .A2(new_n344), .ZN(new_n616));
  OAI21_X1  g430(.A(G472), .B1(new_n361), .B2(G902), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n499), .A2(new_n237), .A3(new_n501), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n590), .B1(new_n599), .B2(KEYINPUT97), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT97), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n598), .A2(new_n622), .A3(new_n572), .A4(new_n573), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(KEYINPUT33), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n626), .B1(new_n600), .B2(new_n601), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n603), .B1(new_n628), .B2(new_n233), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n610), .A2(G478), .ZN(new_n630));
  OAI21_X1  g444(.A(KEYINPUT98), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n630), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT98), .ZN(new_n633));
  AOI21_X1  g447(.A(G902), .B1(new_n625), .B2(new_n627), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n632), .B(new_n633), .C1(new_n634), .C2(new_n603), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n548), .A2(new_n631), .A3(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n451), .A2(new_n452), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT96), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n451), .A2(KEYINPUT96), .A3(new_n452), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n368), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n620), .A2(new_n637), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT34), .B(G104), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G6));
  AOI211_X1 g459(.A(KEYINPUT99), .B(new_n503), .C1(new_n539), .C2(new_n540), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n541), .A2(new_n543), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n646), .B1(new_n647), .B2(KEYINPUT99), .ZN(new_n648));
  INV_X1    g462(.A(new_n538), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n528), .A2(new_n533), .A3(new_n529), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n650), .A2(new_n535), .A3(new_n536), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n505), .B1(new_n651), .B2(new_n532), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n233), .B1(new_n649), .B2(new_n652), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n653), .A2(G475), .B1(new_n611), .B2(new_n606), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n648), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n620), .A2(new_n655), .A3(new_n642), .ZN(new_n656));
  XOR2_X1   g470(.A(new_n656), .B(KEYINPUT100), .Z(new_n657));
  XOR2_X1   g471(.A(KEYINPUT35), .B(G107), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G9));
  NAND2_X1  g473(.A1(new_n236), .A2(new_n226), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n219), .A2(KEYINPUT36), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(new_n213), .ZN(new_n662));
  INV_X1    g476(.A(new_n229), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n616), .A2(new_n617), .A3(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT101), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n616), .A2(new_n617), .A3(new_n665), .A4(KEYINPUT101), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n668), .A2(new_n459), .A3(new_n613), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT37), .B(G110), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT102), .B(KEYINPUT103), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G12));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n365), .B(KEYINPUT104), .Z(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(G900), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n677), .B1(new_n678), .B2(new_n366), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n648), .A2(new_n675), .A3(new_n654), .A4(new_n680), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n502), .B1(new_n640), .B2(new_n641), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n660), .A2(new_n664), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n683), .B1(new_n360), .B2(new_n362), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n539), .A2(new_n540), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(KEYINPUT20), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n539), .A2(new_n503), .A3(new_n540), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n686), .A2(KEYINPUT99), .A3(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT99), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n541), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n688), .A2(new_n690), .A3(new_n654), .A4(new_n680), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(KEYINPUT105), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n681), .A2(new_n682), .A3(new_n684), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G128), .ZN(G30));
  XOR2_X1   g508(.A(new_n679), .B(KEYINPUT39), .Z(new_n695));
  NAND3_X1  g509(.A1(new_n499), .A2(new_n501), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT107), .ZN(new_n697));
  XOR2_X1   g511(.A(new_n697), .B(KEYINPUT40), .Z(new_n698));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n330), .A2(new_n326), .A3(new_n316), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n355), .A2(new_n349), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n233), .ZN(new_n705));
  AOI22_X1  g519(.A1(new_n343), .A2(new_n347), .B1(G472), .B2(new_n705), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n665), .B1(new_n706), .B2(new_n362), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n548), .A2(new_n612), .ZN(new_n708));
  XNOR2_X1  g522(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n451), .B(new_n709), .ZN(new_n710));
  AND4_X1   g524(.A1(new_n452), .A2(new_n707), .A3(new_n708), .A4(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n700), .A2(new_n701), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G143), .ZN(G45));
  NAND4_X1  g527(.A1(new_n548), .A2(new_n631), .A3(new_n635), .A4(new_n680), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n682), .A2(new_n684), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G146), .ZN(G48));
  NAND3_X1  g531(.A1(new_n484), .A2(new_n233), .A3(new_n487), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(G469), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n501), .A3(new_n488), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n363), .A2(new_n637), .A3(new_n642), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT41), .B(G113), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G15));
  NAND4_X1  g538(.A1(new_n655), .A2(new_n363), .A3(new_n642), .A4(new_n721), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G116), .ZN(G18));
  AOI21_X1  g540(.A(new_n720), .B1(new_n640), .B2(new_n641), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n548), .A2(new_n368), .A3(new_n612), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n684), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G119), .ZN(G21));
  AND2_X1   g544(.A1(new_n356), .A2(new_n340), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n332), .B1(new_n311), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n344), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n733), .A2(new_n237), .A3(new_n617), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n640), .A2(new_n641), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n720), .A2(new_n368), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n734), .A2(new_n735), .A3(new_n708), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  NAND3_X1  g552(.A1(new_n733), .A2(new_n617), .A3(new_n665), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n739), .A2(new_n714), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n727), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G125), .ZN(G27));
  XNOR2_X1  g556(.A(KEYINPUT110), .B(KEYINPUT42), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n343), .A2(new_n347), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n359), .A2(G472), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n744), .A2(new_n362), .A3(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n438), .A2(new_n450), .A3(new_n452), .A4(new_n501), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n488), .A2(new_n498), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n493), .A2(KEYINPUT109), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n482), .B1(new_n489), .B2(KEYINPUT83), .ZN(new_n750));
  AOI22_X1  g564(.A1(new_n750), .A2(new_n492), .B1(new_n482), .B2(new_n494), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n749), .B(G469), .C1(new_n751), .C2(KEYINPUT109), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n747), .B1(new_n748), .B2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n746), .A2(new_n753), .A3(new_n237), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n743), .B1(new_n754), .B2(new_n714), .ZN(new_n755));
  NOR2_X1   g569(.A1(KEYINPUT110), .A2(KEYINPUT42), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n363), .A2(new_n715), .A3(new_n753), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT111), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT111), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n755), .A2(new_n761), .A3(new_n758), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G131), .ZN(G33));
  NAND3_X1  g578(.A1(new_n681), .A2(new_n692), .A3(KEYINPUT112), .ZN(new_n765));
  INV_X1    g579(.A(new_n754), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT112), .B1(new_n681), .B2(new_n692), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XOR2_X1   g583(.A(KEYINPUT113), .B(G134), .Z(new_n770));
  XNOR2_X1  g584(.A(new_n769), .B(new_n770), .ZN(G36));
  AOI22_X1  g585(.A1(new_n686), .A2(new_n687), .B1(G475), .B2(new_n653), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(new_n631), .A3(new_n635), .ZN(new_n773));
  XOR2_X1   g587(.A(new_n773), .B(KEYINPUT43), .Z(new_n774));
  NAND3_X1  g588(.A1(new_n774), .A2(new_n618), .A3(new_n665), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT44), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XOR2_X1   g591(.A(new_n777), .B(KEYINPUT114), .Z(new_n778));
  OAI21_X1  g592(.A(G469), .B1(new_n751), .B2(KEYINPUT45), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n751), .A2(KEYINPUT109), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n780), .B1(KEYINPUT109), .B2(new_n493), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n779), .B1(new_n781), .B2(KEYINPUT45), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n782), .A2(new_n497), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n783), .A2(KEYINPUT46), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n488), .B1(new_n783), .B2(KEYINPUT46), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n501), .B(new_n695), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n451), .A2(new_n456), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n789), .B1(new_n775), .B2(new_n776), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n778), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(new_n261), .ZN(G39));
  OAI21_X1  g607(.A(new_n501), .B1(new_n784), .B2(new_n785), .ZN(new_n794));
  XNOR2_X1  g608(.A(KEYINPUT115), .B(KEYINPUT47), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n794), .A2(new_n796), .ZN(new_n798));
  NOR4_X1   g612(.A1(new_n746), .A2(new_n714), .A3(new_n237), .A4(new_n789), .ZN(new_n799));
  XOR2_X1   g613(.A(new_n799), .B(KEYINPUT116), .Z(new_n800));
  NAND3_X1  g614(.A1(new_n797), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G140), .ZN(G42));
  NAND2_X1  g616(.A1(new_n364), .A2(new_n214), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(KEYINPUT123), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT121), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n774), .A2(new_n677), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(new_n734), .ZN(new_n807));
  OR3_X1    g621(.A1(new_n710), .A2(new_n452), .A3(new_n720), .ZN(new_n808));
  OR4_X1    g622(.A1(new_n805), .A2(new_n807), .A3(KEYINPUT50), .A4(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(KEYINPUT121), .B(KEYINPUT50), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n810), .B1(new_n807), .B2(new_n808), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n789), .A2(new_n720), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n806), .A2(new_n812), .ZN(new_n813));
  OR2_X1    g627(.A1(new_n813), .A2(new_n739), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n706), .A2(new_n362), .ZN(new_n815));
  AND4_X1   g629(.A1(new_n237), .A2(new_n815), .A3(new_n365), .A4(new_n812), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n548), .B1(new_n631), .B2(new_n635), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n809), .A2(new_n811), .A3(new_n814), .A4(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT51), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n719), .A2(new_n488), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(new_n501), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n822), .B1(new_n797), .B2(new_n798), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n806), .A2(new_n734), .A3(new_n788), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OR3_X1    g639(.A1(new_n819), .A2(new_n820), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n820), .B1(new_n819), .B2(new_n825), .ZN(new_n827));
  AOI211_X1 g641(.A(new_n364), .B(G953), .C1(new_n816), .C2(new_n637), .ZN(new_n828));
  INV_X1    g642(.A(new_n727), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n828), .B1(new_n807), .B2(new_n829), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n806), .A2(new_n363), .A3(new_n812), .ZN(new_n831));
  AND2_X1   g645(.A1(KEYINPUT122), .A2(KEYINPUT48), .ZN(new_n832));
  NOR2_X1   g646(.A1(KEYINPUT122), .A2(KEYINPUT48), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  AOI211_X1 g648(.A(new_n830), .B(new_n834), .C1(new_n831), .C2(new_n832), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n826), .A2(new_n827), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT119), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n740), .A2(new_n753), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n606), .A2(new_n611), .A3(new_n680), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n839), .B1(G475), .B2(new_n653), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n788), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n688), .A2(new_n690), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n841), .A2(new_n842), .A3(new_n502), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(new_n684), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n838), .A2(new_n844), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n765), .A2(new_n766), .ZN(new_n846));
  INV_X1    g660(.A(new_n768), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n670), .A2(new_n722), .A3(new_n614), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT118), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n636), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n548), .A2(new_n631), .A3(KEYINPUT118), .A4(new_n635), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n772), .A2(new_n612), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n368), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n855), .B1(new_n453), .B2(new_n457), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n856), .A2(new_n618), .A3(new_n619), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n849), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n725), .A2(new_n729), .A3(new_n737), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n848), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n762), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n761), .B1(new_n755), .B2(new_n758), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n837), .B1(new_n862), .B2(new_n865), .ZN(new_n866));
  AOI22_X1  g680(.A1(new_n740), .A2(new_n753), .B1(new_n843), .B2(new_n684), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n867), .B1(new_n767), .B2(new_n768), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n854), .A2(new_n857), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n869), .A2(new_n614), .A3(new_n670), .A4(new_n722), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n868), .A2(new_n870), .A3(new_n860), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n871), .A2(KEYINPUT119), .A3(new_n763), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n693), .A2(new_n741), .A3(new_n716), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n680), .A2(new_n501), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n874), .B1(new_n748), .B2(new_n752), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n707), .A2(new_n735), .A3(new_n708), .A4(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n873), .A2(KEYINPUT120), .A3(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n693), .A2(new_n741), .A3(new_n876), .A4(new_n716), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT120), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT52), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n877), .A2(KEYINPUT52), .A3(new_n880), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n866), .A2(new_n872), .A3(new_n883), .A4(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT53), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n870), .A2(new_n860), .ZN(new_n887));
  AND4_X1   g701(.A1(KEYINPUT119), .A2(new_n763), .A3(new_n887), .A4(new_n848), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT119), .B1(new_n871), .B2(new_n763), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(KEYINPUT52), .B1(new_n877), .B2(new_n880), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n878), .A2(KEYINPUT52), .ZN(new_n893));
  OR3_X1    g707(.A1(new_n892), .A2(KEYINPUT53), .A3(new_n893), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n886), .B(KEYINPUT54), .C1(new_n891), .C2(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n887), .A2(KEYINPUT53), .A3(new_n759), .A4(new_n848), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n892), .A2(new_n896), .A3(new_n893), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT53), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n897), .B1(new_n885), .B2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT54), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n895), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n804), .B1(new_n836), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n821), .A2(KEYINPUT49), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT117), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n237), .A2(new_n452), .A3(new_n501), .ZN(new_n906));
  AOI211_X1 g720(.A(new_n906), .B(new_n710), .C1(KEYINPUT49), .C2(new_n821), .ZN(new_n907));
  INV_X1    g721(.A(new_n773), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n907), .A2(new_n815), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n903), .B1(new_n905), .B2(new_n909), .ZN(G75));
  NOR2_X1   g724(.A1(new_n899), .A2(new_n233), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(G210), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n446), .A2(new_n448), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(new_n445), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT55), .ZN(new_n915));
  XOR2_X1   g729(.A(KEYINPUT124), .B(KEYINPUT56), .Z(new_n916));
  AND3_X1   g730(.A1(new_n912), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT56), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n915), .B1(new_n912), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n214), .A2(G952), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n917), .A2(new_n919), .A3(new_n920), .ZN(G51));
  INV_X1    g735(.A(KEYINPUT125), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(new_n899), .B2(new_n900), .ZN(new_n923));
  INV_X1    g737(.A(new_n884), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n924), .A2(new_n892), .ZN(new_n925));
  AOI21_X1  g739(.A(KEYINPUT53), .B1(new_n890), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(KEYINPUT54), .B1(new_n926), .B2(new_n897), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n922), .B(KEYINPUT54), .C1(new_n926), .C2(new_n897), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n497), .B(KEYINPUT57), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n484), .A2(new_n487), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n911), .A2(new_n782), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n920), .B1(new_n933), .B2(new_n934), .ZN(G54));
  AND2_X1   g749(.A1(KEYINPUT58), .A2(G475), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n911), .A2(new_n539), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n539), .B1(new_n911), .B2(new_n936), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n937), .A2(new_n938), .A3(new_n920), .ZN(G60));
  NAND2_X1  g753(.A1(G478), .A2(G902), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT59), .Z(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n628), .B(KEYINPUT126), .ZN(new_n943));
  AND4_X1   g757(.A1(new_n929), .A2(new_n928), .A3(new_n942), .A4(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n920), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n941), .B1(new_n895), .B2(new_n901), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n945), .B1(new_n946), .B2(new_n943), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n944), .A2(new_n947), .ZN(G63));
  XNOR2_X1  g762(.A(new_n223), .B(KEYINPUT60), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n662), .B(new_n950), .C1(new_n926), .C2(new_n897), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n222), .B1(new_n899), .B2(new_n949), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n951), .A2(new_n952), .A3(new_n945), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT61), .ZN(new_n954));
  OR2_X1    g768(.A1(new_n954), .A2(KEYINPUT127), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(KEYINPUT127), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n953), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n956), .B1(new_n953), .B2(new_n955), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n957), .A2(new_n958), .ZN(G66));
  OAI21_X1  g773(.A(G953), .B1(new_n367), .B2(new_n421), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n960), .B1(new_n887), .B2(G953), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n913), .B1(G898), .B2(new_n214), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(G69));
  AOI21_X1  g777(.A(new_n214), .B1(G227), .B2(G900), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n697), .A2(new_n854), .A3(new_n363), .A4(new_n788), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n801), .B(new_n965), .C1(new_n778), .C2(new_n791), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT62), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n967), .B1(new_n712), .B2(new_n873), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n712), .A2(new_n967), .A3(new_n873), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n966), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n970), .A2(G953), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n321), .A2(new_n325), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(new_n526), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n801), .B1(new_n778), .B2(new_n791), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n787), .A2(new_n363), .A3(new_n735), .A4(new_n708), .ZN(new_n976));
  INV_X1    g790(.A(new_n769), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n976), .A2(new_n763), .A3(new_n977), .A4(new_n873), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n975), .A2(G953), .A3(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n973), .B1(new_n678), .B2(new_n214), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n964), .B1(new_n974), .B2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n964), .ZN(new_n983));
  OAI221_X1 g797(.A(new_n983), .B1(new_n979), .B2(new_n980), .C1(new_n971), .C2(new_n973), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n982), .A2(new_n984), .ZN(G72));
  NOR2_X1   g799(.A1(new_n348), .A2(new_n311), .ZN(new_n986));
  NOR4_X1   g800(.A1(new_n975), .A2(new_n860), .A3(new_n978), .A4(new_n870), .ZN(new_n987));
  NAND2_X1  g801(.A1(G472), .A2(G902), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT63), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n986), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n989), .B1(new_n970), .B2(new_n887), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n348), .A2(new_n311), .ZN(new_n992));
  OAI211_X1 g806(.A(new_n990), .B(new_n945), .C1(new_n991), .C2(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n886), .B1(new_n891), .B2(new_n894), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n348), .A2(new_n349), .ZN(new_n995));
  AOI211_X1 g809(.A(new_n989), .B(new_n994), .C1(new_n702), .C2(new_n995), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n993), .A2(new_n996), .ZN(G57));
endmodule


