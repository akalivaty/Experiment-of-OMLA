//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 0 0 0 0 0 0 1 1 0 0 1 0 0 1 0 0 1 1 1 0 1 0 1 1 1 0 1 0 1 1 1 1 1 1 1 0 0 0 1 1 1 1 0 1 1 1 1 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n530, new_n531, new_n532, new_n533, new_n534, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n544, new_n545,
    new_n546, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n567, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n598, new_n599, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1156, new_n1157;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  XNOR2_X1  g042(.A(new_n467), .B(KEYINPUT67), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n460), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g044(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G137), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n462), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n469), .A2(new_n474), .ZN(G160));
  NAND2_X1  g050(.A1(new_n470), .A2(G136), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n476), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  AND2_X1   g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NOR2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  OAI211_X1 g059(.A(G138), .B(new_n460), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT4), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n465), .A2(new_n487), .A3(G138), .A4(new_n460), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n460), .A2(G114), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n494), .A2(new_n496), .A3(KEYINPUT68), .A4(G2104), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n493), .A2(new_n497), .B1(new_n477), .B2(G126), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n489), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  XNOR2_X1  g075(.A(KEYINPUT5), .B(G543), .ZN(new_n501));
  NOR2_X1   g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  AND2_X1   g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G88), .ZN(new_n505));
  INV_X1    g080(.A(G50), .ZN(new_n506));
  OAI21_X1  g081(.A(G543), .B1(new_n503), .B2(new_n502), .ZN(new_n507));
  OAI22_X1  g082(.A1(new_n504), .A2(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n501), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OR2_X1    g086(.A1(new_n508), .A2(new_n511), .ZN(G303));
  INV_X1    g087(.A(G303), .ZN(G166));
  XOR2_X1   g088(.A(KEYINPUT5), .B(G543), .Z(new_n514));
  NOR2_X1   g089(.A1(new_n503), .A2(new_n502), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G89), .ZN(new_n517));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n518), .B(KEYINPUT7), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT70), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n517), .A2(KEYINPUT70), .A3(new_n519), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n514), .A2(new_n510), .ZN(new_n524));
  INV_X1    g099(.A(new_n507), .ZN(new_n525));
  XOR2_X1   g100(.A(KEYINPUT69), .B(G51), .Z(new_n526));
  AOI22_X1  g101(.A1(new_n524), .A2(G63), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n522), .A2(new_n523), .A3(new_n527), .ZN(G286));
  INV_X1    g103(.A(G286), .ZN(G168));
  XNOR2_X1  g104(.A(KEYINPUT72), .B(G90), .ZN(new_n530));
  XOR2_X1   g105(.A(KEYINPUT71), .B(G52), .Z(new_n531));
  OAI22_X1  g106(.A1(new_n504), .A2(new_n530), .B1(new_n507), .B2(new_n531), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n501), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n510), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n532), .A2(new_n534), .ZN(G171));
  INV_X1    g110(.A(G81), .ZN(new_n536));
  INV_X1    g111(.A(G43), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n504), .A2(new_n536), .B1(new_n537), .B2(new_n507), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n501), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n510), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  NAND4_X1  g117(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g118(.A(KEYINPUT73), .B(KEYINPUT8), .Z(new_n544));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n544), .B(new_n545), .ZN(new_n546));
  NAND4_X1  g121(.A1(G319), .A2(G483), .A3(G661), .A4(new_n546), .ZN(G188));
  INV_X1    g122(.A(KEYINPUT9), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT74), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G53), .ZN(new_n550));
  OR3_X1    g125(.A1(new_n507), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n548), .B1(new_n507), .B2(new_n550), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(KEYINPUT75), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT75), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n551), .A2(new_n555), .A3(new_n552), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n514), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G651), .ZN(new_n561));
  INV_X1    g136(.A(G91), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n562), .B2(new_n504), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n557), .A2(new_n564), .ZN(G299));
  INV_X1    g140(.A(G171), .ZN(G301));
  AOI22_X1  g141(.A1(new_n516), .A2(G87), .B1(new_n525), .B2(G49), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n501), .B2(G74), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n568), .A2(KEYINPUT76), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(KEYINPUT76), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n567), .A2(new_n569), .A3(new_n570), .ZN(G288));
  AOI22_X1  g146(.A1(new_n501), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n572), .A2(new_n510), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n516), .A2(G86), .B1(new_n525), .B2(G48), .ZN(new_n574));
  AND2_X1   g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G305));
  NAND2_X1  g151(.A1(G72), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G60), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n514), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n510), .B1(new_n579), .B2(KEYINPUT77), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n580), .B1(KEYINPUT77), .B2(new_n579), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n516), .A2(G85), .B1(new_n525), .B2(G47), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G290));
  NAND3_X1  g158(.A1(new_n516), .A2(KEYINPUT10), .A3(G92), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT10), .ZN(new_n585));
  INV_X1    g160(.A(G92), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n504), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(G79), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G66), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n514), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n591), .A2(G651), .B1(new_n525), .B2(G54), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(G868), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n595), .B1(new_n594), .B2(G171), .ZN(G284));
  OAI21_X1  g171(.A(new_n595), .B1(new_n594), .B2(G171), .ZN(G321));
  NAND2_X1  g172(.A1(G286), .A2(G868), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n563), .B1(new_n554), .B2(new_n556), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(G868), .B2(new_n599), .ZN(G297));
  OAI21_X1  g175(.A(new_n598), .B1(G868), .B2(new_n599), .ZN(G280));
  INV_X1    g176(.A(new_n593), .ZN(new_n602));
  INV_X1    g177(.A(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(G860), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT78), .ZN(G148));
  OAI21_X1  g180(.A(KEYINPUT79), .B1(new_n541), .B2(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n602), .A2(new_n603), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G868), .ZN(new_n608));
  MUX2_X1   g183(.A(KEYINPUT79), .B(new_n606), .S(new_n608), .Z(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g185(.A1(new_n465), .A2(new_n472), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT12), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT13), .ZN(new_n613));
  INV_X1    g188(.A(G2100), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n613), .A2(new_n614), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n470), .A2(G135), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n477), .A2(G123), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n460), .A2(G111), .ZN(new_n619));
  OAI21_X1  g194(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n617), .B(new_n618), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(G2096), .Z(new_n622));
  NAND3_X1  g197(.A1(new_n615), .A2(new_n616), .A3(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT80), .Z(G156));
  XOR2_X1   g199(.A(KEYINPUT15), .B(G2435), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2438), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2427), .B(G2430), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT81), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n626), .A2(new_n628), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n629), .A2(KEYINPUT14), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2443), .B(G2446), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G1341), .B(G1348), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(G2451), .B(G2454), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT82), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n635), .A2(new_n639), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(G14), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT83), .ZN(G401));
  XOR2_X1   g218(.A(G2084), .B(G2090), .Z(new_n644));
  XNOR2_X1  g219(.A(G2067), .B(G2678), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2072), .B(G2078), .Z(new_n647));
  NOR2_X1   g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT18), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n647), .B(KEYINPUT17), .ZN(new_n650));
  INV_X1    g225(.A(new_n644), .ZN(new_n651));
  INV_X1    g226(.A(new_n645), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n651), .A2(new_n647), .A3(new_n652), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n654), .A2(new_n646), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n649), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2096), .B(G2100), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(G227));
  XOR2_X1   g233(.A(G1971), .B(G1976), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  XOR2_X1   g235(.A(G1956), .B(G2474), .Z(new_n661));
  XOR2_X1   g236(.A(G1961), .B(G1966), .Z(new_n662));
  AND2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT20), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n661), .A2(new_n662), .ZN(new_n666));
  NOR3_X1   g241(.A1(new_n660), .A2(new_n663), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n667), .B1(new_n660), .B2(new_n666), .ZN(new_n668));
  AND2_X1   g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1991), .B(G1996), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1981), .B(G1986), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(G229));
  INV_X1    g250(.A(G16), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(G23), .ZN(new_n677));
  INV_X1    g252(.A(G288), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n677), .B1(new_n678), .B2(new_n676), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT33), .ZN(new_n680));
  INV_X1    g255(.A(G1976), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n676), .A2(G6), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n683), .B1(new_n575), .B2(new_n676), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT32), .B(G1981), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT87), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n684), .B(new_n686), .Z(new_n687));
  NAND2_X1  g262(.A1(new_n676), .A2(G22), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(G166), .B2(new_n676), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G1971), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n680), .A2(new_n681), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n682), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(KEYINPUT34), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT34), .ZN(new_n695));
  NAND4_X1  g270(.A1(new_n682), .A2(new_n691), .A3(new_n695), .A4(new_n692), .ZN(new_n696));
  INV_X1    g271(.A(G29), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G25), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n470), .A2(G131), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n477), .A2(G119), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n460), .A2(G107), .ZN(new_n701));
  OAI21_X1  g276(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n699), .B(new_n700), .C1(new_n701), .C2(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT84), .Z(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n698), .B1(new_n705), .B2(new_n697), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT35), .B(G1991), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT85), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n706), .B(new_n708), .ZN(new_n709));
  MUX2_X1   g284(.A(G24), .B(G290), .S(G16), .Z(new_n710));
  XOR2_X1   g285(.A(KEYINPUT86), .B(G1986), .Z(new_n711));
  XOR2_X1   g286(.A(new_n710), .B(new_n711), .Z(new_n712));
  NAND4_X1  g287(.A1(new_n694), .A2(new_n696), .A3(new_n709), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT36), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT98), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n676), .A2(G21), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G168), .B2(new_n676), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n717), .A2(KEYINPUT94), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n717), .A2(KEYINPUT94), .ZN(new_n719));
  OR3_X1    g294(.A1(new_n718), .A2(new_n719), .A3(G1966), .ZN(new_n720));
  OAI21_X1  g295(.A(G1966), .B1(new_n718), .B2(new_n719), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT30), .B(G28), .ZN(new_n722));
  OR2_X1    g297(.A1(KEYINPUT31), .A2(G11), .ZN(new_n723));
  NAND2_X1  g298(.A1(KEYINPUT31), .A2(G11), .ZN(new_n724));
  AOI22_X1  g299(.A1(new_n722), .A2(new_n697), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(new_n621), .B2(new_n697), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n676), .A2(G5), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G171), .B2(new_n676), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n726), .B1(new_n728), .B2(G1961), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n720), .A2(new_n721), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT95), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT27), .B(G1996), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n470), .A2(G141), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT91), .Z(new_n734));
  AND2_X1   g309(.A1(new_n472), .A2(G105), .ZN(new_n735));
  NAND3_X1  g310(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT26), .ZN(new_n737));
  AOI211_X1 g312(.A(new_n735), .B(new_n737), .C1(G129), .C2(new_n477), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT92), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n740), .A2(new_n697), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(KEYINPUT93), .ZN(new_n742));
  INV_X1    g317(.A(G32), .ZN(new_n743));
  AOI21_X1  g318(.A(KEYINPUT93), .B1(new_n697), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n740), .B2(new_n697), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n732), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  AND2_X1   g321(.A1(KEYINPUT24), .A2(G34), .ZN(new_n747));
  NOR2_X1   g322(.A1(KEYINPUT24), .A2(G34), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n697), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT90), .Z(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G160), .B2(G29), .ZN(new_n751));
  OAI22_X1  g326(.A1(new_n728), .A2(G1961), .B1(new_n751), .B2(G2084), .ZN(new_n752));
  OR3_X1    g327(.A1(new_n746), .A2(KEYINPUT96), .A3(new_n752), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT97), .B(KEYINPUT23), .Z(new_n754));
  NAND2_X1  g329(.A1(new_n676), .A2(G20), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n599), .B2(new_n676), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G1956), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n742), .A2(new_n745), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n758), .B1(new_n759), .B2(new_n732), .ZN(new_n760));
  OAI21_X1  g335(.A(KEYINPUT96), .B1(new_n746), .B2(new_n752), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n697), .A2(G33), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT25), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n465), .A2(G127), .ZN(new_n765));
  NAND2_X1  g340(.A1(G115), .A2(G2104), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n460), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AOI211_X1 g342(.A(new_n764), .B(new_n767), .C1(G139), .C2(new_n470), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n762), .B1(new_n768), .B2(new_n697), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n769), .A2(G2072), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G2084), .B2(new_n751), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n676), .A2(G4), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n602), .B2(new_n676), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n773), .A2(G1348), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(G1348), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n771), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n697), .A2(G27), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G164), .B2(new_n697), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(G2078), .Z(new_n779));
  NAND2_X1  g354(.A1(new_n541), .A2(G16), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G16), .B2(G19), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT88), .B(G1341), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n781), .A2(new_n783), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n769), .A2(G2072), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n779), .A2(new_n784), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n470), .A2(G140), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n477), .A2(G128), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n460), .A2(G116), .ZN(new_n790));
  OAI21_X1  g365(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n788), .B(new_n789), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(G29), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT89), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n697), .A2(G26), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT28), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G2067), .ZN(new_n798));
  NOR2_X1   g373(.A1(G29), .A2(G35), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G162), .B2(G29), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT29), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G2090), .ZN(new_n802));
  NOR4_X1   g377(.A1(new_n776), .A2(new_n787), .A3(new_n798), .A4(new_n802), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n753), .A2(new_n760), .A3(new_n761), .A4(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n731), .A2(new_n804), .ZN(new_n805));
  AND3_X1   g380(.A1(new_n714), .A2(new_n715), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n715), .B1(new_n714), .B2(new_n805), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n806), .A2(new_n807), .ZN(G311));
  NAND2_X1  g383(.A1(new_n714), .A2(new_n805), .ZN(G150));
  NAND2_X1  g384(.A1(new_n516), .A2(G93), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n525), .A2(G55), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(KEYINPUT99), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT99), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n810), .A2(new_n814), .A3(new_n811), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n501), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n817), .A2(new_n510), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(G860), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT37), .Z(new_n821));
  NAND2_X1  g396(.A1(new_n602), .A2(G559), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT38), .ZN(new_n823));
  INV_X1    g398(.A(new_n541), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n819), .A2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n815), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n814), .B1(new_n810), .B2(new_n811), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n541), .B(new_n818), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n823), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n823), .A2(new_n829), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n830), .A2(KEYINPUT39), .A3(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT100), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT101), .ZN(new_n834));
  AOI21_X1  g409(.A(KEYINPUT39), .B1(new_n830), .B2(new_n831), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n835), .A2(G860), .ZN(new_n836));
  AND3_X1   g411(.A1(new_n833), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n834), .B1(new_n833), .B2(new_n836), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n821), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT102), .ZN(G145));
  XOR2_X1   g415(.A(new_n792), .B(KEYINPUT104), .Z(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n703), .B(KEYINPUT106), .Z(new_n843));
  INV_X1    g418(.A(new_n612), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n843), .A2(new_n844), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n470), .A2(G142), .ZN(new_n847));
  INV_X1    g422(.A(new_n477), .ZN(new_n848));
  INV_X1    g423(.A(G130), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n460), .A2(G118), .ZN(new_n850));
  OAI21_X1  g425(.A(KEYINPUT105), .B1(G106), .B2(G2105), .ZN(new_n851));
  AND2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT105), .ZN(new_n853));
  OAI21_X1  g428(.A(G2104), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  OAI221_X1 g429(.A(new_n847), .B1(new_n848), .B2(new_n849), .C1(new_n852), .C2(new_n854), .ZN(new_n855));
  OR3_X1    g430(.A1(new_n845), .A2(new_n846), .A3(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n855), .B1(new_n845), .B2(new_n846), .ZN(new_n857));
  AND3_X1   g432(.A1(new_n856), .A2(new_n499), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n499), .B1(new_n856), .B2(new_n857), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n842), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n856), .A2(new_n857), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(G164), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n856), .A2(new_n499), .A3(new_n857), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n862), .A2(new_n841), .A3(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n739), .A2(new_n768), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n865), .B1(new_n740), .B2(new_n768), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n860), .A2(new_n864), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n867), .B1(new_n860), .B2(new_n864), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XOR2_X1   g445(.A(G160), .B(KEYINPUT103), .Z(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(G162), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n621), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(G37), .B1(new_n870), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n860), .A2(new_n864), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(new_n866), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n860), .A2(new_n864), .A3(new_n867), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n874), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n875), .A2(KEYINPUT40), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT40), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n877), .A2(new_n874), .A3(new_n878), .ZN(new_n883));
  INV_X1    g458(.A(G37), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n882), .B1(new_n885), .B2(new_n879), .ZN(new_n886));
  AND2_X1   g461(.A1(new_n881), .A2(new_n886), .ZN(G395));
  NAND2_X1  g462(.A1(new_n819), .A2(new_n594), .ZN(new_n888));
  XOR2_X1   g463(.A(G303), .B(KEYINPUT108), .Z(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(G288), .ZN(new_n890));
  XNOR2_X1  g465(.A(G290), .B(G305), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n889), .B(new_n678), .ZN(new_n893));
  INV_X1    g468(.A(new_n891), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(KEYINPUT42), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n829), .B(new_n607), .Z(new_n898));
  NAND2_X1  g473(.A1(G299), .A2(new_n602), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT107), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n599), .A2(new_n900), .A3(new_n593), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n900), .B1(new_n599), .B2(new_n593), .ZN(new_n903));
  OAI21_X1  g478(.A(KEYINPUT41), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n903), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT41), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n905), .A2(new_n906), .A3(new_n899), .A4(new_n901), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n898), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n902), .A2(new_n903), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n910), .B1(new_n898), .B2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n897), .B(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n888), .B1(new_n913), .B2(new_n594), .ZN(G295));
  OAI21_X1  g489(.A(new_n888), .B1(new_n913), .B2(new_n594), .ZN(G331));
  AND2_X1   g490(.A1(new_n892), .A2(new_n895), .ZN(new_n916));
  OAI21_X1  g491(.A(KEYINPUT109), .B1(new_n532), .B2(new_n534), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT110), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n523), .A2(new_n527), .ZN(new_n919));
  AOI21_X1  g494(.A(KEYINPUT70), .B1(new_n517), .B2(new_n519), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n917), .B(new_n918), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n918), .B1(G286), .B2(new_n917), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n825), .B(new_n828), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n917), .B1(new_n919), .B2(new_n920), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(KEYINPUT110), .ZN(new_n926));
  INV_X1    g501(.A(new_n828), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n541), .B1(new_n816), .B2(new_n818), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n926), .B(new_n921), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(G301), .A2(KEYINPUT109), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n924), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n930), .B1(new_n924), .B2(new_n929), .ZN(new_n933));
  NOR3_X1   g508(.A1(new_n932), .A2(new_n933), .A3(new_n911), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n924), .A2(new_n929), .ZN(new_n935));
  INV_X1    g510(.A(new_n930), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n908), .B1(new_n937), .B2(new_n931), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n916), .B1(new_n934), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n909), .B1(new_n932), .B2(new_n933), .ZN(new_n940));
  INV_X1    g515(.A(new_n911), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n937), .A2(new_n941), .A3(new_n931), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n940), .A2(new_n896), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n939), .A2(new_n884), .A3(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n944), .A2(KEYINPUT43), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n944), .A2(KEYINPUT43), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n946), .A2(KEYINPUT44), .A3(new_n947), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n944), .A2(KEYINPUT111), .A3(KEYINPUT43), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT111), .B1(new_n944), .B2(KEYINPUT43), .ZN(new_n950));
  NOR3_X1   g525(.A1(new_n949), .A2(new_n950), .A3(new_n945), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n948), .B1(new_n951), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g527(.A(G1384), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n499), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT45), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n466), .A2(new_n468), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(G2105), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n958), .A2(G40), .A3(new_n473), .A4(new_n471), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n792), .B(G2067), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n960), .B1(new_n739), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n960), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n963), .A2(G1996), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n962), .B1(new_n964), .B2(KEYINPUT46), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n965), .B1(KEYINPUT46), .B2(new_n964), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n966), .B(KEYINPUT47), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n961), .B1(G1996), .B2(new_n739), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n968), .B1(new_n740), .B2(G1996), .ZN(new_n969));
  XOR2_X1   g544(.A(new_n703), .B(new_n707), .Z(new_n970));
  OAI21_X1  g545(.A(new_n960), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(G290), .A2(G1986), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n960), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n973), .B(KEYINPUT48), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n967), .B1(new_n971), .B2(new_n974), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n969), .A2(new_n960), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n705), .A2(new_n707), .ZN(new_n977));
  OAI22_X1  g552(.A1(new_n976), .A2(new_n977), .B1(G2067), .B2(new_n792), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT125), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n963), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n980), .B1(new_n979), .B2(new_n978), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n975), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n954), .A2(KEYINPUT50), .ZN(new_n983));
  INV_X1    g558(.A(G2084), .ZN(new_n984));
  INV_X1    g559(.A(G40), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n469), .A2(new_n474), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(G1384), .B1(new_n489), .B2(new_n498), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT50), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n983), .A2(new_n984), .A3(new_n986), .A4(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT119), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n959), .B1(new_n954), .B2(KEYINPUT50), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n993), .A2(KEYINPUT119), .A3(new_n984), .A4(new_n989), .ZN(new_n994));
  INV_X1    g569(.A(G1966), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n955), .A2(G1384), .ZN(new_n996));
  AND2_X1   g571(.A1(new_n486), .A2(new_n488), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n493), .A2(new_n497), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n477), .A2(G126), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n996), .B1(new_n997), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n986), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT45), .B1(new_n499), .B2(new_n953), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n995), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n992), .A2(G168), .A3(new_n994), .A4(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(G8), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT51), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1007), .A2(KEYINPUT123), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(KEYINPUT123), .B(KEYINPUT51), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1005), .A2(G8), .A3(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n992), .A2(new_n994), .A3(new_n1004), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1012), .A2(G8), .A3(G286), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1009), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT62), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1009), .A2(KEYINPUT62), .A3(new_n1011), .A4(new_n1013), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n986), .A2(new_n987), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(G8), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT116), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT116), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  AOI22_X1  g599(.A1(new_n1022), .A2(new_n1024), .B1(G1976), .B2(new_n678), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT52), .B1(G288), .B2(new_n681), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  XOR2_X1   g602(.A(KEYINPUT117), .B(G1981), .Z(new_n1028));
  NAND2_X1  g603(.A1(new_n575), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G1981), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1029), .B1(new_n1030), .B2(new_n575), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT49), .ZN(new_n1032));
  OR2_X1    g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1022), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1024), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1033), .B(new_n1034), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1027), .B(new_n1037), .C1(new_n1038), .C2(new_n1025), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT113), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1001), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n499), .A2(KEYINPUT113), .A3(new_n996), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n956), .A2(new_n1041), .A3(new_n986), .A4(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT114), .ZN(new_n1044));
  INV_X1    g619(.A(G1971), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT113), .B1(new_n499), .B2(new_n996), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1003), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1047), .A2(new_n1048), .A3(new_n986), .A4(new_n1042), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1044), .A2(new_n1045), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n993), .A2(new_n989), .ZN(new_n1051));
  OR2_X1    g626(.A1(new_n1051), .A2(G2090), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n1050), .A2(KEYINPUT115), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT115), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1054));
  INV_X1    g629(.A(G8), .ZN(new_n1055));
  NOR3_X1   g630(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(G303), .A2(G8), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n1057), .B(KEYINPUT55), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1039), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(G8), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1062), .A2(new_n1063), .A3(new_n1058), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1055), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1065));
  OAI21_X1  g640(.A(KEYINPUT118), .B1(new_n1065), .B2(new_n1059), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n1068));
  OR4_X1    g643(.A1(new_n1068), .A2(new_n1002), .A3(G2078), .A4(new_n1003), .ZN(new_n1069));
  INV_X1    g644(.A(G1961), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1051), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(G2078), .B1(new_n1044), .B2(new_n1049), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1069), .B(new_n1071), .C1(new_n1072), .C2(KEYINPUT53), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n1073), .A2(G171), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1018), .A2(new_n1060), .A3(new_n1067), .A4(new_n1074), .ZN(new_n1075));
  XOR2_X1   g650(.A(G171), .B(KEYINPUT54), .Z(new_n1076));
  NAND2_X1  g651(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n1047), .A2(new_n1042), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1068), .A2(new_n985), .A3(G2078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT124), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n958), .B(new_n1079), .C1(new_n474), .C2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1081), .B1(new_n1080), .B2(new_n474), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1076), .B1(new_n1078), .B2(new_n1082), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1071), .B(new_n1083), .C1(new_n1072), .C2(KEYINPUT53), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1014), .A2(new_n1077), .A3(new_n1084), .ZN(new_n1085));
  NOR3_X1   g660(.A1(new_n563), .A2(KEYINPUT57), .A3(new_n553), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1086), .B1(G299), .B2(KEYINPUT57), .ZN(new_n1087));
  XOR2_X1   g662(.A(KEYINPUT56), .B(G2072), .Z(new_n1088));
  OR2_X1    g663(.A1(new_n1043), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G1956), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1051), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1087), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1091), .B(new_n1087), .C1(new_n1043), .C2(new_n1088), .ZN(new_n1093));
  INV_X1    g668(.A(G1348), .ZN(new_n1094));
  INV_X1    g669(.A(new_n989), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1094), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  OR2_X1    g672(.A1(new_n1019), .A2(G2067), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n593), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1092), .B1(new_n1093), .B2(new_n1099), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n1097), .A2(new_n593), .A3(new_n1098), .ZN(new_n1101));
  OAI21_X1  g676(.A(KEYINPUT60), .B1(new_n1101), .B2(new_n1099), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n593), .A2(KEYINPUT60), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1097), .A2(new_n1098), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1019), .ZN(new_n1105));
  XNOR2_X1  g680(.A(KEYINPUT58), .B(G1341), .ZN(new_n1106));
  OAI22_X1  g681(.A1(new_n1043), .A2(G1996), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT59), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n824), .A2(KEYINPUT121), .ZN(new_n1109));
  AND3_X1   g684(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1108), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1102), .B(new_n1104), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1112));
  AND2_X1   g687(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n1093), .B(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1100), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1085), .A2(new_n1060), .A3(new_n1067), .A4(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT115), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1061), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1050), .A2(KEYINPUT115), .A3(new_n1052), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1118), .A2(G8), .A3(new_n1059), .A4(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1120), .A2(new_n1039), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1037), .A2(new_n681), .A3(new_n678), .ZN(new_n1122));
  AOI22_X1  g697(.A1(new_n1122), .A2(new_n1029), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1075), .A2(new_n1116), .A3(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1027), .A2(new_n1037), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1025), .A2(new_n1038), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n1120), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1059), .B1(new_n1130), .B2(new_n1119), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1012), .A2(G8), .A3(G168), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT63), .ZN(new_n1133));
  OR2_X1    g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n1129), .A2(new_n1131), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1063), .B1(new_n1062), .B2(new_n1058), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1065), .A2(KEYINPUT118), .A3(new_n1059), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1128), .B(new_n1120), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1133), .B1(new_n1138), .B2(new_n1132), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT120), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1135), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  OAI211_X1 g716(.A(KEYINPUT120), .B(new_n1133), .C1(new_n1138), .C2(new_n1132), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1125), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  AND2_X1   g718(.A1(G290), .A2(G1986), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n960), .B1(new_n1144), .B2(new_n972), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1145), .B(KEYINPUT112), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n971), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n982), .B1(new_n1143), .B2(new_n1147), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g723(.A1(G227), .A2(new_n458), .ZN(new_n1150));
  AND3_X1   g724(.A1(new_n642), .A2(KEYINPUT126), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g725(.A(KEYINPUT126), .B1(new_n642), .B2(new_n1150), .ZN(new_n1152));
  NOR3_X1   g726(.A1(new_n1151), .A2(G229), .A3(new_n1152), .ZN(new_n1153));
  OAI21_X1  g727(.A(new_n1153), .B1(new_n885), .B2(new_n879), .ZN(new_n1154));
  NOR2_X1   g728(.A1(new_n951), .A2(new_n1154), .ZN(G308));
  NAND2_X1  g729(.A1(new_n875), .A2(new_n880), .ZN(new_n1156));
  OR2_X1    g730(.A1(new_n950), .A2(new_n945), .ZN(new_n1157));
  OAI211_X1 g731(.A(new_n1156), .B(new_n1153), .C1(new_n1157), .C2(new_n949), .ZN(G225));
endmodule


