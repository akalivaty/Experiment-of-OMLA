//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 1 1 0 1 0 1 1 1 0 0 0 1 0 0 0 1 0 0 0 1 0 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:56 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1081, new_n1082, new_n1083, new_n1084, new_n1085,
    new_n1086, new_n1087, new_n1088, new_n1089, new_n1090, new_n1091,
    new_n1092, new_n1093, new_n1094, new_n1095, new_n1096, new_n1097,
    new_n1098, new_n1099, new_n1100, new_n1101, new_n1102, new_n1103,
    new_n1104, new_n1105, new_n1106, new_n1107, new_n1108, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186;
  NOR2_X1   g000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g001(.A(G50), .ZN(new_n202));
  NAND2_X1  g002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g006(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n207));
  XOR2_X1   g007(.A(new_n207), .B(KEYINPUT64), .Z(new_n208));
  AOI22_X1  g008(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n209));
  AOI22_X1  g009(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n210));
  NAND2_X1  g010(.A1(G68), .A2(G238), .ZN(new_n211));
  NAND4_X1  g011(.A1(new_n208), .A2(new_n209), .A3(new_n210), .A4(new_n211), .ZN(new_n212));
  INV_X1    g012(.A(G226), .ZN(new_n213));
  NOR2_X1   g013(.A1(new_n202), .A2(new_n213), .ZN(new_n214));
  OAI21_X1  g014(.A(new_n206), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g015(.A(new_n215), .B(KEYINPUT1), .ZN(new_n216));
  OAI21_X1  g016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  INV_X1    g017(.A(G20), .ZN(new_n218));
  NAND2_X1  g018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR3_X1   g019(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NOR2_X1   g020(.A1(new_n206), .A2(G13), .ZN(new_n221));
  OAI211_X1 g021(.A(new_n221), .B(G250), .C1(G257), .C2(G264), .ZN(new_n222));
  XOR2_X1   g022(.A(new_n222), .B(KEYINPUT0), .Z(new_n223));
  NOR3_X1   g023(.A1(new_n216), .A2(new_n220), .A3(new_n223), .ZN(G361));
  XNOR2_X1  g024(.A(G238), .B(G244), .ZN(new_n225));
  INV_X1    g025(.A(G232), .ZN(new_n226));
  XNOR2_X1  g026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g027(.A(new_n227), .B(KEYINPUT2), .ZN(new_n228));
  XNOR2_X1  g028(.A(new_n228), .B(new_n213), .ZN(new_n229));
  XNOR2_X1  g029(.A(G250), .B(G257), .ZN(new_n230));
  INV_X1    g030(.A(G264), .ZN(new_n231));
  XNOR2_X1  g031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g032(.A(new_n232), .B(G270), .ZN(new_n233));
  XNOR2_X1  g033(.A(new_n229), .B(new_n233), .ZN(G358));
  XNOR2_X1  g034(.A(G50), .B(G68), .ZN(new_n235));
  XNOR2_X1  g035(.A(new_n235), .B(G58), .ZN(new_n236));
  XNOR2_X1  g036(.A(new_n236), .B(G77), .ZN(new_n237));
  XNOR2_X1  g037(.A(G97), .B(G107), .ZN(new_n238));
  XNOR2_X1  g038(.A(new_n238), .B(G87), .ZN(new_n239));
  INV_X1    g039(.A(G116), .ZN(new_n240));
  XNOR2_X1  g040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g041(.A(new_n237), .B(new_n241), .Z(G351));
  INV_X1    g042(.A(G33), .ZN(new_n243));
  AND3_X1   g043(.A1(new_n243), .A2(KEYINPUT70), .A3(KEYINPUT3), .ZN(new_n244));
  XNOR2_X1  g044(.A(KEYINPUT3), .B(G33), .ZN(new_n245));
  INV_X1    g045(.A(KEYINPUT70), .ZN(new_n246));
  AOI21_X1  g046(.A(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g047(.A(KEYINPUT7), .ZN(new_n248));
  NAND2_X1  g048(.A1(new_n248), .A2(KEYINPUT71), .ZN(new_n249));
  NOR2_X1   g049(.A1(new_n248), .A2(KEYINPUT71), .ZN(new_n250));
  INV_X1    g050(.A(new_n250), .ZN(new_n251));
  NAND4_X1  g051(.A1(new_n247), .A2(new_n218), .A3(new_n249), .A4(new_n251), .ZN(new_n252));
  NAND2_X1  g052(.A1(new_n243), .A2(KEYINPUT3), .ZN(new_n253));
  INV_X1    g053(.A(KEYINPUT3), .ZN(new_n254));
  NAND2_X1  g054(.A1(new_n254), .A2(G33), .ZN(new_n255));
  NAND3_X1  g055(.A1(new_n253), .A2(new_n255), .A3(new_n246), .ZN(new_n256));
  NAND3_X1  g056(.A1(new_n243), .A2(KEYINPUT70), .A3(KEYINPUT3), .ZN(new_n257));
  NAND4_X1  g057(.A1(new_n256), .A2(new_n218), .A3(new_n257), .A4(new_n249), .ZN(new_n258));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n250), .ZN(new_n259));
  NAND3_X1  g059(.A1(new_n252), .A2(new_n259), .A3(G68), .ZN(new_n260));
  INV_X1    g060(.A(G58), .ZN(new_n261));
  INV_X1    g061(.A(G68), .ZN(new_n262));
  NOR2_X1   g062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OR2_X1    g063(.A1(new_n263), .A2(new_n201), .ZN(new_n264));
  NOR2_X1   g064(.A1(G20), .A2(G33), .ZN(new_n265));
  AOI22_X1  g065(.A1(new_n264), .A2(G20), .B1(G159), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g066(.A1(new_n260), .A2(KEYINPUT16), .A3(new_n266), .ZN(new_n267));
  OAI21_X1  g067(.A(KEYINPUT7), .B1(new_n245), .B2(G20), .ZN(new_n268));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n255), .ZN(new_n269));
  NAND3_X1  g069(.A1(new_n269), .A2(new_n248), .A3(new_n218), .ZN(new_n270));
  NAND2_X1  g070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g071(.A(new_n266), .B1(new_n271), .B2(new_n262), .ZN(new_n272));
  INV_X1    g072(.A(KEYINPUT16), .ZN(new_n273));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g074(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n275));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n219), .ZN(new_n276));
  NAND3_X1  g076(.A1(new_n267), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  INV_X1    g077(.A(G13), .ZN(new_n278));
  NOR3_X1   g078(.A1(new_n278), .A2(new_n218), .A3(G1), .ZN(new_n279));
  INV_X1    g079(.A(new_n279), .ZN(new_n280));
  XNOR2_X1  g080(.A(KEYINPUT8), .B(G58), .ZN(new_n281));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g082(.A(G1), .ZN(new_n283));
  AOI21_X1  g083(.A(new_n276), .B1(new_n283), .B2(G20), .ZN(new_n284));
  OAI21_X1  g084(.A(new_n282), .B1(new_n284), .B2(new_n281), .ZN(new_n285));
  NAND2_X1  g085(.A1(new_n277), .A2(new_n285), .ZN(new_n286));
  INV_X1    g086(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g087(.A(new_n219), .B1(G33), .B2(G41), .ZN(new_n288));
  INV_X1    g088(.A(G41), .ZN(new_n289));
  INV_X1    g089(.A(G45), .ZN(new_n290));
  AOI21_X1  g090(.A(G1), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NOR2_X1   g091(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  INV_X1    g092(.A(new_n292), .ZN(new_n293));
  OAI21_X1  g093(.A(KEYINPUT74), .B1(new_n293), .B2(new_n226), .ZN(new_n294));
  NAND3_X1  g094(.A1(new_n291), .A2(KEYINPUT65), .A3(G274), .ZN(new_n295));
  INV_X1    g095(.A(KEYINPUT65), .ZN(new_n296));
  OAI21_X1  g096(.A(new_n283), .B1(G41), .B2(G45), .ZN(new_n297));
  INV_X1    g097(.A(G274), .ZN(new_n298));
  OAI21_X1  g098(.A(new_n296), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g099(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  INV_X1    g100(.A(KEYINPUT74), .ZN(new_n301));
  NAND3_X1  g101(.A1(new_n292), .A2(new_n301), .A3(G232), .ZN(new_n302));
  NAND3_X1  g102(.A1(new_n294), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  INV_X1    g103(.A(new_n303), .ZN(new_n304));
  INV_X1    g104(.A(G190), .ZN(new_n305));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g106(.A1(new_n256), .A2(new_n257), .ZN(new_n307));
  NAND3_X1  g107(.A1(new_n307), .A2(G226), .A3(G1698), .ZN(new_n308));
  NAND2_X1  g108(.A1(new_n308), .A2(KEYINPUT72), .ZN(new_n309));
  INV_X1    g109(.A(G87), .ZN(new_n310));
  NOR2_X1   g110(.A1(new_n243), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g111(.A(G1698), .B1(new_n256), .B2(new_n257), .ZN(new_n312));
  AOI21_X1  g112(.A(new_n311), .B1(new_n312), .B2(G223), .ZN(new_n313));
  INV_X1    g113(.A(KEYINPUT72), .ZN(new_n314));
  NAND4_X1  g114(.A1(new_n307), .A2(new_n314), .A3(G226), .A4(G1698), .ZN(new_n315));
  NAND3_X1  g115(.A1(new_n309), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n288), .ZN(new_n317));
  INV_X1    g117(.A(KEYINPUT73), .ZN(new_n318));
  NAND2_X1  g118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g119(.A1(new_n316), .A2(KEYINPUT73), .A3(new_n288), .ZN(new_n320));
  AOI21_X1  g120(.A(new_n306), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g121(.A(G200), .B1(new_n317), .B2(new_n304), .ZN(new_n322));
  OAI21_X1  g122(.A(new_n287), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g123(.A1(new_n323), .A2(KEYINPUT17), .ZN(new_n324));
  NOR2_X1   g124(.A1(new_n303), .A2(G190), .ZN(new_n325));
  AND3_X1   g125(.A1(new_n316), .A2(KEYINPUT73), .A3(new_n288), .ZN(new_n326));
  AOI21_X1  g126(.A(KEYINPUT73), .B1(new_n316), .B2(new_n288), .ZN(new_n327));
  OAI21_X1  g127(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g128(.A1(new_n317), .A2(new_n304), .ZN(new_n329));
  INV_X1    g129(.A(G200), .ZN(new_n330));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g131(.A(new_n286), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  INV_X1    g132(.A(KEYINPUT17), .ZN(new_n333));
  NAND2_X1  g133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NOR2_X1   g134(.A1(new_n303), .A2(G179), .ZN(new_n335));
  OAI21_X1  g135(.A(new_n335), .B1(new_n326), .B2(new_n327), .ZN(new_n336));
  INV_X1    g136(.A(G169), .ZN(new_n337));
  NAND2_X1  g137(.A1(new_n329), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g138(.A1(new_n336), .A2(new_n286), .A3(new_n338), .ZN(new_n339));
  INV_X1    g139(.A(KEYINPUT18), .ZN(new_n340));
  NAND2_X1  g140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND4_X1  g141(.A1(new_n336), .A2(new_n286), .A3(new_n338), .A4(KEYINPUT18), .ZN(new_n342));
  AOI22_X1  g142(.A1(new_n324), .A2(new_n334), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NOR2_X1   g143(.A1(new_n269), .A2(G1698), .ZN(new_n344));
  AOI22_X1  g144(.A1(new_n344), .A2(G222), .B1(G77), .B2(new_n269), .ZN(new_n345));
  INV_X1    g145(.A(G223), .ZN(new_n346));
  NAND2_X1  g146(.A1(new_n245), .A2(G1698), .ZN(new_n347));
  OAI21_X1  g147(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n288), .ZN(new_n349));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n300), .ZN(new_n350));
  AOI21_X1  g150(.A(new_n350), .B1(G226), .B2(new_n292), .ZN(new_n351));
  NAND2_X1  g151(.A1(new_n351), .A2(G190), .ZN(new_n352));
  NAND2_X1  g152(.A1(new_n284), .A2(G50), .ZN(new_n353));
  NAND2_X1  g153(.A1(new_n218), .A2(G33), .ZN(new_n354));
  INV_X1    g154(.A(G150), .ZN(new_n355));
  INV_X1    g155(.A(new_n265), .ZN(new_n356));
  OAI22_X1  g156(.A1(new_n281), .A2(new_n354), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g157(.A(new_n357), .B1(G20), .B2(new_n203), .ZN(new_n358));
  INV_X1    g158(.A(new_n276), .ZN(new_n359));
  OAI221_X1 g159(.A(new_n353), .B1(G50), .B2(new_n280), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  INV_X1    g160(.A(KEYINPUT9), .ZN(new_n361));
  OAI21_X1  g161(.A(KEYINPUT67), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g162(.A(new_n362), .B1(new_n361), .B2(new_n360), .ZN(new_n363));
  OAI211_X1 g163(.A(new_n352), .B(new_n363), .C1(new_n330), .C2(new_n351), .ZN(new_n364));
  XNOR2_X1  g164(.A(new_n364), .B(KEYINPUT10), .ZN(new_n365));
  INV_X1    g165(.A(G179), .ZN(new_n366));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n366), .ZN(new_n367));
  OAI211_X1 g167(.A(new_n367), .B(new_n360), .C1(G169), .C2(new_n351), .ZN(new_n368));
  NAND2_X1  g168(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  INV_X1    g169(.A(G1698), .ZN(new_n370));
  NOR2_X1   g170(.A1(new_n269), .A2(new_n370), .ZN(new_n371));
  AOI22_X1  g171(.A1(G232), .A2(new_n344), .B1(new_n371), .B2(G238), .ZN(new_n372));
  XNOR2_X1  g172(.A(KEYINPUT66), .B(G107), .ZN(new_n373));
  OAI21_X1  g173(.A(new_n372), .B1(new_n245), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n288), .ZN(new_n375));
  NAND2_X1  g175(.A1(new_n292), .A2(G244), .ZN(new_n376));
  NAND3_X1  g176(.A1(new_n375), .A2(new_n300), .A3(new_n376), .ZN(new_n377));
  OR2_X1    g177(.A1(new_n377), .A2(G179), .ZN(new_n378));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n337), .ZN(new_n379));
  INV_X1    g179(.A(new_n281), .ZN(new_n380));
  AOI22_X1  g180(.A1(new_n380), .A2(new_n265), .B1(G20), .B2(G77), .ZN(new_n381));
  XOR2_X1   g181(.A(KEYINPUT15), .B(G87), .Z(new_n382));
  INV_X1    g182(.A(new_n382), .ZN(new_n383));
  OAI21_X1  g183(.A(new_n381), .B1(new_n354), .B2(new_n383), .ZN(new_n384));
  INV_X1    g184(.A(G77), .ZN(new_n385));
  AOI22_X1  g185(.A1(new_n384), .A2(new_n276), .B1(new_n385), .B2(new_n279), .ZN(new_n386));
  INV_X1    g186(.A(new_n284), .ZN(new_n387));
  OAI21_X1  g187(.A(new_n386), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g188(.A1(new_n378), .A2(new_n379), .A3(new_n388), .ZN(new_n389));
  INV_X1    g189(.A(new_n389), .ZN(new_n390));
  NOR2_X1   g190(.A1(new_n369), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g191(.A(new_n388), .B1(new_n377), .B2(G200), .ZN(new_n392));
  OAI21_X1  g192(.A(new_n392), .B1(new_n305), .B2(new_n377), .ZN(new_n393));
  XOR2_X1   g193(.A(new_n300), .B(KEYINPUT68), .Z(new_n394));
  NAND2_X1  g194(.A1(new_n344), .A2(G226), .ZN(new_n395));
  NAND2_X1  g195(.A1(G33), .A2(G97), .ZN(new_n396));
  OAI211_X1 g196(.A(new_n395), .B(new_n396), .C1(new_n226), .C2(new_n347), .ZN(new_n397));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n288), .ZN(new_n398));
  NAND2_X1  g198(.A1(new_n292), .A2(G238), .ZN(new_n399));
  NAND3_X1  g199(.A1(new_n394), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g200(.A1(new_n400), .A2(KEYINPUT13), .ZN(new_n401));
  INV_X1    g201(.A(KEYINPUT13), .ZN(new_n402));
  NAND4_X1  g202(.A1(new_n394), .A2(new_n398), .A3(new_n402), .A4(new_n399), .ZN(new_n403));
  NAND2_X1  g203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g204(.A1(new_n404), .A2(G169), .ZN(new_n405));
  NAND2_X1  g205(.A1(new_n405), .A2(KEYINPUT14), .ZN(new_n406));
  NAND3_X1  g206(.A1(new_n401), .A2(G179), .A3(new_n403), .ZN(new_n407));
  INV_X1    g207(.A(KEYINPUT14), .ZN(new_n408));
  NAND3_X1  g208(.A1(new_n404), .A2(new_n408), .A3(G169), .ZN(new_n409));
  NAND3_X1  g209(.A1(new_n406), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g210(.A1(new_n265), .A2(G50), .ZN(new_n411));
  OAI221_X1 g211(.A(new_n411), .B1(new_n218), .B2(G68), .C1(new_n385), .C2(new_n354), .ZN(new_n412));
  AND2_X1   g212(.A1(new_n412), .A2(new_n276), .ZN(new_n413));
  AOI22_X1  g213(.A1(new_n413), .A2(KEYINPUT11), .B1(G68), .B2(new_n284), .ZN(new_n414));
  NAND2_X1  g214(.A1(new_n279), .A2(new_n262), .ZN(new_n415));
  XNOR2_X1  g215(.A(new_n415), .B(KEYINPUT12), .ZN(new_n416));
  OAI211_X1 g216(.A(new_n414), .B(new_n416), .C1(KEYINPUT11), .C2(new_n413), .ZN(new_n417));
  XNOR2_X1  g217(.A(new_n417), .B(KEYINPUT69), .ZN(new_n418));
  NAND2_X1  g218(.A1(new_n410), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g219(.A(new_n418), .B1(G200), .B2(new_n404), .ZN(new_n420));
  OAI21_X1  g220(.A(new_n420), .B1(new_n305), .B2(new_n404), .ZN(new_n421));
  AND2_X1   g221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  AND4_X1   g222(.A1(new_n343), .A2(new_n391), .A3(new_n393), .A4(new_n422), .ZN(new_n423));
  NAND3_X1  g223(.A1(new_n245), .A2(new_n218), .A3(G87), .ZN(new_n424));
  INV_X1    g224(.A(KEYINPUT22), .ZN(new_n425));
  NAND2_X1  g225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g226(.A1(new_n373), .A2(G20), .ZN(new_n427));
  NAND2_X1  g227(.A1(new_n427), .A2(KEYINPUT23), .ZN(new_n428));
  OR3_X1    g228(.A1(new_n218), .A2(KEYINPUT23), .A3(G107), .ZN(new_n429));
  NAND3_X1  g229(.A1(new_n426), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  INV_X1    g230(.A(new_n430), .ZN(new_n431));
  INV_X1    g231(.A(KEYINPUT80), .ZN(new_n432));
  NAND3_X1  g232(.A1(new_n307), .A2(KEYINPUT22), .A3(G87), .ZN(new_n433));
  NOR2_X1   g233(.A1(new_n243), .A2(new_n240), .ZN(new_n434));
  INV_X1    g234(.A(new_n434), .ZN(new_n435));
  AND2_X1   g235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  OAI211_X1 g236(.A(new_n431), .B(new_n432), .C1(new_n436), .C2(G20), .ZN(new_n437));
  AOI21_X1  g237(.A(G20), .B1(new_n433), .B2(new_n435), .ZN(new_n438));
  OAI21_X1  g238(.A(KEYINPUT80), .B1(new_n438), .B2(new_n430), .ZN(new_n439));
  NAND3_X1  g239(.A1(new_n437), .A2(KEYINPUT24), .A3(new_n439), .ZN(new_n440));
  INV_X1    g240(.A(KEYINPUT24), .ZN(new_n441));
  OAI211_X1 g241(.A(KEYINPUT80), .B(new_n441), .C1(new_n438), .C2(new_n430), .ZN(new_n442));
  NAND3_X1  g242(.A1(new_n440), .A2(new_n442), .A3(new_n276), .ZN(new_n443));
  AOI211_X1 g243(.A(new_n276), .B(new_n279), .C1(new_n283), .C2(G33), .ZN(new_n444));
  NAND2_X1  g244(.A1(new_n444), .A2(G107), .ZN(new_n445));
  NOR2_X1   g245(.A1(new_n280), .A2(G107), .ZN(new_n446));
  XNOR2_X1  g246(.A(new_n446), .B(KEYINPUT25), .ZN(new_n447));
  NAND3_X1  g247(.A1(new_n443), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  OAI21_X1  g248(.A(new_n307), .B1(G250), .B2(G1698), .ZN(new_n449));
  NOR2_X1   g249(.A1(new_n370), .A2(G257), .ZN(new_n450));
  INV_X1    g250(.A(G294), .ZN(new_n451));
  OAI22_X1  g251(.A1(new_n449), .A2(new_n450), .B1(new_n243), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n288), .ZN(new_n453));
  INV_X1    g253(.A(new_n288), .ZN(new_n454));
  AND2_X1   g254(.A1(KEYINPUT5), .A2(G41), .ZN(new_n455));
  NOR2_X1   g255(.A1(KEYINPUT5), .A2(G41), .ZN(new_n456));
  OAI211_X1 g256(.A(new_n283), .B(G45), .C1(new_n455), .C2(new_n456), .ZN(new_n457));
  AND2_X1   g257(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g258(.A1(new_n458), .A2(G264), .ZN(new_n459));
  OR2_X1    g259(.A1(new_n457), .A2(new_n298), .ZN(new_n460));
  NAND3_X1  g260(.A1(new_n453), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NOR2_X1   g261(.A1(new_n461), .A2(G179), .ZN(new_n462));
  AOI21_X1  g262(.A(new_n462), .B1(new_n337), .B2(new_n461), .ZN(new_n463));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g264(.A1(new_n464), .A2(KEYINPUT81), .ZN(new_n465));
  INV_X1    g265(.A(KEYINPUT81), .ZN(new_n466));
  NAND3_X1  g266(.A1(new_n448), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g268(.A1(new_n231), .A2(G1698), .ZN(new_n469));
  OAI211_X1 g269(.A(new_n307), .B(new_n469), .C1(G257), .C2(G1698), .ZN(new_n470));
  INV_X1    g270(.A(G303), .ZN(new_n471));
  OAI21_X1  g271(.A(new_n470), .B1(new_n471), .B2(new_n245), .ZN(new_n472));
  INV_X1    g272(.A(KEYINPUT79), .ZN(new_n473));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g274(.A(new_n470), .B(KEYINPUT79), .C1(new_n471), .C2(new_n245), .ZN(new_n475));
  NAND3_X1  g275(.A1(new_n474), .A2(new_n288), .A3(new_n475), .ZN(new_n476));
  INV_X1    g276(.A(new_n460), .ZN(new_n477));
  AOI21_X1  g277(.A(new_n477), .B1(G270), .B2(new_n458), .ZN(new_n478));
  NAND2_X1  g278(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g279(.A1(new_n444), .A2(G116), .ZN(new_n480));
  NAND2_X1  g280(.A1(G33), .A2(G283), .ZN(new_n481));
  INV_X1    g281(.A(G97), .ZN(new_n482));
  OAI211_X1 g282(.A(new_n481), .B(new_n218), .C1(G33), .C2(new_n482), .ZN(new_n483));
  OAI211_X1 g283(.A(new_n483), .B(new_n276), .C1(new_n218), .C2(G116), .ZN(new_n484));
  INV_X1    g284(.A(KEYINPUT20), .ZN(new_n485));
  AND2_X1   g285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g286(.A1(new_n484), .A2(new_n485), .ZN(new_n487));
  OAI221_X1 g287(.A(new_n480), .B1(G116), .B2(new_n280), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  NAND3_X1  g288(.A1(new_n479), .A2(G169), .A3(new_n488), .ZN(new_n489));
  INV_X1    g289(.A(KEYINPUT21), .ZN(new_n490));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g291(.A1(new_n479), .A2(G200), .ZN(new_n492));
  INV_X1    g292(.A(new_n488), .ZN(new_n493));
  OAI211_X1 g293(.A(new_n492), .B(new_n493), .C1(new_n305), .C2(new_n479), .ZN(new_n494));
  NOR2_X1   g294(.A1(new_n479), .A2(new_n366), .ZN(new_n495));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n488), .ZN(new_n496));
  NAND4_X1  g296(.A1(new_n479), .A2(KEYINPUT21), .A3(G169), .A4(new_n488), .ZN(new_n497));
  AND4_X1   g297(.A1(new_n491), .A2(new_n494), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  AND2_X1   g298(.A1(new_n461), .A2(G200), .ZN(new_n499));
  NOR2_X1   g299(.A1(new_n461), .A2(new_n305), .ZN(new_n500));
  NOR3_X1   g300(.A1(new_n448), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NOR2_X1   g301(.A1(new_n280), .A2(G97), .ZN(new_n502));
  INV_X1    g302(.A(new_n444), .ZN(new_n503));
  NOR2_X1   g303(.A1(new_n503), .A2(new_n482), .ZN(new_n504));
  NOR2_X1   g304(.A1(new_n482), .A2(G107), .ZN(new_n505));
  MUX2_X1   g305(.A(new_n238), .B(new_n505), .S(KEYINPUT6), .Z(new_n506));
  NAND2_X1  g306(.A1(new_n506), .A2(G20), .ZN(new_n507));
  OAI221_X1 g307(.A(new_n507), .B1(new_n385), .B2(new_n356), .C1(new_n271), .C2(new_n373), .ZN(new_n508));
  AOI211_X1 g308(.A(new_n502), .B(new_n504), .C1(new_n508), .C2(new_n276), .ZN(new_n509));
  INV_X1    g309(.A(new_n509), .ZN(new_n510));
  AND2_X1   g310(.A1(new_n307), .A2(G244), .ZN(new_n511));
  AOI21_X1  g311(.A(KEYINPUT4), .B1(new_n511), .B2(new_n370), .ZN(new_n512));
  NAND3_X1  g312(.A1(new_n344), .A2(KEYINPUT4), .A3(G244), .ZN(new_n513));
  INV_X1    g313(.A(KEYINPUT75), .ZN(new_n514));
  NAND3_X1  g314(.A1(new_n371), .A2(new_n514), .A3(G250), .ZN(new_n515));
  INV_X1    g315(.A(G250), .ZN(new_n516));
  OAI21_X1  g316(.A(KEYINPUT75), .B1(new_n347), .B2(new_n516), .ZN(new_n517));
  NAND4_X1  g317(.A1(new_n513), .A2(new_n515), .A3(new_n517), .A4(new_n481), .ZN(new_n518));
  OAI21_X1  g318(.A(new_n288), .B1(new_n512), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g319(.A1(new_n458), .A2(G257), .ZN(new_n520));
  NAND3_X1  g320(.A1(new_n519), .A2(new_n460), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n337), .ZN(new_n522));
  NAND4_X1  g322(.A1(new_n519), .A2(new_n366), .A3(new_n460), .A4(new_n520), .ZN(new_n523));
  NAND3_X1  g323(.A1(new_n510), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g324(.A1(new_n521), .A2(G200), .ZN(new_n525));
  OAI211_X1 g325(.A(new_n525), .B(new_n509), .C1(new_n305), .C2(new_n521), .ZN(new_n526));
  NAND2_X1  g326(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g327(.A1(new_n307), .A2(G238), .A3(new_n370), .ZN(new_n528));
  NAND2_X1  g328(.A1(new_n528), .A2(KEYINPUT77), .ZN(new_n529));
  NAND3_X1  g329(.A1(new_n307), .A2(G244), .A3(G1698), .ZN(new_n530));
  INV_X1    g330(.A(KEYINPUT77), .ZN(new_n531));
  NAND3_X1  g331(.A1(new_n312), .A2(new_n531), .A3(G238), .ZN(new_n532));
  NAND4_X1  g332(.A1(new_n529), .A2(new_n435), .A3(new_n530), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n288), .ZN(new_n534));
  NAND2_X1  g334(.A1(new_n283), .A2(G45), .ZN(new_n535));
  NAND3_X1  g335(.A1(new_n454), .A2(G250), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g336(.A(new_n536), .B1(new_n298), .B2(new_n535), .ZN(new_n537));
  INV_X1    g337(.A(KEYINPUT76), .ZN(new_n538));
  XNOR2_X1  g338(.A(new_n537), .B(new_n538), .ZN(new_n539));
  NAND2_X1  g339(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n337), .ZN(new_n541));
  INV_X1    g341(.A(KEYINPUT19), .ZN(new_n542));
  OAI21_X1  g342(.A(new_n542), .B1(new_n354), .B2(new_n482), .ZN(new_n543));
  XNOR2_X1  g343(.A(new_n543), .B(KEYINPUT78), .ZN(new_n544));
  NAND3_X1  g344(.A1(new_n373), .A2(new_n310), .A3(new_n482), .ZN(new_n545));
  OAI21_X1  g345(.A(new_n218), .B1(new_n396), .B2(new_n542), .ZN(new_n546));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g347(.A1(new_n307), .A2(new_n218), .A3(G68), .ZN(new_n548));
  NAND3_X1  g348(.A1(new_n544), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  AOI22_X1  g349(.A1(new_n549), .A2(new_n276), .B1(new_n279), .B2(new_n383), .ZN(new_n550));
  OAI21_X1  g350(.A(new_n550), .B1(new_n383), .B2(new_n503), .ZN(new_n551));
  OAI211_X1 g351(.A(new_n541), .B(new_n551), .C1(G179), .C2(new_n540), .ZN(new_n552));
  NAND2_X1  g352(.A1(new_n540), .A2(G200), .ZN(new_n553));
  NAND2_X1  g353(.A1(new_n444), .A2(G87), .ZN(new_n554));
  AND2_X1   g354(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g355(.A(new_n553), .B(new_n555), .C1(new_n305), .C2(new_n540), .ZN(new_n556));
  NAND2_X1  g356(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  NOR3_X1   g357(.A1(new_n501), .A2(new_n527), .A3(new_n557), .ZN(new_n558));
  AND4_X1   g358(.A1(new_n423), .A2(new_n468), .A3(new_n498), .A4(new_n558), .ZN(G372));
  INV_X1    g359(.A(new_n552), .ZN(new_n560));
  INV_X1    g360(.A(KEYINPUT26), .ZN(new_n561));
  OR3_X1    g361(.A1(new_n557), .A2(new_n561), .A3(new_n524), .ZN(new_n562));
  OAI21_X1  g362(.A(new_n561), .B1(new_n557), .B2(new_n524), .ZN(new_n563));
  AOI21_X1  g363(.A(new_n560), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g364(.A(new_n464), .ZN(new_n565));
  NAND3_X1  g365(.A1(new_n491), .A2(new_n496), .A3(new_n497), .ZN(new_n566));
  OAI21_X1  g366(.A(new_n558), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g367(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g368(.A1(new_n423), .A2(new_n568), .ZN(new_n569));
  INV_X1    g369(.A(new_n368), .ZN(new_n570));
  NAND2_X1  g370(.A1(new_n341), .A2(new_n342), .ZN(new_n571));
  INV_X1    g371(.A(new_n419), .ZN(new_n572));
  AOI21_X1  g372(.A(new_n572), .B1(new_n421), .B2(new_n390), .ZN(new_n573));
  NAND2_X1  g373(.A1(new_n324), .A2(new_n334), .ZN(new_n574));
  INV_X1    g374(.A(new_n574), .ZN(new_n575));
  OAI21_X1  g375(.A(new_n571), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g376(.A(new_n570), .B1(new_n576), .B2(new_n365), .ZN(new_n577));
  NAND2_X1  g377(.A1(new_n569), .A2(new_n577), .ZN(G369));
  AND2_X1   g378(.A1(new_n465), .A2(new_n467), .ZN(new_n579));
  NOR2_X1   g379(.A1(new_n579), .A2(new_n501), .ZN(new_n580));
  NOR2_X1   g380(.A1(new_n278), .A2(G20), .ZN(new_n581));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n283), .ZN(new_n582));
  OR2_X1    g382(.A1(new_n582), .A2(KEYINPUT27), .ZN(new_n583));
  NAND2_X1  g383(.A1(new_n582), .A2(KEYINPUT27), .ZN(new_n584));
  NAND3_X1  g384(.A1(new_n583), .A2(G213), .A3(new_n584), .ZN(new_n585));
  INV_X1    g385(.A(G343), .ZN(new_n586));
  NOR2_X1   g386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g387(.A(new_n587), .ZN(new_n588));
  AND2_X1   g388(.A1(new_n566), .A2(new_n588), .ZN(new_n589));
  AOI22_X1  g389(.A1(new_n580), .A2(new_n589), .B1(new_n565), .B2(new_n588), .ZN(new_n590));
  NAND2_X1  g390(.A1(new_n488), .A2(new_n587), .ZN(new_n591));
  MUX2_X1   g391(.A(new_n566), .B(new_n498), .S(new_n591), .Z(new_n592));
  XNOR2_X1  g392(.A(new_n592), .B(KEYINPUT82), .ZN(new_n593));
  NAND2_X1  g393(.A1(new_n593), .A2(G330), .ZN(new_n594));
  NAND2_X1  g394(.A1(new_n448), .A2(new_n587), .ZN(new_n595));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g396(.A1(new_n565), .A2(new_n587), .ZN(new_n597));
  NAND2_X1  g397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g398(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g399(.A(new_n590), .B1(new_n594), .B2(new_n599), .ZN(G399));
  INV_X1    g400(.A(new_n221), .ZN(new_n601));
  NOR2_X1   g401(.A1(new_n601), .A2(G41), .ZN(new_n602));
  INV_X1    g402(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g403(.A1(new_n603), .A2(G1), .ZN(new_n604));
  OR2_X1    g404(.A1(new_n545), .A2(G116), .ZN(new_n605));
  OAI22_X1  g405(.A1(new_n604), .A2(new_n605), .B1(new_n217), .B2(new_n603), .ZN(new_n606));
  XNOR2_X1  g406(.A(new_n606), .B(KEYINPUT28), .ZN(new_n607));
  INV_X1    g407(.A(G330), .ZN(new_n608));
  NAND4_X1  g408(.A1(new_n558), .A2(new_n468), .A3(new_n498), .A4(new_n588), .ZN(new_n609));
  NAND2_X1  g409(.A1(new_n609), .A2(KEYINPUT31), .ZN(new_n610));
  NAND2_X1  g410(.A1(new_n519), .A2(new_n520), .ZN(new_n611));
  NOR2_X1   g411(.A1(new_n611), .A2(new_n461), .ZN(new_n612));
  NAND4_X1  g412(.A1(new_n495), .A2(new_n534), .A3(new_n539), .A4(new_n612), .ZN(new_n613));
  XNOR2_X1  g413(.A(new_n613), .B(KEYINPUT30), .ZN(new_n614));
  NAND3_X1  g414(.A1(new_n479), .A2(new_n366), .A3(new_n521), .ZN(new_n615));
  NAND2_X1  g415(.A1(new_n540), .A2(new_n461), .ZN(new_n616));
  NOR2_X1   g416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g417(.A(new_n617), .B(KEYINPUT83), .ZN(new_n618));
  AOI21_X1  g418(.A(new_n588), .B1(new_n614), .B2(new_n618), .ZN(new_n619));
  INV_X1    g419(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g420(.A1(new_n610), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g421(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n622));
  NAND3_X1  g422(.A1(new_n622), .A2(KEYINPUT31), .A3(new_n587), .ZN(new_n623));
  AOI21_X1  g423(.A(new_n608), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g424(.A(new_n587), .B1(new_n564), .B2(new_n567), .ZN(new_n625));
  INV_X1    g425(.A(KEYINPUT29), .ZN(new_n626));
  AND2_X1   g426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g427(.A(new_n558), .B1(new_n579), .B2(new_n566), .ZN(new_n628));
  AOI21_X1  g428(.A(new_n587), .B1(new_n628), .B2(new_n564), .ZN(new_n629));
  NOR2_X1   g429(.A1(new_n629), .A2(new_n626), .ZN(new_n630));
  NOR3_X1   g430(.A1(new_n624), .A2(new_n627), .A3(new_n630), .ZN(new_n631));
  OAI21_X1  g431(.A(new_n607), .B1(new_n631), .B2(G1), .ZN(G364));
  AOI21_X1  g432(.A(new_n283), .B1(new_n581), .B2(G45), .ZN(new_n633));
  INV_X1    g433(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g434(.A1(new_n602), .A2(new_n634), .ZN(new_n635));
  INV_X1    g435(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g436(.A1(G179), .A2(G200), .ZN(new_n637));
  NAND3_X1  g437(.A1(new_n637), .A2(G20), .A3(new_n305), .ZN(new_n638));
  INV_X1    g438(.A(G329), .ZN(new_n639));
  OAI21_X1  g439(.A(new_n269), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g440(.A1(new_n218), .A2(new_n366), .ZN(new_n641));
  NAND2_X1  g441(.A1(new_n641), .A2(G200), .ZN(new_n642));
  NOR2_X1   g442(.A1(new_n642), .A2(G190), .ZN(new_n643));
  INV_X1    g443(.A(G317), .ZN(new_n644));
  NAND2_X1  g444(.A1(new_n644), .A2(KEYINPUT33), .ZN(new_n645));
  OR2_X1    g445(.A1(new_n644), .A2(KEYINPUT33), .ZN(new_n646));
  NAND3_X1  g446(.A1(new_n643), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  INV_X1    g447(.A(G283), .ZN(new_n648));
  NOR2_X1   g448(.A1(new_n218), .A2(G179), .ZN(new_n649));
  NAND3_X1  g449(.A1(new_n649), .A2(new_n305), .A3(G200), .ZN(new_n650));
  NAND3_X1  g450(.A1(new_n649), .A2(G190), .A3(G200), .ZN(new_n651));
  OAI221_X1 g451(.A(new_n647), .B1(new_n648), .B2(new_n650), .C1(new_n471), .C2(new_n651), .ZN(new_n652));
  NAND3_X1  g452(.A1(new_n641), .A2(G190), .A3(new_n330), .ZN(new_n653));
  OR2_X1    g453(.A1(new_n653), .A2(KEYINPUT85), .ZN(new_n654));
  NAND2_X1  g454(.A1(new_n653), .A2(KEYINPUT85), .ZN(new_n655));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AOI211_X1 g456(.A(new_n640), .B(new_n652), .C1(G322), .C2(new_n656), .ZN(new_n657));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n305), .ZN(new_n658));
  AOI21_X1  g458(.A(new_n218), .B1(new_n637), .B2(G190), .ZN(new_n659));
  INV_X1    g459(.A(new_n659), .ZN(new_n660));
  AOI22_X1  g460(.A1(new_n658), .A2(G326), .B1(G294), .B2(new_n660), .ZN(new_n661));
  XOR2_X1   g461(.A(new_n661), .B(KEYINPUT87), .Z(new_n662));
  INV_X1    g462(.A(G311), .ZN(new_n663));
  NAND3_X1  g463(.A1(new_n641), .A2(new_n305), .A3(new_n330), .ZN(new_n664));
  OAI211_X1 g464(.A(new_n657), .B(new_n662), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  XNOR2_X1  g465(.A(new_n665), .B(KEYINPUT88), .ZN(new_n666));
  NOR2_X1   g466(.A1(new_n659), .A2(new_n482), .ZN(new_n667));
  INV_X1    g467(.A(new_n664), .ZN(new_n668));
  AOI21_X1  g468(.A(new_n667), .B1(G77), .B2(new_n668), .ZN(new_n669));
  INV_X1    g469(.A(new_n658), .ZN(new_n670));
  INV_X1    g470(.A(new_n643), .ZN(new_n671));
  OAI221_X1 g471(.A(new_n669), .B1(new_n670), .B2(new_n202), .C1(new_n262), .C2(new_n671), .ZN(new_n672));
  AOI21_X1  g472(.A(new_n672), .B1(G58), .B2(new_n656), .ZN(new_n673));
  INV_X1    g473(.A(new_n650), .ZN(new_n674));
  NAND2_X1  g474(.A1(new_n674), .A2(G107), .ZN(new_n675));
  OAI211_X1 g475(.A(new_n675), .B(new_n245), .C1(new_n310), .C2(new_n651), .ZN(new_n676));
  OR2_X1    g476(.A1(new_n676), .A2(KEYINPUT86), .ZN(new_n677));
  NAND2_X1  g477(.A1(new_n676), .A2(KEYINPUT86), .ZN(new_n678));
  NAND3_X1  g478(.A1(new_n673), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  INV_X1    g479(.A(new_n638), .ZN(new_n680));
  NAND2_X1  g480(.A1(new_n680), .A2(G159), .ZN(new_n681));
  XNOR2_X1  g481(.A(new_n681), .B(KEYINPUT32), .ZN(new_n682));
  OAI21_X1  g482(.A(new_n666), .B1(new_n679), .B2(new_n682), .ZN(new_n683));
  AOI21_X1  g483(.A(new_n219), .B1(G20), .B2(new_n337), .ZN(new_n684));
  AOI21_X1  g484(.A(new_n636), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NOR2_X1   g485(.A1(G13), .A2(G33), .ZN(new_n686));
  XOR2_X1   g486(.A(new_n686), .B(KEYINPUT84), .Z(new_n687));
  INV_X1    g487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g488(.A1(new_n688), .A2(G20), .ZN(new_n689));
  INV_X1    g489(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g490(.A(new_n685), .B1(new_n593), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g491(.A1(new_n689), .A2(new_n684), .ZN(new_n692));
  NAND2_X1  g492(.A1(new_n237), .A2(G45), .ZN(new_n693));
  NOR2_X1   g493(.A1(new_n307), .A2(new_n601), .ZN(new_n694));
  OAI211_X1 g494(.A(new_n693), .B(new_n694), .C1(G45), .C2(new_n217), .ZN(new_n695));
  NOR2_X1   g495(.A1(new_n601), .A2(new_n269), .ZN(new_n696));
  NAND2_X1  g496(.A1(new_n696), .A2(G355), .ZN(new_n697));
  OAI211_X1 g497(.A(new_n695), .B(new_n697), .C1(G116), .C2(new_n221), .ZN(new_n698));
  AOI21_X1  g498(.A(new_n691), .B1(new_n692), .B2(new_n698), .ZN(new_n699));
  XNOR2_X1  g499(.A(new_n699), .B(KEYINPUT89), .ZN(new_n700));
  NOR2_X1   g500(.A1(new_n593), .A2(G330), .ZN(new_n701));
  NAND2_X1  g501(.A1(new_n594), .A2(new_n636), .ZN(new_n702));
  OAI21_X1  g502(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(G396));
  NOR2_X1   g503(.A1(new_n389), .A2(new_n587), .ZN(new_n704));
  INV_X1    g504(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g505(.A1(new_n388), .A2(new_n587), .ZN(new_n706));
  AND2_X1   g506(.A1(new_n393), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g507(.A(new_n705), .B1(new_n707), .B2(new_n390), .ZN(new_n708));
  OR2_X1    g508(.A1(new_n708), .A2(KEYINPUT90), .ZN(new_n709));
  NAND2_X1  g509(.A1(new_n708), .A2(KEYINPUT90), .ZN(new_n710));
  NAND2_X1  g510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g511(.A(new_n625), .B(new_n711), .ZN(new_n712));
  XNOR2_X1  g512(.A(new_n712), .B(new_n624), .ZN(new_n713));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n636), .ZN(new_n714));
  AOI22_X1  g514(.A1(new_n643), .A2(G150), .B1(new_n658), .B2(G137), .ZN(new_n715));
  INV_X1    g515(.A(G159), .ZN(new_n716));
  INV_X1    g516(.A(new_n656), .ZN(new_n717));
  INV_X1    g517(.A(G143), .ZN(new_n718));
  OAI221_X1 g518(.A(new_n715), .B1(new_n716), .B2(new_n664), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  XNOR2_X1  g519(.A(new_n719), .B(KEYINPUT34), .ZN(new_n720));
  OAI22_X1  g520(.A1(new_n202), .A2(new_n651), .B1(new_n650), .B2(new_n262), .ZN(new_n721));
  AOI211_X1 g521(.A(new_n247), .B(new_n721), .C1(G132), .C2(new_n680), .ZN(new_n722));
  OAI211_X1 g522(.A(new_n720), .B(new_n722), .C1(new_n261), .C2(new_n659), .ZN(new_n723));
  NOR2_X1   g523(.A1(new_n638), .A2(new_n663), .ZN(new_n724));
  NOR2_X1   g524(.A1(new_n650), .A2(new_n310), .ZN(new_n725));
  NOR2_X1   g525(.A1(new_n671), .A2(new_n648), .ZN(new_n726));
  INV_X1    g526(.A(new_n651), .ZN(new_n727));
  AOI211_X1 g527(.A(new_n725), .B(new_n726), .C1(G107), .C2(new_n727), .ZN(new_n728));
  OAI21_X1  g528(.A(new_n269), .B1(new_n664), .B2(new_n240), .ZN(new_n729));
  AOI211_X1 g529(.A(new_n667), .B(new_n729), .C1(G303), .C2(new_n658), .ZN(new_n730));
  OAI211_X1 g530(.A(new_n728), .B(new_n730), .C1(new_n451), .C2(new_n717), .ZN(new_n731));
  OAI21_X1  g531(.A(new_n723), .B1(new_n724), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g532(.A1(new_n684), .A2(new_n686), .ZN(new_n733));
  AOI22_X1  g533(.A1(new_n732), .A2(new_n684), .B1(new_n385), .B2(new_n733), .ZN(new_n734));
  OAI211_X1 g534(.A(new_n635), .B(new_n734), .C1(new_n711), .C2(new_n688), .ZN(new_n735));
  AND2_X1   g535(.A1(new_n714), .A2(new_n735), .ZN(new_n736));
  INV_X1    g536(.A(new_n736), .ZN(G384));
  NAND2_X1  g537(.A1(new_n418), .A2(new_n587), .ZN(new_n738));
  NAND3_X1  g538(.A1(new_n419), .A2(new_n421), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g539(.A(KEYINPUT91), .B1(new_n572), .B2(new_n587), .ZN(new_n740));
  INV_X1    g540(.A(KEYINPUT91), .ZN(new_n741));
  NOR3_X1   g541(.A1(new_n419), .A2(new_n741), .A3(new_n588), .ZN(new_n742));
  OAI21_X1  g542(.A(new_n739), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g543(.A(new_n619), .B1(new_n609), .B2(KEYINPUT31), .ZN(new_n744));
  NAND2_X1  g544(.A1(new_n619), .A2(KEYINPUT31), .ZN(new_n745));
  INV_X1    g545(.A(new_n745), .ZN(new_n746));
  OAI211_X1 g546(.A(new_n711), .B(new_n743), .C1(new_n744), .C2(new_n746), .ZN(new_n747));
  INV_X1    g547(.A(new_n747), .ZN(new_n748));
  INV_X1    g548(.A(KEYINPUT40), .ZN(new_n749));
  NAND2_X1  g549(.A1(new_n574), .A2(new_n571), .ZN(new_n750));
  NAND2_X1  g550(.A1(new_n267), .A2(new_n276), .ZN(new_n751));
  AOI21_X1  g551(.A(KEYINPUT16), .B1(new_n260), .B2(new_n266), .ZN(new_n752));
  OAI21_X1  g552(.A(new_n285), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g553(.A(new_n585), .ZN(new_n754));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g555(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g556(.A(KEYINPUT92), .B1(new_n750), .B2(new_n756), .ZN(new_n757));
  INV_X1    g557(.A(KEYINPUT92), .ZN(new_n758));
  NOR3_X1   g558(.A1(new_n343), .A2(new_n758), .A3(new_n755), .ZN(new_n759));
  INV_X1    g559(.A(KEYINPUT37), .ZN(new_n760));
  NAND2_X1  g560(.A1(new_n286), .A2(new_n754), .ZN(new_n761));
  NAND4_X1  g561(.A1(new_n323), .A2(new_n760), .A3(new_n339), .A4(new_n761), .ZN(new_n762));
  INV_X1    g562(.A(new_n762), .ZN(new_n763));
  NAND3_X1  g563(.A1(new_n336), .A2(new_n753), .A3(new_n338), .ZN(new_n764));
  NAND2_X1  g564(.A1(new_n323), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g565(.A(new_n756), .B1(new_n765), .B2(KEYINPUT93), .ZN(new_n766));
  INV_X1    g566(.A(KEYINPUT93), .ZN(new_n767));
  NAND3_X1  g567(.A1(new_n323), .A2(new_n767), .A3(new_n764), .ZN(new_n768));
  AOI21_X1  g568(.A(new_n760), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  OAI22_X1  g569(.A1(new_n757), .A2(new_n759), .B1(new_n763), .B2(new_n769), .ZN(new_n770));
  INV_X1    g570(.A(KEYINPUT38), .ZN(new_n771));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g572(.A1(new_n750), .A2(KEYINPUT92), .A3(new_n756), .ZN(new_n773));
  OAI21_X1  g573(.A(new_n758), .B1(new_n343), .B2(new_n755), .ZN(new_n774));
  AND3_X1   g574(.A1(new_n336), .A2(new_n753), .A3(new_n338), .ZN(new_n775));
  OAI21_X1  g575(.A(KEYINPUT93), .B1(new_n775), .B2(new_n332), .ZN(new_n776));
  NAND3_X1  g576(.A1(new_n776), .A2(new_n768), .A3(new_n755), .ZN(new_n777));
  NAND2_X1  g577(.A1(new_n777), .A2(KEYINPUT37), .ZN(new_n778));
  AOI22_X1  g578(.A1(new_n773), .A2(new_n774), .B1(new_n778), .B2(new_n762), .ZN(new_n779));
  NAND2_X1  g579(.A1(new_n779), .A2(KEYINPUT38), .ZN(new_n780));
  NAND3_X1  g580(.A1(new_n772), .A2(new_n780), .A3(KEYINPUT94), .ZN(new_n781));
  INV_X1    g581(.A(KEYINPUT94), .ZN(new_n782));
  NAND3_X1  g582(.A1(new_n779), .A2(new_n782), .A3(KEYINPUT38), .ZN(new_n783));
  NAND4_X1  g583(.A1(new_n748), .A2(new_n749), .A3(new_n781), .A4(new_n783), .ZN(new_n784));
  INV_X1    g584(.A(new_n761), .ZN(new_n785));
  INV_X1    g585(.A(KEYINPUT95), .ZN(new_n786));
  NAND2_X1  g586(.A1(new_n319), .A2(new_n320), .ZN(new_n787));
  AOI21_X1  g587(.A(new_n322), .B1(new_n787), .B2(new_n325), .ZN(new_n788));
  OAI211_X1 g588(.A(new_n339), .B(new_n761), .C1(new_n788), .C2(new_n286), .ZN(new_n789));
  AOI21_X1  g589(.A(new_n786), .B1(new_n789), .B2(KEYINPUT37), .ZN(new_n790));
  AOI22_X1  g590(.A1(new_n750), .A2(new_n785), .B1(new_n790), .B2(new_n762), .ZN(new_n791));
  NAND2_X1  g591(.A1(new_n763), .A2(new_n786), .ZN(new_n792));
  AOI21_X1  g592(.A(KEYINPUT38), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g593(.A(new_n793), .B1(KEYINPUT38), .B2(new_n779), .ZN(new_n794));
  OAI21_X1  g594(.A(KEYINPUT40), .B1(new_n747), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g595(.A1(new_n784), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g596(.A1(new_n621), .A2(new_n745), .ZN(new_n797));
  NAND2_X1  g597(.A1(new_n423), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g598(.A(new_n796), .B(new_n798), .ZN(new_n799));
  NAND2_X1  g599(.A1(new_n799), .A2(G330), .ZN(new_n800));
  AOI21_X1  g600(.A(new_n704), .B1(new_n625), .B2(new_n711), .ZN(new_n801));
  INV_X1    g601(.A(new_n801), .ZN(new_n802));
  NAND4_X1  g602(.A1(new_n802), .A2(new_n781), .A3(new_n743), .A4(new_n783), .ZN(new_n803));
  NAND3_X1  g603(.A1(new_n341), .A2(new_n342), .A3(new_n585), .ZN(new_n804));
  INV_X1    g604(.A(new_n793), .ZN(new_n805));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n780), .ZN(new_n806));
  INV_X1    g606(.A(KEYINPUT96), .ZN(new_n807));
  NOR3_X1   g607(.A1(new_n806), .A2(new_n807), .A3(KEYINPUT39), .ZN(new_n808));
  NAND3_X1  g608(.A1(new_n805), .A2(new_n780), .A3(new_n807), .ZN(new_n809));
  OAI21_X1  g609(.A(KEYINPUT94), .B1(new_n779), .B2(KEYINPUT38), .ZN(new_n810));
  NAND2_X1  g610(.A1(new_n773), .A2(new_n774), .ZN(new_n811));
  NAND2_X1  g611(.A1(new_n778), .A2(new_n762), .ZN(new_n812));
  AND3_X1   g612(.A1(new_n811), .A2(KEYINPUT38), .A3(new_n812), .ZN(new_n813));
  NOR2_X1   g613(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  INV_X1    g614(.A(new_n783), .ZN(new_n815));
  OAI21_X1  g615(.A(new_n809), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g616(.A(new_n808), .B1(new_n816), .B2(KEYINPUT39), .ZN(new_n817));
  NOR2_X1   g617(.A1(new_n419), .A2(new_n587), .ZN(new_n818));
  INV_X1    g618(.A(new_n818), .ZN(new_n819));
  OAI211_X1 g619(.A(new_n803), .B(new_n804), .C1(new_n817), .C2(new_n819), .ZN(new_n820));
  XOR2_X1   g620(.A(new_n800), .B(new_n820), .Z(new_n821));
  OAI21_X1  g621(.A(new_n423), .B1(new_n627), .B2(new_n630), .ZN(new_n822));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n577), .ZN(new_n823));
  XNOR2_X1  g623(.A(new_n821), .B(new_n823), .ZN(new_n824));
  OAI21_X1  g624(.A(new_n824), .B1(new_n283), .B2(new_n581), .ZN(new_n825));
  AOI21_X1  g625(.A(new_n240), .B1(new_n506), .B2(KEYINPUT35), .ZN(new_n826));
  NOR2_X1   g626(.A1(new_n219), .A2(new_n218), .ZN(new_n827));
  OAI211_X1 g627(.A(new_n826), .B(new_n827), .C1(KEYINPUT35), .C2(new_n506), .ZN(new_n828));
  XNOR2_X1  g628(.A(new_n828), .B(KEYINPUT36), .ZN(new_n829));
  OAI21_X1  g629(.A(G77), .B1(new_n261), .B2(new_n262), .ZN(new_n830));
  OAI22_X1  g630(.A1(new_n830), .A2(new_n217), .B1(G50), .B2(new_n262), .ZN(new_n831));
  NAND3_X1  g631(.A1(new_n831), .A2(G1), .A3(new_n278), .ZN(new_n832));
  NAND3_X1  g632(.A1(new_n825), .A2(new_n829), .A3(new_n832), .ZN(G367));
  INV_X1    g633(.A(new_n694), .ZN(new_n834));
  OAI221_X1 g634(.A(new_n692), .B1(new_n221), .B2(new_n383), .C1(new_n233), .C2(new_n834), .ZN(new_n835));
  NAND2_X1  g635(.A1(new_n643), .A2(G294), .ZN(new_n836));
  OAI221_X1 g636(.A(new_n836), .B1(new_n373), .B2(new_n659), .C1(new_n670), .C2(new_n663), .ZN(new_n837));
  AOI21_X1  g637(.A(new_n837), .B1(G97), .B2(new_n674), .ZN(new_n838));
  NAND2_X1  g638(.A1(new_n680), .A2(G317), .ZN(new_n839));
  AOI21_X1  g639(.A(KEYINPUT46), .B1(new_n727), .B2(G116), .ZN(new_n840));
  AOI21_X1  g640(.A(new_n840), .B1(new_n656), .B2(G303), .ZN(new_n841));
  AND3_X1   g641(.A1(new_n727), .A2(KEYINPUT46), .A3(G116), .ZN(new_n842));
  AOI211_X1 g642(.A(new_n307), .B(new_n842), .C1(G283), .C2(new_n668), .ZN(new_n843));
  NAND4_X1  g643(.A1(new_n838), .A2(new_n839), .A3(new_n841), .A4(new_n843), .ZN(new_n844));
  OAI22_X1  g644(.A1(new_n718), .A2(new_n670), .B1(new_n671), .B2(new_n716), .ZN(new_n845));
  AOI211_X1 g645(.A(new_n269), .B(new_n845), .C1(G137), .C2(new_n680), .ZN(new_n846));
  NOR2_X1   g646(.A1(new_n659), .A2(new_n262), .ZN(new_n847));
  NOR2_X1   g647(.A1(new_n650), .A2(new_n385), .ZN(new_n848));
  AOI211_X1 g648(.A(new_n847), .B(new_n848), .C1(G58), .C2(new_n727), .ZN(new_n849));
  OAI211_X1 g649(.A(new_n846), .B(new_n849), .C1(new_n355), .C2(new_n717), .ZN(new_n850));
  NOR2_X1   g650(.A1(new_n664), .A2(new_n202), .ZN(new_n851));
  OAI21_X1  g651(.A(new_n844), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  XNOR2_X1  g652(.A(new_n852), .B(KEYINPUT47), .ZN(new_n853));
  AOI21_X1  g653(.A(new_n636), .B1(new_n853), .B2(new_n684), .ZN(new_n854));
  OR2_X1    g654(.A1(new_n555), .A2(new_n588), .ZN(new_n855));
  NAND3_X1  g655(.A1(new_n552), .A2(new_n556), .A3(new_n855), .ZN(new_n856));
  OR2_X1    g656(.A1(new_n856), .A2(KEYINPUT97), .ZN(new_n857));
  NAND2_X1  g657(.A1(new_n856), .A2(KEYINPUT97), .ZN(new_n858));
  OAI211_X1 g658(.A(new_n857), .B(new_n858), .C1(new_n552), .C2(new_n855), .ZN(new_n859));
  OAI211_X1 g659(.A(new_n835), .B(new_n854), .C1(new_n859), .C2(new_n690), .ZN(new_n860));
  OAI211_X1 g660(.A(new_n524), .B(new_n526), .C1(new_n509), .C2(new_n588), .ZN(new_n861));
  OAI21_X1  g661(.A(new_n861), .B1(new_n524), .B2(new_n588), .ZN(new_n862));
  OR2_X1    g662(.A1(new_n590), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g663(.A1(new_n863), .A2(KEYINPUT100), .ZN(new_n864));
  AND2_X1   g664(.A1(KEYINPUT99), .A2(KEYINPUT44), .ZN(new_n865));
  NOR2_X1   g665(.A1(KEYINPUT99), .A2(KEYINPUT44), .ZN(new_n866));
  NOR3_X1   g666(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g667(.A1(new_n863), .A2(KEYINPUT100), .ZN(new_n868));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI211_X1 g669(.A(new_n863), .B(KEYINPUT100), .C1(new_n865), .C2(new_n866), .ZN(new_n870));
  NAND2_X1  g670(.A1(new_n590), .A2(new_n862), .ZN(new_n871));
  XOR2_X1   g671(.A(new_n871), .B(KEYINPUT45), .Z(new_n872));
  NAND3_X1  g672(.A1(new_n869), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  NOR2_X1   g673(.A1(new_n594), .A2(new_n599), .ZN(new_n874));
  OR2_X1    g674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g675(.A(KEYINPUT101), .ZN(new_n876));
  NAND3_X1  g676(.A1(new_n873), .A2(new_n876), .A3(new_n874), .ZN(new_n877));
  NAND2_X1  g677(.A1(new_n580), .A2(new_n589), .ZN(new_n878));
  OAI21_X1  g678(.A(new_n878), .B1(new_n598), .B2(new_n589), .ZN(new_n879));
  XOR2_X1   g679(.A(new_n594), .B(new_n879), .Z(new_n880));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n631), .ZN(new_n881));
  NAND2_X1  g681(.A1(new_n881), .A2(KEYINPUT102), .ZN(new_n882));
  OR2_X1    g682(.A1(new_n881), .A2(KEYINPUT102), .ZN(new_n883));
  NAND4_X1  g683(.A1(new_n875), .A2(new_n877), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  NOR2_X1   g684(.A1(new_n874), .A2(new_n876), .ZN(new_n885));
  OAI21_X1  g685(.A(new_n631), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  XNOR2_X1  g686(.A(new_n602), .B(KEYINPUT41), .ZN(new_n887));
  AOI21_X1  g687(.A(new_n634), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g688(.A1(new_n580), .A2(new_n589), .A3(new_n862), .ZN(new_n889));
  XOR2_X1   g689(.A(new_n889), .B(KEYINPUT42), .Z(new_n890));
  OAI21_X1  g690(.A(new_n524), .B1(new_n468), .B2(new_n861), .ZN(new_n891));
  XNOR2_X1  g691(.A(new_n891), .B(KEYINPUT98), .ZN(new_n892));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n588), .ZN(new_n893));
  AOI22_X1  g693(.A1(new_n890), .A2(new_n893), .B1(KEYINPUT43), .B2(new_n859), .ZN(new_n894));
  NOR2_X1   g694(.A1(new_n859), .A2(KEYINPUT43), .ZN(new_n895));
  XNOR2_X1  g695(.A(new_n894), .B(new_n895), .ZN(new_n896));
  NAND2_X1  g696(.A1(new_n874), .A2(new_n862), .ZN(new_n897));
  XOR2_X1   g697(.A(new_n896), .B(new_n897), .Z(new_n898));
  OAI21_X1  g698(.A(new_n860), .B1(new_n888), .B2(new_n898), .ZN(G387));
  OR2_X1    g699(.A1(new_n880), .A2(new_n631), .ZN(new_n900));
  NAND3_X1  g700(.A1(new_n900), .A2(new_n602), .A3(new_n881), .ZN(new_n901));
  NAND2_X1  g701(.A1(new_n880), .A2(new_n634), .ZN(new_n902));
  XOR2_X1   g702(.A(KEYINPUT106), .B(G322), .Z(new_n903));
  OAI22_X1  g703(.A1(new_n670), .A2(new_n903), .B1(new_n671), .B2(new_n663), .ZN(new_n904));
  AOI21_X1  g704(.A(new_n904), .B1(G317), .B2(new_n656), .ZN(new_n905));
  OAI21_X1  g705(.A(new_n905), .B1(new_n471), .B2(new_n664), .ZN(new_n906));
  XNOR2_X1  g706(.A(new_n906), .B(KEYINPUT48), .ZN(new_n907));
  OAI22_X1  g707(.A1(new_n651), .A2(new_n451), .B1(new_n659), .B2(new_n648), .ZN(new_n908));
  XOR2_X1   g708(.A(new_n908), .B(KEYINPUT105), .Z(new_n909));
  NAND2_X1  g709(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g710(.A(KEYINPUT107), .B(KEYINPUT49), .ZN(new_n911));
  OR2_X1    g711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g712(.A1(new_n680), .A2(G326), .ZN(new_n913));
  NAND2_X1  g713(.A1(new_n910), .A2(new_n911), .ZN(new_n914));
  AOI21_X1  g714(.A(new_n307), .B1(G116), .B2(new_n674), .ZN(new_n915));
  NAND4_X1  g715(.A1(new_n912), .A2(new_n913), .A3(new_n914), .A4(new_n915), .ZN(new_n916));
  OAI22_X1  g716(.A1(new_n651), .A2(new_n385), .B1(new_n355), .B2(new_n638), .ZN(new_n917));
  INV_X1    g717(.A(KEYINPUT103), .ZN(new_n918));
  AOI21_X1  g718(.A(new_n247), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI221_X1 g719(.A(new_n919), .B1(new_n918), .B2(new_n917), .C1(new_n482), .C2(new_n650), .ZN(new_n920));
  XOR2_X1   g720(.A(new_n920), .B(KEYINPUT104), .Z(new_n921));
  AOI22_X1  g721(.A1(new_n668), .A2(G68), .B1(new_n660), .B2(new_n382), .ZN(new_n922));
  OAI21_X1  g722(.A(new_n922), .B1(new_n716), .B2(new_n670), .ZN(new_n923));
  AOI21_X1  g723(.A(new_n923), .B1(G50), .B2(new_n656), .ZN(new_n924));
  OAI211_X1 g724(.A(new_n921), .B(new_n924), .C1(new_n281), .C2(new_n671), .ZN(new_n925));
  NAND2_X1  g725(.A1(new_n916), .A2(new_n925), .ZN(new_n926));
  OR2_X1    g726(.A1(new_n229), .A2(new_n290), .ZN(new_n927));
  AOI22_X1  g727(.A1(new_n927), .A2(new_n694), .B1(new_n605), .B2(new_n696), .ZN(new_n928));
  NOR2_X1   g728(.A1(new_n281), .A2(G50), .ZN(new_n929));
  XNOR2_X1  g729(.A(new_n929), .B(KEYINPUT50), .ZN(new_n930));
  OAI21_X1  g730(.A(new_n930), .B1(new_n262), .B2(new_n385), .ZN(new_n931));
  NOR3_X1   g731(.A1(new_n931), .A2(G45), .A3(new_n605), .ZN(new_n932));
  OAI22_X1  g732(.A1(new_n928), .A2(new_n932), .B1(G107), .B2(new_n221), .ZN(new_n933));
  AOI22_X1  g733(.A1(new_n926), .A2(new_n684), .B1(new_n692), .B2(new_n933), .ZN(new_n934));
  OAI211_X1 g734(.A(new_n934), .B(new_n635), .C1(new_n598), .C2(new_n690), .ZN(new_n935));
  NAND3_X1  g735(.A1(new_n901), .A2(new_n902), .A3(new_n935), .ZN(G393));
  NAND2_X1  g736(.A1(new_n873), .A2(new_n874), .ZN(new_n937));
  NAND2_X1  g737(.A1(new_n875), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n881), .ZN(new_n939));
  OAI211_X1 g739(.A(new_n939), .B(new_n602), .C1(new_n884), .C2(new_n885), .ZN(new_n940));
  AOI22_X1  g740(.A1(new_n656), .A2(G311), .B1(G317), .B2(new_n658), .ZN(new_n941));
  XNOR2_X1  g741(.A(new_n941), .B(KEYINPUT111), .ZN(new_n942));
  XNOR2_X1  g742(.A(new_n942), .B(KEYINPUT52), .ZN(new_n943));
  OAI221_X1 g743(.A(new_n269), .B1(new_n903), .B2(new_n638), .C1(new_n451), .C2(new_n664), .ZN(new_n944));
  OAI21_X1  g744(.A(new_n675), .B1(new_n671), .B2(new_n471), .ZN(new_n945));
  AOI211_X1 g745(.A(new_n944), .B(new_n945), .C1(G283), .C2(new_n727), .ZN(new_n946));
  OAI211_X1 g746(.A(new_n943), .B(new_n946), .C1(new_n240), .C2(new_n659), .ZN(new_n947));
  AOI22_X1  g747(.A1(G50), .A2(new_n643), .B1(new_n668), .B2(new_n380), .ZN(new_n948));
  XNOR2_X1  g748(.A(new_n948), .B(KEYINPUT110), .ZN(new_n949));
  AOI21_X1  g749(.A(new_n725), .B1(G68), .B2(new_n727), .ZN(new_n950));
  NOR2_X1   g750(.A1(new_n659), .A2(new_n385), .ZN(new_n951));
  AOI211_X1 g751(.A(new_n951), .B(new_n247), .C1(G143), .C2(new_n680), .ZN(new_n952));
  NAND3_X1  g752(.A1(new_n949), .A2(new_n950), .A3(new_n952), .ZN(new_n953));
  AOI22_X1  g753(.A1(new_n656), .A2(G159), .B1(G150), .B2(new_n658), .ZN(new_n954));
  XNOR2_X1  g754(.A(KEYINPUT109), .B(KEYINPUT51), .ZN(new_n955));
  XOR2_X1   g755(.A(new_n954), .B(new_n955), .Z(new_n956));
  OAI21_X1  g756(.A(new_n947), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g757(.A(new_n636), .B1(new_n957), .B2(new_n684), .ZN(new_n958));
  OAI221_X1 g758(.A(new_n692), .B1(new_n482), .B2(new_n221), .C1(new_n241), .C2(new_n834), .ZN(new_n959));
  OAI211_X1 g759(.A(new_n958), .B(new_n959), .C1(new_n690), .C2(new_n862), .ZN(new_n960));
  INV_X1    g760(.A(KEYINPUT108), .ZN(new_n961));
  NAND2_X1  g761(.A1(new_n938), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g762(.A1(new_n875), .A2(KEYINPUT108), .A3(new_n937), .ZN(new_n963));
  NAND3_X1  g763(.A1(new_n962), .A2(new_n634), .A3(new_n963), .ZN(new_n964));
  NAND3_X1  g764(.A1(new_n940), .A2(new_n960), .A3(new_n964), .ZN(G390));
  INV_X1    g765(.A(KEYINPUT39), .ZN(new_n966));
  NAND3_X1  g766(.A1(new_n794), .A2(KEYINPUT96), .A3(new_n966), .ZN(new_n967));
  INV_X1    g767(.A(new_n743), .ZN(new_n968));
  OAI21_X1  g768(.A(new_n819), .B1(new_n801), .B2(new_n968), .ZN(new_n969));
  AOI22_X1  g769(.A1(new_n781), .A2(new_n783), .B1(new_n794), .B2(new_n807), .ZN(new_n970));
  OAI211_X1 g770(.A(new_n967), .B(new_n969), .C1(new_n970), .C2(new_n966), .ZN(new_n971));
  AOI21_X1  g771(.A(new_n704), .B1(new_n629), .B2(new_n711), .ZN(new_n972));
  OAI211_X1 g772(.A(new_n806), .B(new_n819), .C1(new_n972), .C2(new_n968), .ZN(new_n973));
  NAND3_X1  g773(.A1(new_n624), .A2(new_n711), .A3(new_n743), .ZN(new_n974));
  INV_X1    g774(.A(new_n974), .ZN(new_n975));
  AND3_X1   g775(.A1(new_n971), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  NOR2_X1   g776(.A1(new_n747), .A2(new_n608), .ZN(new_n977));
  AOI21_X1  g777(.A(new_n977), .B1(new_n971), .B2(new_n973), .ZN(new_n978));
  NOR2_X1   g778(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g779(.A1(new_n423), .A2(new_n797), .A3(G330), .ZN(new_n980));
  NAND3_X1  g780(.A1(new_n822), .A2(new_n980), .A3(new_n577), .ZN(new_n981));
  INV_X1    g781(.A(new_n981), .ZN(new_n982));
  INV_X1    g782(.A(new_n623), .ZN(new_n983));
  OAI211_X1 g783(.A(G330), .B(new_n711), .C1(new_n983), .C2(new_n744), .ZN(new_n984));
  AOI22_X1  g784(.A1(new_n748), .A2(G330), .B1(new_n968), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g785(.A1(new_n985), .A2(new_n801), .ZN(new_n986));
  OAI211_X1 g786(.A(G330), .B(new_n711), .C1(new_n744), .C2(new_n746), .ZN(new_n987));
  NAND2_X1  g787(.A1(new_n987), .A2(new_n968), .ZN(new_n988));
  NAND3_X1  g788(.A1(new_n974), .A2(new_n988), .A3(new_n972), .ZN(new_n989));
  INV_X1    g789(.A(new_n989), .ZN(new_n990));
  OAI21_X1  g790(.A(new_n982), .B1(new_n986), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g791(.A(new_n602), .B1(new_n979), .B2(new_n991), .ZN(new_n992));
  AOI21_X1  g792(.A(new_n992), .B1(new_n979), .B2(new_n991), .ZN(new_n993));
  INV_X1    g793(.A(G128), .ZN(new_n994));
  NOR2_X1   g794(.A1(new_n670), .A2(new_n994), .ZN(new_n995));
  INV_X1    g795(.A(G137), .ZN(new_n996));
  OAI22_X1  g796(.A1(new_n671), .A2(new_n996), .B1(new_n202), .B2(new_n650), .ZN(new_n997));
  AOI211_X1 g797(.A(new_n995), .B(new_n997), .C1(G159), .C2(new_n660), .ZN(new_n998));
  NAND2_X1  g798(.A1(new_n680), .A2(G125), .ZN(new_n999));
  NOR2_X1   g799(.A1(new_n651), .A2(new_n355), .ZN(new_n1000));
  XOR2_X1   g800(.A(KEYINPUT112), .B(KEYINPUT53), .Z(new_n1001));
  XNOR2_X1  g801(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g802(.A(KEYINPUT54), .B(G143), .ZN(new_n1003));
  OAI21_X1  g803(.A(new_n245), .B1(new_n664), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g804(.A(new_n1004), .B1(new_n656), .B2(G132), .ZN(new_n1005));
  NAND4_X1  g805(.A1(new_n998), .A2(new_n999), .A3(new_n1002), .A4(new_n1005), .ZN(new_n1006));
  NOR2_X1   g806(.A1(new_n671), .A2(new_n373), .ZN(new_n1007));
  AOI211_X1 g807(.A(new_n951), .B(new_n1007), .C1(G283), .C2(new_n658), .ZN(new_n1008));
  OAI22_X1  g808(.A1(new_n262), .A2(new_n650), .B1(new_n651), .B2(new_n310), .ZN(new_n1009));
  AOI211_X1 g809(.A(new_n245), .B(new_n1009), .C1(G97), .C2(new_n668), .ZN(new_n1010));
  OAI211_X1 g810(.A(new_n1008), .B(new_n1010), .C1(new_n240), .C2(new_n717), .ZN(new_n1011));
  NOR2_X1   g811(.A1(new_n638), .A2(new_n451), .ZN(new_n1012));
  OAI21_X1  g812(.A(new_n1006), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AOI22_X1  g813(.A1(new_n1013), .A2(new_n684), .B1(new_n281), .B2(new_n733), .ZN(new_n1014));
  OAI21_X1  g814(.A(new_n967), .B1(new_n970), .B2(new_n966), .ZN(new_n1015));
  OAI211_X1 g815(.A(new_n635), .B(new_n1014), .C1(new_n1015), .C2(new_n688), .ZN(new_n1016));
  OAI21_X1  g816(.A(new_n1016), .B1(new_n979), .B2(new_n633), .ZN(new_n1017));
  NOR2_X1   g817(.A1(new_n993), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g818(.A(new_n1018), .ZN(G378));
  INV_X1    g819(.A(KEYINPUT57), .ZN(new_n1020));
  NAND2_X1  g820(.A1(new_n971), .A2(new_n973), .ZN(new_n1021));
  INV_X1    g821(.A(new_n977), .ZN(new_n1022));
  NAND2_X1  g822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g823(.A1(new_n971), .A2(new_n973), .A3(new_n975), .ZN(new_n1024));
  AOI21_X1  g824(.A(new_n991), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g825(.A(KEYINPUT117), .B1(new_n1025), .B2(new_n981), .ZN(new_n1026));
  INV_X1    g826(.A(KEYINPUT117), .ZN(new_n1027));
  OAI211_X1 g827(.A(new_n1027), .B(new_n982), .C1(new_n979), .C2(new_n991), .ZN(new_n1028));
  NAND2_X1  g828(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g829(.A1(new_n796), .A2(G330), .ZN(new_n1030));
  INV_X1    g830(.A(new_n1030), .ZN(new_n1031));
  NAND2_X1  g831(.A1(new_n820), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g832(.A1(new_n360), .A2(new_n754), .ZN(new_n1033));
  XNOR2_X1  g833(.A(new_n369), .B(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g834(.A(new_n1034), .B(KEYINPUT55), .ZN(new_n1035));
  INV_X1    g835(.A(KEYINPUT56), .ZN(new_n1036));
  XNOR2_X1  g836(.A(new_n1035), .B(new_n1036), .ZN(new_n1037));
  NAND2_X1  g837(.A1(new_n1015), .A2(new_n818), .ZN(new_n1038));
  NAND4_X1  g838(.A1(new_n1038), .A2(new_n1030), .A3(new_n803), .A4(new_n804), .ZN(new_n1039));
  AND3_X1   g839(.A1(new_n1032), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g840(.A(new_n1037), .B1(new_n1032), .B2(new_n1039), .ZN(new_n1041));
  NOR2_X1   g841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g842(.A(new_n1020), .B1(new_n1029), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g843(.A1(new_n1032), .A2(new_n1039), .ZN(new_n1044));
  INV_X1    g844(.A(new_n1037), .ZN(new_n1045));
  NAND2_X1  g845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g846(.A1(new_n1032), .A2(new_n1039), .A3(new_n1037), .ZN(new_n1047));
  NAND2_X1  g847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g848(.A1(new_n1048), .A2(KEYINPUT57), .A3(new_n1026), .A4(new_n1028), .ZN(new_n1049));
  NAND3_X1  g849(.A1(new_n1043), .A2(new_n602), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g850(.A1(new_n733), .A2(new_n202), .ZN(new_n1051));
  OAI22_X1  g851(.A1(new_n670), .A2(new_n240), .B1(new_n651), .B2(new_n385), .ZN(new_n1052));
  AOI21_X1  g852(.A(new_n1052), .B1(G97), .B2(new_n643), .ZN(new_n1053));
  NOR2_X1   g853(.A1(new_n638), .A2(new_n648), .ZN(new_n1054));
  AOI211_X1 g854(.A(new_n847), .B(new_n1054), .C1(new_n656), .C2(G107), .ZN(new_n1055));
  NAND2_X1  g855(.A1(new_n674), .A2(G58), .ZN(new_n1056));
  AOI211_X1 g856(.A(G41), .B(new_n307), .C1(new_n382), .C2(new_n668), .ZN(new_n1057));
  NAND4_X1  g857(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g858(.A(new_n1058), .B(KEYINPUT58), .ZN(new_n1059));
  NOR2_X1   g859(.A1(G33), .A2(G41), .ZN(new_n1060));
  XNOR2_X1  g860(.A(new_n1060), .B(KEYINPUT113), .ZN(new_n1061));
  OAI211_X1 g861(.A(new_n202), .B(new_n1061), .C1(new_n307), .C2(G41), .ZN(new_n1062));
  AOI21_X1  g862(.A(new_n1061), .B1(G159), .B2(new_n674), .ZN(new_n1063));
  INV_X1    g863(.A(G124), .ZN(new_n1064));
  OAI21_X1  g864(.A(new_n1063), .B1(new_n1064), .B2(new_n638), .ZN(new_n1065));
  XNOR2_X1  g865(.A(new_n1065), .B(KEYINPUT114), .ZN(new_n1066));
  AOI22_X1  g866(.A1(new_n656), .A2(G128), .B1(G125), .B2(new_n658), .ZN(new_n1067));
  OAI22_X1  g867(.A1(new_n651), .A2(new_n1003), .B1(new_n659), .B2(new_n355), .ZN(new_n1068));
  AOI21_X1  g868(.A(new_n1068), .B1(G132), .B2(new_n643), .ZN(new_n1069));
  OAI211_X1 g869(.A(new_n1067), .B(new_n1069), .C1(new_n996), .C2(new_n664), .ZN(new_n1070));
  XNOR2_X1  g870(.A(new_n1070), .B(KEYINPUT59), .ZN(new_n1071));
  OAI211_X1 g871(.A(new_n1059), .B(new_n1062), .C1(new_n1066), .C2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g872(.A(new_n636), .B1(new_n1072), .B2(new_n684), .ZN(new_n1073));
  OAI211_X1 g873(.A(new_n1051), .B(new_n1073), .C1(new_n1045), .C2(new_n688), .ZN(new_n1074));
  INV_X1    g874(.A(KEYINPUT115), .ZN(new_n1075));
  XNOR2_X1  g875(.A(new_n1074), .B(new_n1075), .ZN(new_n1076));
  NAND2_X1  g876(.A1(new_n1076), .A2(KEYINPUT116), .ZN(new_n1077));
  NOR2_X1   g877(.A1(new_n1076), .A2(KEYINPUT116), .ZN(new_n1078));
  AOI21_X1  g878(.A(new_n1078), .B1(new_n634), .B2(new_n1048), .ZN(new_n1079));
  NAND3_X1  g879(.A1(new_n1050), .A2(new_n1077), .A3(new_n1079), .ZN(G375));
  OAI21_X1  g880(.A(new_n634), .B1(new_n986), .B2(new_n990), .ZN(new_n1081));
  INV_X1    g881(.A(KEYINPUT118), .ZN(new_n1082));
  NAND2_X1  g882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g883(.A1(new_n733), .A2(new_n262), .ZN(new_n1084));
  NOR2_X1   g884(.A1(new_n717), .A2(new_n648), .ZN(new_n1085));
  OAI22_X1  g885(.A1(new_n670), .A2(new_n451), .B1(new_n659), .B2(new_n383), .ZN(new_n1086));
  OAI21_X1  g886(.A(new_n269), .B1(new_n638), .B2(new_n471), .ZN(new_n1087));
  NOR4_X1   g887(.A1(new_n1085), .A2(new_n848), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  OAI22_X1  g888(.A1(new_n671), .A2(new_n240), .B1(new_n664), .B2(new_n373), .ZN(new_n1089));
  XNOR2_X1  g889(.A(new_n1089), .B(KEYINPUT119), .ZN(new_n1090));
  OAI211_X1 g890(.A(new_n1088), .B(new_n1090), .C1(new_n482), .C2(new_n651), .ZN(new_n1091));
  XOR2_X1   g891(.A(new_n1091), .B(KEYINPUT120), .Z(new_n1092));
  AOI22_X1  g892(.A1(new_n727), .A2(G159), .B1(new_n674), .B2(G58), .ZN(new_n1093));
  NAND2_X1  g893(.A1(new_n658), .A2(G132), .ZN(new_n1094));
  OAI211_X1 g894(.A(new_n1093), .B(new_n1094), .C1(new_n671), .C2(new_n1003), .ZN(new_n1095));
  AOI211_X1 g895(.A(new_n247), .B(new_n1095), .C1(G137), .C2(new_n656), .ZN(new_n1096));
  OAI22_X1  g896(.A1(new_n664), .A2(new_n355), .B1(new_n659), .B2(new_n202), .ZN(new_n1097));
  XNOR2_X1  g897(.A(new_n1097), .B(KEYINPUT121), .ZN(new_n1098));
  OAI211_X1 g898(.A(new_n1096), .B(new_n1098), .C1(new_n994), .C2(new_n638), .ZN(new_n1099));
  NAND2_X1  g899(.A1(new_n1092), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g900(.A(new_n636), .B1(new_n1100), .B2(new_n684), .ZN(new_n1101));
  INV_X1    g901(.A(new_n686), .ZN(new_n1102));
  OAI211_X1 g902(.A(new_n1084), .B(new_n1101), .C1(new_n743), .C2(new_n1102), .ZN(new_n1103));
  OAI211_X1 g903(.A(KEYINPUT118), .B(new_n634), .C1(new_n986), .C2(new_n990), .ZN(new_n1104));
  NAND3_X1  g904(.A1(new_n1083), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g905(.A(new_n1105), .ZN(new_n1106));
  OAI211_X1 g906(.A(new_n989), .B(new_n981), .C1(new_n985), .C2(new_n801), .ZN(new_n1107));
  NAND3_X1  g907(.A1(new_n991), .A2(new_n887), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g908(.A1(new_n1106), .A2(new_n1108), .ZN(G381));
  OR2_X1    g909(.A1(G375), .A2(G378), .ZN(new_n1110));
  OR3_X1    g910(.A1(G390), .A2(G396), .A3(G393), .ZN(new_n1111));
  NOR4_X1   g911(.A1(new_n1111), .A2(G384), .A3(G387), .A4(G381), .ZN(new_n1112));
  AOI21_X1  g912(.A(new_n1110), .B1(new_n1112), .B2(KEYINPUT122), .ZN(new_n1113));
  OAI21_X1  g913(.A(new_n1113), .B1(KEYINPUT122), .B2(new_n1112), .ZN(G407));
  OAI211_X1 g914(.A(G407), .B(G213), .C1(G343), .C2(new_n1110), .ZN(G409));
  NAND2_X1  g915(.A1(G375), .A2(G378), .ZN(new_n1116));
  NAND4_X1  g916(.A1(new_n1048), .A2(new_n887), .A3(new_n1026), .A4(new_n1028), .ZN(new_n1117));
  NAND2_X1  g917(.A1(new_n1048), .A2(new_n634), .ZN(new_n1118));
  NAND4_X1  g918(.A1(new_n1018), .A2(new_n1076), .A3(new_n1117), .A4(new_n1118), .ZN(new_n1119));
  NAND2_X1  g919(.A1(new_n586), .A2(G213), .ZN(new_n1120));
  NAND2_X1  g920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g921(.A(new_n1121), .ZN(new_n1122));
  INV_X1    g922(.A(KEYINPUT125), .ZN(new_n1123));
  NAND2_X1  g923(.A1(new_n1107), .A2(KEYINPUT123), .ZN(new_n1124));
  NAND2_X1  g924(.A1(new_n1124), .A2(KEYINPUT60), .ZN(new_n1125));
  INV_X1    g925(.A(KEYINPUT60), .ZN(new_n1126));
  NAND3_X1  g926(.A1(new_n1107), .A2(KEYINPUT123), .A3(new_n1126), .ZN(new_n1127));
  NAND4_X1  g927(.A1(new_n1125), .A2(new_n602), .A3(new_n991), .A4(new_n1127), .ZN(new_n1128));
  NAND2_X1  g928(.A1(new_n1128), .A2(KEYINPUT124), .ZN(new_n1129));
  AND2_X1   g929(.A1(new_n1127), .A2(new_n991), .ZN(new_n1130));
  INV_X1    g930(.A(KEYINPUT124), .ZN(new_n1131));
  AOI21_X1  g931(.A(new_n603), .B1(new_n1124), .B2(KEYINPUT60), .ZN(new_n1132));
  NAND3_X1  g932(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g933(.A(new_n1105), .B1(new_n1129), .B2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g934(.A1(new_n1134), .A2(G384), .ZN(new_n1135));
  AOI211_X1 g935(.A(new_n736), .B(new_n1105), .C1(new_n1129), .C2(new_n1133), .ZN(new_n1136));
  OAI21_X1  g936(.A(new_n1123), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g937(.A1(new_n1128), .A2(KEYINPUT124), .ZN(new_n1138));
  AOI21_X1  g938(.A(new_n1131), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1139));
  OAI21_X1  g939(.A(new_n1106), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g940(.A1(new_n1140), .A2(new_n736), .ZN(new_n1141));
  NAND2_X1  g941(.A1(new_n1134), .A2(G384), .ZN(new_n1142));
  NAND3_X1  g942(.A1(new_n1141), .A2(KEYINPUT125), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g943(.A1(new_n1137), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g944(.A1(new_n1116), .A2(new_n1122), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g945(.A(KEYINPUT127), .ZN(new_n1146));
  INV_X1    g946(.A(KEYINPUT62), .ZN(new_n1147));
  NAND2_X1  g947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g948(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1149));
  NAND3_X1  g949(.A1(new_n1145), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g950(.A1(new_n1116), .A2(new_n1122), .ZN(new_n1151));
  NAND3_X1  g951(.A1(new_n586), .A2(G213), .A3(G2897), .ZN(new_n1152));
  AOI21_X1  g952(.A(new_n1152), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1153));
  AOI21_X1  g953(.A(new_n1153), .B1(new_n1144), .B2(new_n1152), .ZN(new_n1154));
  AOI21_X1  g954(.A(KEYINPUT61), .B1(new_n1151), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g955(.A(new_n1121), .B1(G375), .B2(G378), .ZN(new_n1156));
  NAND4_X1  g956(.A1(new_n1156), .A2(new_n1146), .A3(new_n1147), .A4(new_n1144), .ZN(new_n1157));
  NAND3_X1  g957(.A1(new_n1150), .A2(new_n1155), .A3(new_n1157), .ZN(new_n1158));
  XOR2_X1   g958(.A(G393), .B(G396), .Z(new_n1159));
  INV_X1    g959(.A(G390), .ZN(new_n1160));
  NAND2_X1  g960(.A1(G387), .A2(new_n1160), .ZN(new_n1161));
  OAI211_X1 g961(.A(G390), .B(new_n860), .C1(new_n888), .C2(new_n898), .ZN(new_n1162));
  AOI21_X1  g962(.A(new_n1159), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g963(.A(new_n1163), .ZN(new_n1164));
  NAND3_X1  g964(.A1(new_n1161), .A2(new_n1159), .A3(new_n1162), .ZN(new_n1165));
  NAND2_X1  g965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g966(.A1(new_n1158), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g967(.A1(new_n1154), .A2(KEYINPUT126), .ZN(new_n1168));
  INV_X1    g968(.A(KEYINPUT126), .ZN(new_n1169));
  INV_X1    g969(.A(new_n1152), .ZN(new_n1170));
  AOI21_X1  g970(.A(new_n1170), .B1(new_n1137), .B2(new_n1143), .ZN(new_n1171));
  OAI21_X1  g971(.A(new_n1169), .B1(new_n1171), .B2(new_n1153), .ZN(new_n1172));
  NAND3_X1  g972(.A1(new_n1168), .A2(new_n1172), .A3(new_n1151), .ZN(new_n1173));
  AND2_X1   g973(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1174));
  INV_X1    g974(.A(KEYINPUT63), .ZN(new_n1175));
  AOI21_X1  g975(.A(KEYINPUT61), .B1(new_n1145), .B2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g976(.A1(new_n1156), .A2(KEYINPUT63), .A3(new_n1144), .ZN(new_n1177));
  NAND4_X1  g977(.A1(new_n1173), .A2(new_n1174), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  NAND2_X1  g978(.A1(new_n1167), .A2(new_n1178), .ZN(G405));
  AND3_X1   g979(.A1(new_n1110), .A2(new_n1116), .A3(new_n1144), .ZN(new_n1180));
  NOR2_X1   g980(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1181));
  AOI21_X1  g981(.A(new_n1181), .B1(new_n1110), .B2(new_n1116), .ZN(new_n1182));
  OAI21_X1  g982(.A(new_n1174), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g983(.A1(new_n1110), .A2(new_n1116), .A3(new_n1144), .ZN(new_n1184));
  AND2_X1   g984(.A1(new_n1110), .A2(new_n1116), .ZN(new_n1185));
  OAI211_X1 g985(.A(new_n1166), .B(new_n1184), .C1(new_n1185), .C2(new_n1181), .ZN(new_n1186));
  AND2_X1   g986(.A1(new_n1183), .A2(new_n1186), .ZN(G402));
endmodule


