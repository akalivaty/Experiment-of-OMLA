

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592;

  AND2_X1 U324 ( .A1(G230GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U325 ( .A(n426), .B(n334), .ZN(n338) );
  XNOR2_X1 U326 ( .A(n394), .B(n342), .ZN(n343) );
  XNOR2_X1 U327 ( .A(n344), .B(n343), .ZN(n582) );
  XOR2_X1 U328 ( .A(n420), .B(n419), .Z(n533) );
  XNOR2_X1 U329 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U330 ( .A(n463), .B(n462), .ZN(G1351GAT) );
  XOR2_X1 U331 ( .A(KEYINPUT75), .B(KEYINPUT11), .Z(n294) );
  XNOR2_X1 U332 ( .A(G134GAT), .B(KEYINPUT74), .ZN(n293) );
  XNOR2_X1 U333 ( .A(n294), .B(n293), .ZN(n302) );
  XNOR2_X1 U334 ( .A(G36GAT), .B(G190GAT), .ZN(n296) );
  INV_X1 U335 ( .A(n296), .ZN(n383) );
  XNOR2_X1 U336 ( .A(G99GAT), .B(G85GAT), .ZN(n295) );
  NAND2_X1 U337 ( .A1(n383), .A2(n295), .ZN(n298) );
  INV_X1 U338 ( .A(n295), .ZN(n333) );
  NAND2_X1 U339 ( .A1(n296), .A2(n333), .ZN(n297) );
  NAND2_X1 U340 ( .A1(n298), .A2(n297), .ZN(n300) );
  NAND2_X1 U341 ( .A1(G232GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U342 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U343 ( .A(n302), .B(n301), .Z(n307) );
  XOR2_X1 U344 ( .A(G50GAT), .B(G162GAT), .Z(n434) );
  XOR2_X1 U345 ( .A(KEYINPUT9), .B(KEYINPUT76), .Z(n304) );
  XNOR2_X1 U346 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n303) );
  XNOR2_X1 U347 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U348 ( .A(n434), .B(n305), .ZN(n306) );
  XNOR2_X1 U349 ( .A(n307), .B(n306), .ZN(n309) );
  INV_X1 U350 ( .A(G92GAT), .ZN(n308) );
  XNOR2_X1 U351 ( .A(n309), .B(n308), .ZN(n313) );
  XOR2_X1 U352 ( .A(G29GAT), .B(G43GAT), .Z(n311) );
  XNOR2_X1 U353 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n310) );
  XNOR2_X1 U354 ( .A(n311), .B(n310), .ZN(n323) );
  XNOR2_X1 U355 ( .A(n323), .B(G106GAT), .ZN(n312) );
  XNOR2_X1 U356 ( .A(n313), .B(n312), .ZN(n549) );
  INV_X1 U357 ( .A(n549), .ZN(n561) );
  INV_X1 U358 ( .A(KEYINPUT54), .ZN(n399) );
  XOR2_X1 U359 ( .A(KEYINPUT70), .B(KEYINPUT30), .Z(n315) );
  XNOR2_X1 U360 ( .A(G197GAT), .B(KEYINPUT29), .ZN(n314) );
  XNOR2_X1 U361 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U362 ( .A(KEYINPUT68), .B(KEYINPUT67), .Z(n317) );
  XNOR2_X1 U363 ( .A(KEYINPUT69), .B(KEYINPUT66), .ZN(n316) );
  XNOR2_X1 U364 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U365 ( .A(n319), .B(n318), .ZN(n330) );
  XOR2_X1 U366 ( .A(G50GAT), .B(G36GAT), .Z(n321) );
  XOR2_X1 U367 ( .A(G141GAT), .B(G22GAT), .Z(n435) );
  XOR2_X1 U368 ( .A(G113GAT), .B(G1GAT), .Z(n412) );
  XNOR2_X1 U369 ( .A(n435), .B(n412), .ZN(n320) );
  XNOR2_X1 U370 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U371 ( .A(n322), .B(G15GAT), .Z(n328) );
  XOR2_X1 U372 ( .A(n323), .B(G8GAT), .Z(n325) );
  NAND2_X1 U373 ( .A1(G229GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U374 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U375 ( .A(G169GAT), .B(n326), .ZN(n327) );
  XNOR2_X1 U376 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U377 ( .A(n330), .B(n329), .ZN(n577) );
  INV_X1 U378 ( .A(n577), .ZN(n538) );
  XNOR2_X1 U379 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n345) );
  XOR2_X1 U380 ( .A(G78GAT), .B(G148GAT), .Z(n332) );
  XNOR2_X1 U381 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n331) );
  XNOR2_X1 U382 ( .A(n332), .B(n331), .ZN(n426) );
  XNOR2_X1 U383 ( .A(n333), .B(n292), .ZN(n334) );
  XOR2_X1 U384 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n336) );
  XNOR2_X1 U385 ( .A(KEYINPUT73), .B(KEYINPUT33), .ZN(n335) );
  XNOR2_X1 U386 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U387 ( .A(n338), .B(n337), .Z(n344) );
  XOR2_X1 U388 ( .A(KEYINPUT72), .B(G64GAT), .Z(n340) );
  XNOR2_X1 U389 ( .A(G176GAT), .B(G92GAT), .ZN(n339) );
  XNOR2_X1 U390 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U391 ( .A(G204GAT), .B(n341), .Z(n394) );
  XOR2_X1 U392 ( .A(G120GAT), .B(G71GAT), .Z(n444) );
  XOR2_X1 U393 ( .A(G57GAT), .B(KEYINPUT13), .Z(n362) );
  XNOR2_X1 U394 ( .A(n444), .B(n362), .ZN(n342) );
  XOR2_X1 U395 ( .A(n345), .B(n582), .Z(n565) );
  INV_X1 U396 ( .A(n565), .ZN(n540) );
  NAND2_X1 U397 ( .A1(n538), .A2(n540), .ZN(n346) );
  XNOR2_X1 U398 ( .A(KEYINPUT46), .B(n346), .ZN(n367) );
  XOR2_X1 U399 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n348) );
  XNOR2_X1 U400 ( .A(KEYINPUT82), .B(KEYINPUT12), .ZN(n347) );
  XNOR2_X1 U401 ( .A(n348), .B(n347), .ZN(n366) );
  XOR2_X1 U402 ( .A(G78GAT), .B(G155GAT), .Z(n350) );
  XNOR2_X1 U403 ( .A(G22GAT), .B(G71GAT), .ZN(n349) );
  XNOR2_X1 U404 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U405 ( .A(KEYINPUT81), .B(G64GAT), .Z(n352) );
  XNOR2_X1 U406 ( .A(G1GAT), .B(G211GAT), .ZN(n351) );
  XNOR2_X1 U407 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U408 ( .A(n354), .B(n353), .Z(n359) );
  XOR2_X1 U409 ( .A(KEYINPUT79), .B(KEYINPUT78), .Z(n356) );
  NAND2_X1 U410 ( .A1(G231GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U412 ( .A(KEYINPUT80), .B(n357), .ZN(n358) );
  XNOR2_X1 U413 ( .A(n359), .B(n358), .ZN(n361) );
  XNOR2_X1 U414 ( .A(G8GAT), .B(G183GAT), .ZN(n360) );
  XNOR2_X1 U415 ( .A(n360), .B(KEYINPUT77), .ZN(n386) );
  XOR2_X1 U416 ( .A(n361), .B(n386), .Z(n364) );
  XOR2_X1 U417 ( .A(G15GAT), .B(G127GAT), .Z(n448) );
  XNOR2_X1 U418 ( .A(n448), .B(n362), .ZN(n363) );
  XNOR2_X1 U419 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U420 ( .A(n366), .B(n365), .Z(n585) );
  NAND2_X1 U421 ( .A1(n367), .A2(n585), .ZN(n368) );
  NOR2_X1 U422 ( .A1(n368), .A2(n549), .ZN(n370) );
  XNOR2_X1 U423 ( .A(KEYINPUT111), .B(KEYINPUT47), .ZN(n369) );
  XNOR2_X1 U424 ( .A(n370), .B(n369), .ZN(n376) );
  INV_X1 U425 ( .A(n582), .ZN(n464) );
  XOR2_X1 U426 ( .A(n549), .B(KEYINPUT36), .Z(n590) );
  NOR2_X1 U427 ( .A1(n585), .A2(n590), .ZN(n371) );
  XOR2_X1 U428 ( .A(KEYINPUT45), .B(n371), .Z(n372) );
  NOR2_X1 U429 ( .A1(n464), .A2(n372), .ZN(n373) );
  XOR2_X1 U430 ( .A(KEYINPUT112), .B(n373), .Z(n374) );
  NOR2_X1 U431 ( .A1(n538), .A2(n374), .ZN(n375) );
  NOR2_X1 U432 ( .A1(n376), .A2(n375), .ZN(n378) );
  XNOR2_X1 U433 ( .A(KEYINPUT113), .B(KEYINPUT48), .ZN(n377) );
  XNOR2_X1 U434 ( .A(n378), .B(n377), .ZN(n531) );
  XOR2_X1 U435 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n385) );
  XNOR2_X1 U436 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n379) );
  XNOR2_X1 U437 ( .A(n379), .B(KEYINPUT85), .ZN(n380) );
  XOR2_X1 U438 ( .A(n380), .B(KEYINPUT86), .Z(n382) );
  XNOR2_X1 U439 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n381) );
  XNOR2_X1 U440 ( .A(n382), .B(n381), .ZN(n456) );
  XNOR2_X1 U441 ( .A(n456), .B(n383), .ZN(n384) );
  XNOR2_X1 U442 ( .A(n385), .B(n384), .ZN(n390) );
  XOR2_X1 U443 ( .A(n386), .B(KEYINPUT96), .Z(n388) );
  NAND2_X1 U444 ( .A1(G226GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U445 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U446 ( .A(n390), .B(n389), .Z(n397) );
  XOR2_X1 U447 ( .A(KEYINPUT90), .B(G218GAT), .Z(n392) );
  XNOR2_X1 U448 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n391) );
  XNOR2_X1 U449 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U450 ( .A(G197GAT), .B(n393), .ZN(n438) );
  INV_X1 U451 ( .A(n438), .ZN(n395) );
  XNOR2_X1 U452 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U453 ( .A(n397), .B(n396), .ZN(n485) );
  NAND2_X1 U454 ( .A1(n531), .A2(n485), .ZN(n398) );
  XNOR2_X1 U455 ( .A(n399), .B(n398), .ZN(n421) );
  XOR2_X1 U456 ( .A(KEYINPUT93), .B(KEYINPUT1), .Z(n401) );
  XNOR2_X1 U457 ( .A(KEYINPUT95), .B(KEYINPUT6), .ZN(n400) );
  XNOR2_X1 U458 ( .A(n401), .B(n400), .ZN(n420) );
  XOR2_X1 U459 ( .A(G162GAT), .B(G120GAT), .Z(n403) );
  XNOR2_X1 U460 ( .A(G141GAT), .B(G127GAT), .ZN(n402) );
  XNOR2_X1 U461 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U462 ( .A(KEYINPUT94), .B(KEYINPUT5), .Z(n405) );
  XNOR2_X1 U463 ( .A(G148GAT), .B(G57GAT), .ZN(n404) );
  XNOR2_X1 U464 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U465 ( .A(n407), .B(n406), .Z(n418) );
  XNOR2_X1 U466 ( .A(G134GAT), .B(KEYINPUT83), .ZN(n408) );
  XNOR2_X1 U467 ( .A(n408), .B(KEYINPUT0), .ZN(n447) );
  XOR2_X1 U468 ( .A(KEYINPUT4), .B(n447), .Z(n410) );
  NAND2_X1 U469 ( .A1(G225GAT), .A2(G233GAT), .ZN(n409) );
  XNOR2_X1 U470 ( .A(n410), .B(n409), .ZN(n416) );
  XNOR2_X1 U471 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n411) );
  XNOR2_X1 U472 ( .A(n411), .B(KEYINPUT2), .ZN(n427) );
  XOR2_X1 U473 ( .A(G85GAT), .B(n427), .Z(n414) );
  XNOR2_X1 U474 ( .A(G29GAT), .B(n412), .ZN(n413) );
  XNOR2_X1 U475 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U476 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U477 ( .A(n418), .B(n417), .ZN(n419) );
  NAND2_X1 U478 ( .A1(n421), .A2(n533), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n422), .B(KEYINPUT65), .ZN(n576) );
  XOR2_X1 U480 ( .A(KEYINPUT24), .B(KEYINPUT92), .Z(n424) );
  NAND2_X1 U481 ( .A1(G228GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U482 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U483 ( .A(n425), .B(KEYINPUT91), .Z(n429) );
  XNOR2_X1 U484 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U485 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U486 ( .A(G204GAT), .B(KEYINPUT23), .Z(n431) );
  XNOR2_X1 U487 ( .A(KEYINPUT22), .B(KEYINPUT89), .ZN(n430) );
  XNOR2_X1 U488 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U489 ( .A(n433), .B(n432), .Z(n437) );
  XNOR2_X1 U490 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n439) );
  XNOR2_X1 U492 ( .A(n439), .B(n438), .ZN(n471) );
  NAND2_X1 U493 ( .A1(n576), .A2(n471), .ZN(n440) );
  XNOR2_X1 U494 ( .A(n440), .B(KEYINPUT55), .ZN(n459) );
  XOR2_X1 U495 ( .A(G183GAT), .B(KEYINPUT87), .Z(n442) );
  XNOR2_X1 U496 ( .A(G99GAT), .B(KEYINPUT88), .ZN(n441) );
  XNOR2_X1 U497 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U498 ( .A(n443), .B(G190GAT), .Z(n446) );
  XNOR2_X1 U499 ( .A(G43GAT), .B(n444), .ZN(n445) );
  XNOR2_X1 U500 ( .A(n446), .B(n445), .ZN(n452) );
  XOR2_X1 U501 ( .A(n448), .B(n447), .Z(n450) );
  NAND2_X1 U502 ( .A1(G227GAT), .A2(G233GAT), .ZN(n449) );
  XNOR2_X1 U503 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U504 ( .A(n452), .B(n451), .Z(n458) );
  XOR2_X1 U505 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n454) );
  XNOR2_X1 U506 ( .A(G113GAT), .B(G176GAT), .ZN(n453) );
  XNOR2_X1 U507 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U508 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U509 ( .A(n458), .B(n457), .ZN(n534) );
  NAND2_X1 U510 ( .A1(n459), .A2(n534), .ZN(n571) );
  NOR2_X1 U511 ( .A1(n561), .A2(n571), .ZN(n463) );
  XNOR2_X1 U512 ( .A(KEYINPUT122), .B(KEYINPUT58), .ZN(n461) );
  INV_X1 U513 ( .A(G190GAT), .ZN(n460) );
  NOR2_X1 U514 ( .A1(n577), .A2(n464), .ZN(n495) );
  NOR2_X1 U515 ( .A1(n549), .A2(n585), .ZN(n465) );
  XNOR2_X1 U516 ( .A(KEYINPUT16), .B(n465), .ZN(n480) );
  NAND2_X1 U517 ( .A1(n534), .A2(n485), .ZN(n466) );
  XNOR2_X1 U518 ( .A(KEYINPUT100), .B(n466), .ZN(n467) );
  NAND2_X1 U519 ( .A1(n467), .A2(n471), .ZN(n468) );
  XNOR2_X1 U520 ( .A(KEYINPUT25), .B(n468), .ZN(n469) );
  NAND2_X1 U521 ( .A1(n533), .A2(n469), .ZN(n479) );
  XOR2_X1 U522 ( .A(n471), .B(KEYINPUT28), .Z(n537) );
  NOR2_X1 U523 ( .A1(n534), .A2(n537), .ZN(n470) );
  NOR2_X1 U524 ( .A1(n533), .A2(n470), .ZN(n476) );
  NOR2_X1 U525 ( .A1(n534), .A2(n471), .ZN(n472) );
  XOR2_X1 U526 ( .A(KEYINPUT26), .B(n472), .Z(n473) );
  XNOR2_X1 U527 ( .A(KEYINPUT99), .B(n473), .ZN(n575) );
  INV_X1 U528 ( .A(n533), .ZN(n474) );
  NOR2_X1 U529 ( .A1(n575), .A2(n474), .ZN(n475) );
  NOR2_X1 U530 ( .A1(n476), .A2(n475), .ZN(n477) );
  XNOR2_X1 U531 ( .A(n485), .B(KEYINPUT27), .ZN(n530) );
  NAND2_X1 U532 ( .A1(n477), .A2(n530), .ZN(n478) );
  NAND2_X1 U533 ( .A1(n479), .A2(n478), .ZN(n491) );
  NAND2_X1 U534 ( .A1(n480), .A2(n491), .ZN(n481) );
  XNOR2_X1 U535 ( .A(n481), .B(KEYINPUT101), .ZN(n507) );
  NAND2_X1 U536 ( .A1(n495), .A2(n507), .ZN(n489) );
  NOR2_X1 U537 ( .A1(n533), .A2(n489), .ZN(n483) );
  XNOR2_X1 U538 ( .A(KEYINPUT34), .B(KEYINPUT102), .ZN(n482) );
  XNOR2_X1 U539 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U540 ( .A(G1GAT), .B(n484), .Z(G1324GAT) );
  INV_X1 U541 ( .A(n485), .ZN(n520) );
  NOR2_X1 U542 ( .A1(n520), .A2(n489), .ZN(n486) );
  XOR2_X1 U543 ( .A(G8GAT), .B(n486), .Z(G1325GAT) );
  INV_X1 U544 ( .A(n534), .ZN(n522) );
  NOR2_X1 U545 ( .A1(n522), .A2(n489), .ZN(n488) );
  XNOR2_X1 U546 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n488), .B(n487), .ZN(G1326GAT) );
  INV_X1 U548 ( .A(n537), .ZN(n526) );
  NOR2_X1 U549 ( .A1(n526), .A2(n489), .ZN(n490) );
  XOR2_X1 U550 ( .A(G22GAT), .B(n490), .Z(G1327GAT) );
  XNOR2_X1 U551 ( .A(KEYINPUT38), .B(KEYINPUT104), .ZN(n497) );
  NAND2_X1 U552 ( .A1(n585), .A2(n491), .ZN(n492) );
  NOR2_X1 U553 ( .A1(n590), .A2(n492), .ZN(n494) );
  XNOR2_X1 U554 ( .A(KEYINPUT103), .B(KEYINPUT37), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(n517) );
  NAND2_X1 U556 ( .A1(n517), .A2(n495), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n497), .B(n496), .ZN(n504) );
  NOR2_X1 U558 ( .A1(n533), .A2(n504), .ZN(n499) );
  XNOR2_X1 U559 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n499), .B(n498), .ZN(G1328GAT) );
  NOR2_X1 U561 ( .A1(n520), .A2(n504), .ZN(n500) );
  XOR2_X1 U562 ( .A(G36GAT), .B(n500), .Z(G1329GAT) );
  NOR2_X1 U563 ( .A1(n522), .A2(n504), .ZN(n502) );
  XNOR2_X1 U564 ( .A(KEYINPUT105), .B(KEYINPUT40), .ZN(n501) );
  XNOR2_X1 U565 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U566 ( .A(G43GAT), .B(n503), .ZN(G1330GAT) );
  NOR2_X1 U567 ( .A1(n526), .A2(n504), .ZN(n505) );
  XOR2_X1 U568 ( .A(G50GAT), .B(n505), .Z(n506) );
  XNOR2_X1 U569 ( .A(KEYINPUT106), .B(n506), .ZN(G1331GAT) );
  NOR2_X1 U570 ( .A1(n565), .A2(n538), .ZN(n516) );
  NAND2_X1 U571 ( .A1(n507), .A2(n516), .ZN(n512) );
  NOR2_X1 U572 ( .A1(n533), .A2(n512), .ZN(n508) );
  XOR2_X1 U573 ( .A(G57GAT), .B(n508), .Z(n509) );
  XNOR2_X1 U574 ( .A(KEYINPUT42), .B(n509), .ZN(G1332GAT) );
  NOR2_X1 U575 ( .A1(n520), .A2(n512), .ZN(n510) );
  XOR2_X1 U576 ( .A(G64GAT), .B(n510), .Z(G1333GAT) );
  NOR2_X1 U577 ( .A1(n522), .A2(n512), .ZN(n511) );
  XOR2_X1 U578 ( .A(G71GAT), .B(n511), .Z(G1334GAT) );
  NOR2_X1 U579 ( .A1(n526), .A2(n512), .ZN(n514) );
  XNOR2_X1 U580 ( .A(KEYINPUT107), .B(KEYINPUT43), .ZN(n513) );
  XNOR2_X1 U581 ( .A(n514), .B(n513), .ZN(n515) );
  XOR2_X1 U582 ( .A(G78GAT), .B(n515), .Z(G1335GAT) );
  NAND2_X1 U583 ( .A1(n517), .A2(n516), .ZN(n525) );
  NOR2_X1 U584 ( .A1(n533), .A2(n525), .ZN(n518) );
  XOR2_X1 U585 ( .A(G85GAT), .B(n518), .Z(n519) );
  XNOR2_X1 U586 ( .A(KEYINPUT108), .B(n519), .ZN(G1336GAT) );
  NOR2_X1 U587 ( .A1(n520), .A2(n525), .ZN(n521) );
  XOR2_X1 U588 ( .A(G92GAT), .B(n521), .Z(G1337GAT) );
  NOR2_X1 U589 ( .A1(n522), .A2(n525), .ZN(n524) );
  XNOR2_X1 U590 ( .A(G99GAT), .B(KEYINPUT109), .ZN(n523) );
  XNOR2_X1 U591 ( .A(n524), .B(n523), .ZN(G1338GAT) );
  NOR2_X1 U592 ( .A1(n526), .A2(n525), .ZN(n528) );
  XNOR2_X1 U593 ( .A(KEYINPUT110), .B(KEYINPUT44), .ZN(n527) );
  XNOR2_X1 U594 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U595 ( .A(G106GAT), .B(n529), .Z(G1339GAT) );
  NAND2_X1 U596 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U597 ( .A1(n533), .A2(n532), .ZN(n553) );
  NAND2_X1 U598 ( .A1(n534), .A2(n553), .ZN(n535) );
  XNOR2_X1 U599 ( .A(KEYINPUT114), .B(n535), .ZN(n536) );
  NOR2_X1 U600 ( .A1(n537), .A2(n536), .ZN(n550) );
  NAND2_X1 U601 ( .A1(n538), .A2(n550), .ZN(n539) );
  XNOR2_X1 U602 ( .A(n539), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n542) );
  NAND2_X1 U604 ( .A1(n550), .A2(n540), .ZN(n541) );
  XNOR2_X1 U605 ( .A(n542), .B(n541), .ZN(n544) );
  XOR2_X1 U606 ( .A(G120GAT), .B(KEYINPUT115), .Z(n543) );
  XNOR2_X1 U607 ( .A(n544), .B(n543), .ZN(G1341GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n547) );
  INV_X1 U609 ( .A(n585), .ZN(n545) );
  NAND2_X1 U610 ( .A1(n550), .A2(n545), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U612 ( .A(G127GAT), .B(n548), .ZN(G1342GAT) );
  XOR2_X1 U613 ( .A(G134GAT), .B(KEYINPUT51), .Z(n552) );
  NAND2_X1 U614 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U615 ( .A(n552), .B(n551), .ZN(G1343GAT) );
  NAND2_X1 U616 ( .A1(n553), .A2(n575), .ZN(n560) );
  NOR2_X1 U617 ( .A1(n577), .A2(n560), .ZN(n554) );
  XOR2_X1 U618 ( .A(G141GAT), .B(n554), .Z(G1344GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT118), .B(KEYINPUT52), .Z(n556) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n556), .B(n555), .ZN(n558) );
  NOR2_X1 U622 ( .A1(n565), .A2(n560), .ZN(n557) );
  XOR2_X1 U623 ( .A(n558), .B(n557), .Z(G1345GAT) );
  NOR2_X1 U624 ( .A1(n585), .A2(n560), .ZN(n559) );
  XOR2_X1 U625 ( .A(G155GAT), .B(n559), .Z(G1346GAT) );
  NOR2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U627 ( .A(G162GAT), .B(n562), .Z(G1347GAT) );
  NOR2_X1 U628 ( .A1(n577), .A2(n571), .ZN(n564) );
  XNOR2_X1 U629 ( .A(G169GAT), .B(KEYINPUT119), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(G1348GAT) );
  NOR2_X1 U631 ( .A1(n565), .A2(n571), .ZN(n570) );
  XOR2_X1 U632 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n567) );
  XNOR2_X1 U633 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U635 ( .A(KEYINPUT56), .B(n568), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(G1349GAT) );
  NOR2_X1 U637 ( .A1(n585), .A2(n571), .ZN(n572) );
  XOR2_X1 U638 ( .A(G183GAT), .B(n572), .Z(G1350GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT125), .B(KEYINPUT124), .Z(n574) );
  XNOR2_X1 U640 ( .A(KEYINPUT123), .B(KEYINPUT60), .ZN(n573) );
  XNOR2_X1 U641 ( .A(n574), .B(n573), .ZN(n581) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n589) );
  NOR2_X1 U643 ( .A1(n577), .A2(n589), .ZN(n579) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n580) );
  XOR2_X1 U646 ( .A(n581), .B(n580), .Z(G1352GAT) );
  NOR2_X1 U647 ( .A1(n582), .A2(n589), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  NOR2_X1 U650 ( .A1(n585), .A2(n589), .ZN(n586) );
  XOR2_X1 U651 ( .A(G211GAT), .B(n586), .Z(G1354GAT) );
  XOR2_X1 U652 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n588) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n587) );
  XNOR2_X1 U654 ( .A(n588), .B(n587), .ZN(n592) );
  NOR2_X1 U655 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U656 ( .A(n592), .B(n591), .Z(G1355GAT) );
endmodule

