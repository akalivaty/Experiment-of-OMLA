

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603;

  INV_X1 U328 ( .A(n574), .ZN(n586) );
  OR2_X1 U329 ( .A1(n297), .A2(n587), .ZN(n578) );
  AND2_X1 U330 ( .A1(n590), .A2(n577), .ZN(n470) );
  XNOR2_X1 U331 ( .A(KEYINPUT93), .B(KEYINPUT27), .ZN(n340) );
  XNOR2_X1 U332 ( .A(n327), .B(n326), .ZN(n353) );
  NOR2_X2 U333 ( .A1(n559), .A2(n488), .ZN(n600) );
  XNOR2_X1 U334 ( .A(n403), .B(n402), .ZN(n599) );
  XNOR2_X1 U335 ( .A(n460), .B(KEYINPUT38), .ZN(n461) );
  NAND2_X1 U336 ( .A1(n586), .A2(n585), .ZN(n296) );
  NAND2_X1 U337 ( .A1(n586), .A2(n577), .ZN(n297) );
  AND2_X1 U338 ( .A1(G231GAT), .A2(G233GAT), .ZN(n298) );
  INV_X1 U339 ( .A(KEYINPUT45), .ZN(n475) );
  XNOR2_X1 U340 ( .A(n475), .B(KEYINPUT112), .ZN(n476) );
  XNOR2_X1 U341 ( .A(n477), .B(n476), .ZN(n478) );
  INV_X1 U342 ( .A(n453), .ZN(n454) );
  INV_X1 U343 ( .A(G211GAT), .ZN(n324) );
  XNOR2_X1 U344 ( .A(n393), .B(n298), .ZN(n394) );
  XNOR2_X1 U345 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U346 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U347 ( .A(n395), .B(n394), .ZN(n401) );
  XNOR2_X1 U348 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U349 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U350 ( .A(n337), .B(n336), .ZN(n338) );
  INV_X1 U351 ( .A(G218GAT), .ZN(n491) );
  XOR2_X1 U352 ( .A(n595), .B(n467), .Z(n577) );
  XNOR2_X1 U353 ( .A(n462), .B(n461), .ZN(n515) );
  XNOR2_X1 U354 ( .A(n491), .B(KEYINPUT62), .ZN(n492) );
  XNOR2_X1 U355 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U356 ( .A(n493), .B(n492), .ZN(G1355GAT) );
  XNOR2_X1 U357 ( .A(n466), .B(n465), .ZN(G1328GAT) );
  XOR2_X1 U358 ( .A(KEYINPUT1), .B(G57GAT), .Z(n300) );
  XNOR2_X1 U359 ( .A(G1GAT), .B(G148GAT), .ZN(n299) );
  XNOR2_X1 U360 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U361 ( .A(KEYINPUT4), .B(KEYINPUT88), .Z(n302) );
  XNOR2_X1 U362 ( .A(KEYINPUT91), .B(KEYINPUT90), .ZN(n301) );
  XNOR2_X1 U363 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U364 ( .A(n304), .B(n303), .Z(n309) );
  XOR2_X1 U365 ( .A(KEYINPUT89), .B(KEYINPUT6), .Z(n306) );
  NAND2_X1 U366 ( .A1(G225GAT), .A2(G233GAT), .ZN(n305) );
  XNOR2_X1 U367 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U368 ( .A(KEYINPUT5), .B(n307), .ZN(n308) );
  XNOR2_X1 U369 ( .A(n309), .B(n308), .ZN(n313) );
  XOR2_X1 U370 ( .A(G85GAT), .B(G162GAT), .Z(n311) );
  XNOR2_X1 U371 ( .A(G29GAT), .B(G120GAT), .ZN(n310) );
  XNOR2_X1 U372 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U373 ( .A(n313), .B(n312), .Z(n321) );
  XOR2_X1 U374 ( .A(G127GAT), .B(KEYINPUT0), .Z(n315) );
  XNOR2_X1 U375 ( .A(G113GAT), .B(G134GAT), .ZN(n314) );
  XNOR2_X1 U376 ( .A(n315), .B(n314), .ZN(n365) );
  XNOR2_X1 U377 ( .A(KEYINPUT86), .B(KEYINPUT85), .ZN(n316) );
  XNOR2_X1 U378 ( .A(n316), .B(KEYINPUT3), .ZN(n317) );
  XOR2_X1 U379 ( .A(n317), .B(KEYINPUT2), .Z(n319) );
  XNOR2_X1 U380 ( .A(G141GAT), .B(G155GAT), .ZN(n318) );
  XNOR2_X1 U381 ( .A(n319), .B(n318), .ZN(n349) );
  XNOR2_X1 U382 ( .A(n365), .B(n349), .ZN(n320) );
  XNOR2_X1 U383 ( .A(n321), .B(n320), .ZN(n543) );
  XOR2_X1 U384 ( .A(G169GAT), .B(G8GAT), .Z(n428) );
  XOR2_X1 U385 ( .A(G176GAT), .B(G64GAT), .Z(n451) );
  XNOR2_X1 U386 ( .A(n428), .B(n451), .ZN(n339) );
  XOR2_X1 U387 ( .A(G36GAT), .B(G190GAT), .Z(n407) );
  XOR2_X1 U388 ( .A(KEYINPUT21), .B(KEYINPUT83), .Z(n323) );
  XNOR2_X1 U389 ( .A(G218GAT), .B(KEYINPUT84), .ZN(n322) );
  XNOR2_X1 U390 ( .A(n323), .B(n322), .ZN(n327) );
  XNOR2_X1 U391 ( .A(G197GAT), .B(G204GAT), .ZN(n325) );
  XNOR2_X1 U392 ( .A(n407), .B(n353), .ZN(n329) );
  AND2_X1 U393 ( .A1(G226GAT), .A2(G233GAT), .ZN(n328) );
  NAND2_X1 U394 ( .A1(n329), .A2(n328), .ZN(n331) );
  OR2_X1 U395 ( .A1(n329), .A2(n328), .ZN(n330) );
  NAND2_X1 U396 ( .A1(n331), .A2(n330), .ZN(n337) );
  XOR2_X1 U397 ( .A(G183GAT), .B(KEYINPUT17), .Z(n333) );
  XNOR2_X1 U398 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n332) );
  XNOR2_X1 U399 ( .A(n333), .B(n332), .ZN(n363) );
  XNOR2_X1 U400 ( .A(n363), .B(G92GAT), .ZN(n335) );
  INV_X1 U401 ( .A(KEYINPUT92), .ZN(n334) );
  XNOR2_X1 U402 ( .A(n339), .B(n338), .ZN(n513) );
  XNOR2_X1 U403 ( .A(n513), .B(n340), .ZN(n545) );
  INV_X1 U404 ( .A(n545), .ZN(n376) );
  XNOR2_X1 U405 ( .A(KEYINPUT28), .B(KEYINPUT67), .ZN(n354) );
  XOR2_X1 U406 ( .A(KEYINPUT87), .B(KEYINPUT23), .Z(n342) );
  XNOR2_X1 U407 ( .A(KEYINPUT22), .B(KEYINPUT24), .ZN(n341) );
  XNOR2_X1 U408 ( .A(n342), .B(n341), .ZN(n344) );
  XNOR2_X1 U409 ( .A(G106GAT), .B(G78GAT), .ZN(n343) );
  XNOR2_X1 U410 ( .A(n343), .B(G148GAT), .ZN(n448) );
  XOR2_X1 U411 ( .A(n344), .B(n448), .Z(n351) );
  XNOR2_X1 U412 ( .A(G50GAT), .B(KEYINPUT76), .ZN(n345) );
  XNOR2_X1 U413 ( .A(n345), .B(G162GAT), .ZN(n416) );
  XOR2_X1 U414 ( .A(n416), .B(G22GAT), .Z(n347) );
  NAND2_X1 U415 ( .A1(G228GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U416 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U417 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U418 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U419 ( .A(n353), .B(n352), .ZN(n571) );
  XNOR2_X1 U420 ( .A(n354), .B(n571), .ZN(n548) );
  NOR2_X1 U421 ( .A1(n376), .A2(n548), .ZN(n356) );
  INV_X1 U422 ( .A(n543), .ZN(n531) );
  AND2_X1 U423 ( .A1(n531), .A2(KEYINPUT94), .ZN(n355) );
  AND2_X1 U424 ( .A1(n356), .A2(n355), .ZN(n358) );
  NOR2_X1 U425 ( .A1(KEYINPUT94), .A2(n356), .ZN(n357) );
  NOR2_X1 U426 ( .A1(n358), .A2(n357), .ZN(n373) );
  XOR2_X1 U427 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n360) );
  XNOR2_X1 U428 ( .A(G99GAT), .B(KEYINPUT81), .ZN(n359) );
  XNOR2_X1 U429 ( .A(n360), .B(n359), .ZN(n372) );
  XOR2_X1 U430 ( .A(G176GAT), .B(G15GAT), .Z(n362) );
  NAND2_X1 U431 ( .A1(G227GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U432 ( .A(n362), .B(n361), .ZN(n364) );
  XOR2_X1 U433 ( .A(n364), .B(n363), .Z(n367) );
  XNOR2_X1 U434 ( .A(G169GAT), .B(n365), .ZN(n366) );
  XNOR2_X1 U435 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U436 ( .A(G120GAT), .B(G71GAT), .Z(n452) );
  XOR2_X1 U437 ( .A(n368), .B(n452), .Z(n370) );
  XNOR2_X1 U438 ( .A(G43GAT), .B(G190GAT), .ZN(n369) );
  XNOR2_X1 U439 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U440 ( .A(n372), .B(n371), .ZN(n574) );
  NOR2_X1 U441 ( .A1(n373), .A2(n586), .ZN(n387) );
  NOR2_X1 U442 ( .A1(n586), .A2(n571), .ZN(n375) );
  XNOR2_X1 U443 ( .A(KEYINPUT26), .B(KEYINPUT95), .ZN(n374) );
  XNOR2_X1 U444 ( .A(n375), .B(n374), .ZN(n559) );
  NOR2_X1 U445 ( .A1(n376), .A2(n559), .ZN(n377) );
  XNOR2_X1 U446 ( .A(n377), .B(KEYINPUT96), .ZN(n384) );
  INV_X1 U447 ( .A(n513), .ZN(n533) );
  NAND2_X1 U448 ( .A1(n533), .A2(n586), .ZN(n378) );
  NAND2_X1 U449 ( .A1(n378), .A2(n571), .ZN(n379) );
  XNOR2_X1 U450 ( .A(n379), .B(KEYINPUT97), .ZN(n380) );
  XNOR2_X1 U451 ( .A(n380), .B(KEYINPUT25), .ZN(n382) );
  OR2_X1 U452 ( .A1(n586), .A2(KEYINPUT94), .ZN(n381) );
  NAND2_X1 U453 ( .A1(n382), .A2(n381), .ZN(n383) );
  NOR2_X1 U454 ( .A1(n384), .A2(n383), .ZN(n385) );
  NOR2_X1 U455 ( .A1(n385), .A2(n531), .ZN(n386) );
  NOR2_X1 U456 ( .A1(n387), .A2(n386), .ZN(n499) );
  XOR2_X1 U457 ( .A(G64GAT), .B(G155GAT), .Z(n389) );
  XNOR2_X1 U458 ( .A(G8GAT), .B(G211GAT), .ZN(n388) );
  XNOR2_X1 U459 ( .A(n389), .B(n388), .ZN(n403) );
  XNOR2_X1 U460 ( .A(G15GAT), .B(G22GAT), .ZN(n390) );
  XNOR2_X1 U461 ( .A(n390), .B(G1GAT), .ZN(n427) );
  XOR2_X1 U462 ( .A(n427), .B(KEYINPUT80), .Z(n395) );
  XOR2_X1 U463 ( .A(G78GAT), .B(G71GAT), .Z(n392) );
  XNOR2_X1 U464 ( .A(G127GAT), .B(G183GAT), .ZN(n391) );
  XNOR2_X1 U465 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U466 ( .A(G57GAT), .B(KEYINPUT71), .ZN(n396) );
  XNOR2_X1 U467 ( .A(n396), .B(KEYINPUT13), .ZN(n453) );
  XOR2_X1 U468 ( .A(KEYINPUT15), .B(KEYINPUT79), .Z(n398) );
  XNOR2_X1 U469 ( .A(KEYINPUT12), .B(KEYINPUT14), .ZN(n397) );
  XNOR2_X1 U470 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U471 ( .A(n453), .B(n399), .ZN(n400) );
  XNOR2_X1 U472 ( .A(n401), .B(n400), .ZN(n402) );
  NOR2_X1 U473 ( .A1(n499), .A2(n599), .ZN(n404) );
  XNOR2_X1 U474 ( .A(n404), .B(KEYINPUT101), .ZN(n425) );
  XOR2_X1 U475 ( .A(KEYINPUT10), .B(KEYINPUT66), .Z(n406) );
  XNOR2_X1 U476 ( .A(G218GAT), .B(KEYINPUT78), .ZN(n405) );
  XNOR2_X1 U477 ( .A(n406), .B(n405), .ZN(n408) );
  XOR2_X1 U478 ( .A(n408), .B(n407), .Z(n410) );
  XNOR2_X1 U479 ( .A(G134GAT), .B(G106GAT), .ZN(n409) );
  XNOR2_X1 U480 ( .A(n410), .B(n409), .ZN(n420) );
  XOR2_X1 U481 ( .A(KEYINPUT9), .B(KEYINPUT77), .Z(n412) );
  NAND2_X1 U482 ( .A1(G232GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U483 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U484 ( .A(n413), .B(KEYINPUT11), .Z(n418) );
  XOR2_X1 U485 ( .A(G92GAT), .B(KEYINPUT73), .Z(n415) );
  XNOR2_X1 U486 ( .A(G99GAT), .B(G85GAT), .ZN(n414) );
  XNOR2_X1 U487 ( .A(n415), .B(n414), .ZN(n447) );
  XNOR2_X1 U488 ( .A(n416), .B(n447), .ZN(n417) );
  XNOR2_X1 U489 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U490 ( .A(n420), .B(n419), .ZN(n424) );
  XOR2_X1 U491 ( .A(KEYINPUT69), .B(KEYINPUT7), .Z(n422) );
  XNOR2_X1 U492 ( .A(G43GAT), .B(G29GAT), .ZN(n421) );
  XNOR2_X1 U493 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U494 ( .A(KEYINPUT8), .B(n423), .ZN(n440) );
  XNOR2_X1 U495 ( .A(n424), .B(n440), .ZN(n585) );
  XOR2_X1 U496 ( .A(n585), .B(KEYINPUT36), .Z(n490) );
  NOR2_X1 U497 ( .A1(n425), .A2(n490), .ZN(n426) );
  XNOR2_X1 U498 ( .A(n426), .B(KEYINPUT37), .ZN(n529) );
  XOR2_X1 U499 ( .A(n428), .B(n427), .Z(n430) );
  XNOR2_X1 U500 ( .A(G50GAT), .B(G36GAT), .ZN(n429) );
  XNOR2_X1 U501 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U502 ( .A(KEYINPUT30), .B(KEYINPUT70), .Z(n432) );
  NAND2_X1 U503 ( .A1(G229GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U504 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U505 ( .A(n434), .B(n433), .Z(n439) );
  XOR2_X1 U506 ( .A(KEYINPUT68), .B(G141GAT), .Z(n436) );
  XNOR2_X1 U507 ( .A(G113GAT), .B(G197GAT), .ZN(n435) );
  XNOR2_X1 U508 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U509 ( .A(n437), .B(KEYINPUT29), .ZN(n438) );
  XNOR2_X1 U510 ( .A(n439), .B(n438), .ZN(n441) );
  XNOR2_X1 U511 ( .A(n441), .B(n440), .ZN(n590) );
  INV_X1 U512 ( .A(n590), .ZN(n518) );
  XOR2_X1 U513 ( .A(KEYINPUT74), .B(KEYINPUT31), .Z(n443) );
  XNOR2_X1 U514 ( .A(G204GAT), .B(KEYINPUT32), .ZN(n442) );
  XNOR2_X1 U515 ( .A(n443), .B(n442), .ZN(n459) );
  XOR2_X1 U516 ( .A(KEYINPUT72), .B(KEYINPUT33), .Z(n445) );
  NAND2_X1 U517 ( .A1(G230GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U518 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U519 ( .A(n446), .B(KEYINPUT75), .Z(n450) );
  XNOR2_X1 U520 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U521 ( .A(n450), .B(n449), .ZN(n457) );
  XNOR2_X1 U522 ( .A(n452), .B(n451), .ZN(n455) );
  XNOR2_X1 U523 ( .A(n459), .B(n458), .ZN(n595) );
  OR2_X1 U524 ( .A1(n518), .A2(n595), .ZN(n502) );
  NOR2_X1 U525 ( .A1(n529), .A2(n502), .ZN(n462) );
  INV_X1 U526 ( .A(KEYINPUT102), .ZN(n460) );
  NOR2_X1 U527 ( .A1(n543), .A2(n515), .ZN(n466) );
  XNOR2_X1 U528 ( .A(KEYINPUT103), .B(KEYINPUT39), .ZN(n464) );
  INV_X1 U529 ( .A(G29GAT), .ZN(n463) );
  INV_X1 U530 ( .A(n599), .ZN(n497) );
  XNOR2_X1 U531 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n467) );
  XOR2_X1 U532 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n468) );
  XOR2_X1 U533 ( .A(KEYINPUT46), .B(n468), .Z(n469) );
  XNOR2_X1 U534 ( .A(n470), .B(n469), .ZN(n471) );
  AND2_X1 U535 ( .A1(n497), .A2(n471), .ZN(n472) );
  XNOR2_X1 U536 ( .A(n472), .B(KEYINPUT111), .ZN(n473) );
  NOR2_X1 U537 ( .A1(n473), .A2(n585), .ZN(n474) );
  XOR2_X1 U538 ( .A(n474), .B(KEYINPUT47), .Z(n483) );
  NOR2_X1 U539 ( .A1(n497), .A2(n490), .ZN(n477) );
  NOR2_X1 U540 ( .A1(n595), .A2(n478), .ZN(n479) );
  XNOR2_X1 U541 ( .A(n479), .B(KEYINPUT113), .ZN(n480) );
  NOR2_X1 U542 ( .A1(n590), .A2(n480), .ZN(n481) );
  XNOR2_X1 U543 ( .A(KEYINPUT114), .B(n481), .ZN(n482) );
  NOR2_X1 U544 ( .A1(n483), .A2(n482), .ZN(n484) );
  XNOR2_X1 U545 ( .A(n484), .B(KEYINPUT48), .ZN(n542) );
  NOR2_X1 U546 ( .A1(n513), .A2(n542), .ZN(n485) );
  XNOR2_X1 U547 ( .A(n485), .B(KEYINPUT54), .ZN(n486) );
  NAND2_X1 U548 ( .A1(n486), .A2(n543), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n487), .B(KEYINPUT65), .ZN(n572) );
  INV_X1 U550 ( .A(n572), .ZN(n488) );
  INV_X1 U551 ( .A(n600), .ZN(n489) );
  NOR2_X1 U552 ( .A1(n490), .A2(n489), .ZN(n493) );
  NOR2_X1 U553 ( .A1(n574), .A2(n515), .ZN(n494) );
  XNOR2_X1 U554 ( .A(n494), .B(KEYINPUT40), .ZN(n496) );
  INV_X1 U555 ( .A(G43GAT), .ZN(n495) );
  XNOR2_X1 U556 ( .A(n496), .B(n495), .ZN(G1330GAT) );
  NOR2_X1 U557 ( .A1(n497), .A2(n585), .ZN(n498) );
  XNOR2_X1 U558 ( .A(n498), .B(KEYINPUT16), .ZN(n501) );
  INV_X1 U559 ( .A(n499), .ZN(n500) );
  NAND2_X1 U560 ( .A1(n501), .A2(n500), .ZN(n519) );
  NOR2_X1 U561 ( .A1(n502), .A2(n519), .ZN(n509) );
  NAND2_X1 U562 ( .A1(n531), .A2(n509), .ZN(n503) );
  XNOR2_X1 U563 ( .A(n503), .B(KEYINPUT34), .ZN(n504) );
  XNOR2_X1 U564 ( .A(G1GAT), .B(n504), .ZN(G1324GAT) );
  NAND2_X1 U565 ( .A1(n533), .A2(n509), .ZN(n505) );
  XNOR2_X1 U566 ( .A(n505), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT35), .B(KEYINPUT98), .Z(n507) );
  NAND2_X1 U568 ( .A1(n509), .A2(n586), .ZN(n506) );
  XNOR2_X1 U569 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U570 ( .A(G15GAT), .B(n508), .ZN(G1326GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n511) );
  NAND2_X1 U572 ( .A1(n509), .A2(n548), .ZN(n510) );
  XNOR2_X1 U573 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U574 ( .A(G22GAT), .B(n512), .ZN(G1327GAT) );
  NOR2_X1 U575 ( .A1(n513), .A2(n515), .ZN(n514) );
  XOR2_X1 U576 ( .A(G36GAT), .B(n514), .Z(G1329GAT) );
  INV_X1 U577 ( .A(n548), .ZN(n516) );
  NOR2_X1 U578 ( .A1(n516), .A2(n515), .ZN(n517) );
  XOR2_X1 U579 ( .A(G50GAT), .B(n517), .Z(G1331GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT104), .B(KEYINPUT42), .Z(n521) );
  NAND2_X1 U581 ( .A1(n577), .A2(n518), .ZN(n528) );
  NOR2_X1 U582 ( .A1(n528), .A2(n519), .ZN(n525) );
  NAND2_X1 U583 ( .A1(n525), .A2(n531), .ZN(n520) );
  XNOR2_X1 U584 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U585 ( .A(G57GAT), .B(n522), .Z(G1332GAT) );
  NAND2_X1 U586 ( .A1(n533), .A2(n525), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n523), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U588 ( .A1(n525), .A2(n586), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n524), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U590 ( .A(G78GAT), .B(KEYINPUT43), .Z(n527) );
  NAND2_X1 U591 ( .A1(n525), .A2(n548), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n527), .B(n526), .ZN(G1335GAT) );
  NOR2_X1 U593 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U594 ( .A(KEYINPUT105), .B(n530), .Z(n538) );
  NAND2_X1 U595 ( .A1(n531), .A2(n538), .ZN(n532) );
  XNOR2_X1 U596 ( .A(n532), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U597 ( .A1(n533), .A2(n538), .ZN(n534) );
  XNOR2_X1 U598 ( .A(n534), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n536) );
  NAND2_X1 U600 ( .A1(n538), .A2(n586), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U602 ( .A(G99GAT), .B(n537), .ZN(G1338GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT108), .B(KEYINPUT44), .Z(n540) );
  NAND2_X1 U604 ( .A1(n538), .A2(n548), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U606 ( .A(G106GAT), .B(n541), .Z(G1339GAT) );
  NOR2_X1 U607 ( .A1(n543), .A2(n542), .ZN(n544) );
  NAND2_X1 U608 ( .A1(n545), .A2(n544), .ZN(n560) );
  NOR2_X1 U609 ( .A1(n574), .A2(n560), .ZN(n546) );
  XNOR2_X1 U610 ( .A(n546), .B(KEYINPUT115), .ZN(n547) );
  NOR2_X1 U611 ( .A1(n548), .A2(n547), .ZN(n556) );
  NAND2_X1 U612 ( .A1(n556), .A2(n590), .ZN(n549) );
  XNOR2_X1 U613 ( .A(n549), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U614 ( .A(G120GAT), .B(KEYINPUT49), .Z(n551) );
  NAND2_X1 U615 ( .A1(n556), .A2(n577), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n551), .B(n550), .ZN(G1341GAT) );
  XNOR2_X1 U617 ( .A(G127GAT), .B(KEYINPUT117), .ZN(n555) );
  XOR2_X1 U618 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n553) );
  NAND2_X1 U619 ( .A1(n556), .A2(n599), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(G1342GAT) );
  XOR2_X1 U622 ( .A(G134GAT), .B(KEYINPUT51), .Z(n558) );
  NAND2_X1 U623 ( .A1(n556), .A2(n585), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1343GAT) );
  XOR2_X1 U625 ( .A(G141GAT), .B(KEYINPUT119), .Z(n563) );
  NOR2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(KEYINPUT118), .ZN(n568) );
  NAND2_X1 U628 ( .A1(n590), .A2(n568), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1344GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n565) );
  NAND2_X1 U631 ( .A1(n577), .A2(n568), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U633 ( .A(G148GAT), .B(n566), .ZN(G1345GAT) );
  NAND2_X1 U634 ( .A1(n568), .A2(n599), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n567), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U636 ( .A1(n568), .A2(n585), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n569), .B(KEYINPUT120), .ZN(n570) );
  XNOR2_X1 U638 ( .A(G162GAT), .B(n570), .ZN(G1347GAT) );
  XOR2_X1 U639 ( .A(G169GAT), .B(KEYINPUT121), .Z(n576) );
  AND2_X1 U640 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U641 ( .A(n573), .B(KEYINPUT55), .ZN(n587) );
  NOR2_X1 U642 ( .A1(n574), .A2(n587), .ZN(n582) );
  NAND2_X1 U643 ( .A1(n582), .A2(n590), .ZN(n575) );
  XNOR2_X1 U644 ( .A(n576), .B(n575), .ZN(G1348GAT) );
  XNOR2_X1 U645 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n581) );
  XOR2_X1 U646 ( .A(KEYINPUT122), .B(KEYINPUT56), .Z(n579) );
  XNOR2_X1 U647 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U648 ( .A(n581), .B(n580), .ZN(G1349GAT) );
  XOR2_X1 U649 ( .A(G183GAT), .B(KEYINPUT123), .Z(n584) );
  NAND2_X1 U650 ( .A1(n582), .A2(n599), .ZN(n583) );
  XNOR2_X1 U651 ( .A(n584), .B(n583), .ZN(G1350GAT) );
  OR2_X1 U652 ( .A1(n587), .A2(n296), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n588), .B(KEYINPUT58), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n589), .B(G190GAT), .ZN(G1351GAT) );
  XNOR2_X1 U655 ( .A(KEYINPUT60), .B(KEYINPUT124), .ZN(n594) );
  XOR2_X1 U656 ( .A(G197GAT), .B(KEYINPUT59), .Z(n592) );
  NAND2_X1 U657 ( .A1(n600), .A2(n590), .ZN(n591) );
  XNOR2_X1 U658 ( .A(n592), .B(n591), .ZN(n593) );
  XNOR2_X1 U659 ( .A(n594), .B(n593), .ZN(G1352GAT) );
  XOR2_X1 U660 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n597) );
  NAND2_X1 U661 ( .A1(n600), .A2(n595), .ZN(n596) );
  XNOR2_X1 U662 ( .A(n597), .B(n596), .ZN(n598) );
  XOR2_X1 U663 ( .A(G204GAT), .B(n598), .Z(G1353GAT) );
  XOR2_X1 U664 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n602) );
  NAND2_X1 U665 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U666 ( .A(n602), .B(n601), .ZN(n603) );
  XNOR2_X1 U667 ( .A(G211GAT), .B(n603), .ZN(G1354GAT) );
endmodule

