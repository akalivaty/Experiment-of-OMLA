//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 1 0 1 0 0 0 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 0 1 1 0 0 0 0 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n774, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n872, new_n873, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n950, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT13), .Z(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT14), .B(G29gat), .ZN(new_n204));
  INV_X1    g003(.A(G36gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(G43gat), .B(G50gat), .Z(new_n207));
  INV_X1    g006(.A(G29gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n208), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n206), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  AOI22_X1  g010(.A1(new_n206), .A2(new_n209), .B1(new_n207), .B2(KEYINPUT86), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT15), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G15gat), .B(G22gat), .ZN(new_n214));
  INV_X1    g013(.A(G1gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT16), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(G1gat), .B2(new_n214), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G8gat), .ZN(new_n219));
  INV_X1    g018(.A(G8gat), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n217), .B(new_n220), .C1(G1gat), .C2(new_n214), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n209), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n207), .A2(KEYINPUT86), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT15), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AND3_X1   g026(.A1(new_n213), .A2(new_n222), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n222), .B1(new_n213), .B2(new_n227), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n203), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT87), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT87), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n232), .B(new_n203), .C1(new_n228), .C2(new_n229), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n226), .B1(new_n225), .B2(new_n210), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n212), .A2(KEYINPUT15), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT17), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT17), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n213), .A2(new_n238), .A3(new_n227), .ZN(new_n239));
  INV_X1    g038(.A(new_n222), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n237), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n228), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n241), .A2(new_n242), .A3(KEYINPUT18), .A4(new_n202), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n241), .A2(new_n242), .A3(new_n202), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT18), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G113gat), .B(G141gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT85), .B(G197gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT11), .B(G169gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(KEYINPUT12), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n234), .A2(new_n243), .A3(new_n246), .A4(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT88), .ZN(new_n254));
  AOI22_X1  g053(.A1(new_n231), .A2(new_n233), .B1(new_n244), .B2(new_n245), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n252), .B1(new_n255), .B2(new_n243), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  AOI211_X1 g056(.A(KEYINPUT88), .B(new_n252), .C1(new_n255), .C2(new_n243), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(G127gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n261), .A2(G134gat), .ZN(new_n262));
  INV_X1    g061(.A(G134gat), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n263), .A2(G127gat), .ZN(new_n264));
  OAI21_X1  g063(.A(KEYINPUT70), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(G127gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n261), .A2(G134gat), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(G113gat), .ZN(new_n270));
  INV_X1    g069(.A(G120gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT1), .ZN(new_n273));
  NAND2_X1  g072(.A1(G113gat), .A2(G120gat), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  AND3_X1   g074(.A1(new_n265), .A2(new_n269), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n266), .A2(new_n267), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT1), .B1(new_n270), .B2(new_n271), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n277), .A2(KEYINPUT70), .A3(new_n274), .A4(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G155gat), .A2(G162gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT2), .ZN(new_n282));
  INV_X1    g081(.A(G141gat), .ZN(new_n283));
  INV_X1    g082(.A(G148gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G141gat), .A2(G148gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n282), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT75), .ZN(new_n288));
  XNOR2_X1  g087(.A(G155gat), .B(G162gat), .ZN(new_n289));
  AND3_X1   g088(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n289), .B1(new_n287), .B2(new_n288), .ZN(new_n291));
  OAI22_X1  g090(.A1(new_n276), .A2(new_n280), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G225gat), .A2(G233gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n265), .A2(new_n269), .A3(new_n275), .ZN(new_n296));
  AND3_X1   g095(.A1(new_n296), .A2(KEYINPUT76), .A3(new_n279), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT76), .B1(new_n296), .B2(new_n279), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n287), .A2(new_n288), .ZN(new_n300));
  INV_X1    g099(.A(new_n289), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n292), .B(new_n295), .C1(new_n299), .C2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT3), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n306), .B1(new_n290), .B2(new_n291), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT77), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n304), .A2(KEYINPUT77), .A3(new_n306), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n296), .A2(new_n279), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT76), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n296), .A2(new_n279), .A3(KEYINPUT76), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n290), .A2(new_n291), .ZN(new_n316));
  AOI22_X1  g115(.A1(new_n314), .A2(new_n315), .B1(new_n316), .B2(KEYINPUT3), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT4), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n304), .A2(new_n318), .A3(new_n312), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n292), .A2(KEYINPUT4), .ZN(new_n320));
  AOI22_X1  g119(.A1(new_n311), .A2(new_n317), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n293), .B1(new_n321), .B2(KEYINPUT5), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n294), .B1(new_n311), .B2(new_n317), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT79), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT78), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n302), .A2(new_n303), .B1(new_n296), .B2(new_n279), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n326), .B1(new_n327), .B2(new_n318), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n292), .A2(KEYINPUT78), .A3(KEYINPUT4), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n327), .A2(KEYINPUT79), .A3(new_n318), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n325), .A2(new_n328), .A3(new_n329), .A4(new_n330), .ZN(new_n331));
  AND2_X1   g130(.A1(new_n323), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n305), .B1(new_n322), .B2(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(G1gat), .B(G29gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n334), .B(KEYINPUT0), .ZN(new_n335));
  XNOR2_X1  g134(.A(G57gat), .B(G85gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n335), .B(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT6), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n302), .A2(KEYINPUT3), .A3(new_n303), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n339), .B1(new_n297), .B2(new_n298), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n340), .B1(new_n309), .B2(new_n310), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n320), .A2(new_n319), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n294), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n323), .A2(new_n331), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n344), .A2(new_n345), .A3(new_n293), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT80), .ZN(new_n347));
  INV_X1    g146(.A(new_n337), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n346), .A2(new_n347), .A3(new_n348), .A4(new_n305), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n348), .B(new_n305), .C1(new_n322), .C2(new_n332), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT80), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n338), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n348), .B1(new_n346), .B2(new_n305), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT6), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G8gat), .B(G36gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(G64gat), .B(G92gat), .ZN(new_n357));
  XOR2_X1   g156(.A(new_n356), .B(new_n357), .Z(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(G226gat), .A2(G233gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(G169gat), .ZN(new_n362));
  INV_X1    g161(.A(G176gat), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT26), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n362), .B(new_n363), .C1(new_n364), .C2(KEYINPUT69), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(KEYINPUT69), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NOR2_X1   g166(.A1(G169gat), .A2(G176gat), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n368), .A2(KEYINPUT69), .A3(new_n364), .ZN(new_n369));
  NAND2_X1  g168(.A1(G169gat), .A2(G176gat), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n367), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(G183gat), .A2(G190gat), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT27), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(G183gat), .ZN(new_n375));
  INV_X1    g174(.A(G183gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT27), .ZN(new_n377));
  INV_X1    g176(.A(G190gat), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n375), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n373), .B1(new_n379), .B2(KEYINPUT28), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT67), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(new_n376), .ZN(new_n382));
  NAND2_X1  g181(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n382), .A2(KEYINPUT27), .A3(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n374), .A2(KEYINPUT68), .A3(G183gat), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT68), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n375), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g186(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n384), .A2(new_n385), .A3(new_n387), .A4(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n371), .A2(new_n380), .A3(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n376), .A2(new_n378), .A3(KEYINPUT64), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT64), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n392), .B1(G183gat), .B2(G190gat), .ZN(new_n393));
  AND2_X1   g192(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n372), .A2(KEYINPUT24), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT24), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n396), .A2(G183gat), .A3(G190gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(KEYINPUT66), .B1(new_n368), .B2(KEYINPUT23), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT66), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT23), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n400), .B(new_n401), .C1(G169gat), .C2(G176gat), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n394), .A2(new_n398), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n362), .A2(new_n363), .A3(KEYINPUT23), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT65), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n368), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n406), .A2(new_n370), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT25), .B1(new_n403), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n382), .A2(new_n383), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n398), .B1(new_n411), .B2(G190gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n399), .A2(new_n402), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n404), .A2(KEYINPUT25), .A3(new_n370), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n390), .B1(new_n410), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT29), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n361), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AND3_X1   g218(.A1(new_n371), .A2(new_n380), .A3(new_n389), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT25), .ZN(new_n421));
  INV_X1    g220(.A(new_n398), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n391), .A2(new_n393), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n413), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n421), .B1(new_n424), .B2(new_n408), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n420), .B1(new_n425), .B2(new_n415), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n426), .A2(new_n360), .ZN(new_n427));
  XNOR2_X1  g226(.A(G197gat), .B(G204gat), .ZN(new_n428));
  INV_X1    g227(.A(G211gat), .ZN(new_n429));
  INV_X1    g228(.A(G218gat), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n428), .B1(KEYINPUT22), .B2(new_n431), .ZN(new_n432));
  XOR2_X1   g231(.A(G211gat), .B(G218gat), .Z(new_n433));
  XOR2_X1   g232(.A(new_n432), .B(new_n433), .Z(new_n434));
  NOR3_X1   g233(.A1(new_n419), .A2(new_n427), .A3(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n434), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n360), .B1(new_n426), .B2(KEYINPUT29), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n417), .A2(new_n361), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n359), .B1(new_n435), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n434), .B1(new_n419), .B2(new_n427), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n437), .A2(new_n436), .A3(new_n438), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n441), .A2(new_n442), .A3(new_n358), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n440), .A2(KEYINPUT30), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT30), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n441), .A2(new_n442), .A3(new_n445), .A4(new_n358), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n355), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT81), .ZN(new_n449));
  NAND2_X1  g248(.A1(G227gat), .A2(G233gat), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT72), .B1(new_n426), .B2(new_n312), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT72), .ZN(new_n452));
  INV_X1    g251(.A(new_n312), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n417), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n312), .B(new_n390), .C1(new_n410), .C2(new_n416), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT71), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n425), .A2(new_n415), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n459), .A2(KEYINPUT71), .A3(new_n312), .A4(new_n390), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n450), .B1(new_n455), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT32), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT73), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  XOR2_X1   g263(.A(G71gat), .B(G99gat), .Z(new_n465));
  XNOR2_X1  g264(.A(G15gat), .B(G43gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n465), .B(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT73), .ZN(new_n468));
  AOI22_X1  g267(.A1(new_n451), .A2(new_n454), .B1(new_n458), .B2(new_n460), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n468), .B(KEYINPUT32), .C1(new_n469), .C2(new_n450), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT33), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n471), .B1(new_n469), .B2(new_n450), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n464), .A2(new_n467), .A3(new_n470), .A4(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n469), .A2(new_n450), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT74), .ZN(new_n475));
  OR2_X1    g274(.A1(new_n475), .A2(KEYINPUT34), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(KEYINPUT34), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n474), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n478), .B1(new_n474), .B2(new_n477), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n467), .A2(KEYINPUT33), .ZN(new_n480));
  OAI211_X1 g279(.A(KEYINPUT32), .B(new_n480), .C1(new_n469), .C2(new_n450), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n473), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n479), .B1(new_n473), .B2(new_n481), .ZN(new_n484));
  NAND2_X1  g283(.A1(G228gat), .A2(G233gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n485), .B(G22gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(KEYINPUT31), .B(G50gat), .ZN(new_n487));
  XOR2_X1   g286(.A(new_n486), .B(new_n487), .Z(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n311), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n434), .B1(new_n490), .B2(KEYINPUT29), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n306), .B1(new_n434), .B2(KEYINPUT29), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(new_n316), .ZN(new_n493));
  XNOR2_X1  g292(.A(G78gat), .B(G106gat), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n491), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n495), .B1(new_n491), .B2(new_n493), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n489), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n498), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n500), .A2(new_n496), .A3(new_n488), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NOR3_X1   g301(.A1(new_n483), .A2(new_n484), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT81), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n355), .A2(new_n504), .A3(new_n447), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n449), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(KEYINPUT35), .ZN(new_n507));
  AND3_X1   g306(.A1(new_n444), .A2(KEYINPUT83), .A3(new_n446), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT83), .B1(new_n444), .B2(new_n446), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n502), .A2(KEYINPUT35), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n510), .A2(new_n355), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n473), .A2(new_n481), .ZN(new_n513));
  INV_X1    g312(.A(new_n479), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n482), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n507), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n443), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT37), .B1(new_n435), .B2(new_n439), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT37), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n441), .A2(new_n442), .A3(new_n522), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n521), .A2(new_n359), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(KEYINPUT84), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT38), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n520), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n521), .A2(new_n359), .A3(new_n523), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n528), .A2(KEYINPUT38), .A3(new_n525), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n527), .A2(new_n352), .A3(new_n354), .A4(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n509), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n444), .A2(KEYINPUT83), .A3(new_n446), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n311), .A2(new_n317), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n293), .B1(new_n534), .B2(new_n342), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT39), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n337), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n292), .B(new_n293), .C1(new_n299), .C2(new_n304), .ZN(new_n538));
  OAI211_X1 g337(.A(KEYINPUT39), .B(new_n538), .C1(new_n321), .C2(new_n293), .ZN(new_n539));
  AND3_X1   g338(.A1(new_n537), .A2(KEYINPUT40), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT40), .B1(new_n537), .B2(new_n539), .ZN(new_n541));
  NOR3_X1   g340(.A1(new_n540), .A2(new_n353), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n502), .B1(new_n533), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT36), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n544), .B1(new_n483), .B2(new_n484), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n515), .A2(KEYINPUT36), .A3(new_n482), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n530), .A2(new_n543), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n502), .B(KEYINPUT82), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n355), .A2(new_n504), .A3(new_n447), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n504), .B1(new_n355), .B2(new_n447), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n260), .B1(new_n519), .B2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G120gat), .B(G148gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(KEYINPUT101), .ZN(new_n555));
  XNOR2_X1  g354(.A(G176gat), .B(G204gat), .ZN(new_n556));
  XOR2_X1   g355(.A(new_n555), .B(new_n556), .Z(new_n557));
  XOR2_X1   g356(.A(G57gat), .B(G64gat), .Z(new_n558));
  INV_X1    g357(.A(KEYINPUT9), .ZN(new_n559));
  INV_X1    g358(.A(G71gat), .ZN(new_n560));
  INV_X1    g359(.A(G78gat), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G71gat), .B(G78gat), .ZN(new_n564));
  AND2_X1   g363(.A1(new_n564), .A2(KEYINPUT89), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n564), .A2(KEYINPUT89), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n563), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT90), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT90), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n569), .B(new_n563), .C1(new_n565), .C2(new_n566), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n558), .A2(new_n562), .A3(new_n564), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT91), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT96), .B(G92gat), .ZN(new_n574));
  INV_X1    g373(.A(G85gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(G99gat), .A2(G106gat), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT8), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(KEYINPUT94), .A2(G85gat), .A3(G92gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(KEYINPUT93), .ZN(new_n581));
  NAND2_X1  g380(.A1(G85gat), .A2(G92gat), .ZN(new_n582));
  OAI211_X1 g381(.A(new_n581), .B(KEYINPUT7), .C1(KEYINPUT93), .C2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT7), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n580), .A2(KEYINPUT93), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(KEYINPUT95), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT95), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n583), .A2(new_n588), .A3(new_n585), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n579), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G99gat), .B(G106gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT99), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n571), .B(new_n573), .C1(new_n590), .C2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n579), .ZN(new_n594));
  INV_X1    g393(.A(new_n589), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n588), .B1(new_n583), .B2(new_n585), .ZN(new_n596));
  OAI211_X1 g395(.A(new_n591), .B(new_n594), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT97), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n590), .A2(KEYINPUT97), .A3(new_n591), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n593), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n597), .A2(new_n598), .ZN(new_n603));
  AOI21_X1  g402(.A(KEYINPUT97), .B1(new_n590), .B2(new_n591), .ZN(new_n604));
  OAI22_X1  g403(.A1(new_n603), .A2(new_n604), .B1(new_n591), .B2(new_n590), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n571), .A2(new_n573), .ZN(new_n606));
  AOI21_X1  g405(.A(KEYINPUT98), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n590), .A2(new_n591), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n608), .B1(new_n599), .B2(new_n600), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT98), .ZN(new_n610));
  INV_X1    g409(.A(new_n606), .ZN(new_n611));
  NOR3_X1   g410(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n602), .B1(new_n607), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G230gat), .A2(G233gat), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n613), .A2(KEYINPUT100), .A3(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT100), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n605), .A2(KEYINPUT98), .A3(new_n606), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n610), .B1(new_n609), .B2(new_n611), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n601), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n617), .B1(new_n620), .B2(new_n614), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT10), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n623), .B(new_n602), .C1(new_n607), .C2(new_n612), .ZN(new_n624));
  NOR3_X1   g423(.A1(new_n605), .A2(new_n623), .A3(new_n606), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n615), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n557), .B1(new_n622), .B2(new_n627), .ZN(new_n628));
  AOI211_X1 g427(.A(KEYINPUT10), .B(new_n601), .C1(new_n618), .C2(new_n619), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n614), .B1(new_n629), .B2(new_n625), .ZN(new_n630));
  INV_X1    g429(.A(new_n557), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n630), .A2(new_n631), .A3(new_n621), .A4(new_n616), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n611), .A2(KEYINPUT21), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  OR3_X1    g435(.A1(new_n636), .A2(KEYINPUT92), .A3(new_n222), .ZN(new_n637));
  OAI21_X1  g436(.A(KEYINPUT92), .B1(new_n636), .B2(new_n222), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n640));
  INV_X1    g439(.A(G155gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n642), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n637), .A2(new_n638), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT21), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n606), .A2(new_n647), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n648), .A2(G231gat), .A3(G233gat), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n648), .B1(G231gat), .B2(G233gat), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(new_n261), .ZN(new_n652));
  XNOR2_X1  g451(.A(G183gat), .B(G211gat), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(G127gat), .B1(new_n649), .B2(new_n650), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n652), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n654), .B1(new_n652), .B2(new_n655), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n646), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n658), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n660), .A2(new_n656), .A3(new_n645), .A4(new_n643), .ZN(new_n661));
  NOR3_X1   g460(.A1(new_n605), .A2(new_n235), .A3(new_n236), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n237), .A2(new_n239), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT41), .ZN(new_n664));
  NAND2_X1  g463(.A1(G232gat), .A2(G233gat), .ZN(new_n665));
  OAI22_X1  g464(.A1(new_n609), .A2(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g466(.A(G190gat), .B(G218gat), .Z(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(G134gat), .B(G162gat), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n665), .A2(new_n664), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n672), .B(new_n673), .Z(new_n674));
  NAND2_X1  g473(.A1(new_n667), .A2(new_n669), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n671), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n674), .ZN(new_n677));
  INV_X1    g476(.A(new_n675), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n677), .B1(new_n678), .B2(new_n670), .ZN(new_n679));
  AOI22_X1  g478(.A1(new_n659), .A2(new_n661), .B1(new_n676), .B2(new_n679), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n634), .A2(new_n680), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n553), .A2(new_n681), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n355), .A2(KEYINPUT102), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n355), .A2(KEYINPUT102), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g487(.A1(new_n682), .A2(new_n533), .ZN(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT16), .B(G8gat), .ZN(new_n690));
  OAI21_X1  g489(.A(KEYINPUT103), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  OR2_X1    g490(.A1(new_n691), .A2(KEYINPUT42), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n689), .A2(G8gat), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(KEYINPUT42), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(G1325gat));
  INV_X1    g494(.A(new_n682), .ZN(new_n696));
  OR3_X1    g495(.A1(new_n696), .A2(G15gat), .A3(new_n516), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n483), .A2(new_n484), .A3(new_n544), .ZN(new_n698));
  AOI21_X1  g497(.A(KEYINPUT36), .B1(new_n515), .B2(new_n482), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(G15gat), .B1(new_n696), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n697), .A2(new_n702), .ZN(G1326gat));
  NAND2_X1  g502(.A1(new_n682), .A2(new_n548), .ZN(new_n704));
  XNOR2_X1  g503(.A(KEYINPUT43), .B(G22gat), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1327gat));
  NAND2_X1  g505(.A1(new_n659), .A2(new_n661), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n679), .A2(new_n676), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n553), .A2(new_n708), .A3(new_n710), .A4(new_n634), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n711), .A2(G29gat), .A3(new_n685), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n712), .B(KEYINPUT45), .Z(new_n713));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n714));
  INV_X1    g513(.A(new_n548), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n715), .B1(new_n449), .B2(new_n505), .ZN(new_n716));
  INV_X1    g515(.A(new_n502), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n542), .B1(new_n508), .B2(new_n509), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n530), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n698), .B2(new_n699), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n714), .B1(new_n716), .B2(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n547), .A2(new_n551), .A3(KEYINPUT105), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n709), .B1(new_n723), .B2(new_n519), .ZN(new_n724));
  XNOR2_X1  g523(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n519), .A2(new_n552), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(new_n710), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(KEYINPUT44), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n634), .A2(KEYINPUT104), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n634), .A2(KEYINPUT104), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n734), .A2(new_n260), .A3(new_n707), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n731), .A2(new_n685), .A3(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n713), .B1(new_n208), .B2(new_n737), .ZN(G1328gat));
  NOR3_X1   g537(.A1(new_n711), .A2(G36gat), .A3(new_n510), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT46), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n731), .A2(new_n510), .A3(new_n736), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n741), .B2(new_n205), .ZN(G1329gat));
  OR3_X1    g541(.A1(new_n711), .A2(G43gat), .A3(new_n516), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n731), .A2(new_n701), .A3(new_n736), .ZN(new_n744));
  INV_X1    g543(.A(G43gat), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT47), .B1(new_n743), .B2(KEYINPUT107), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(G1330gat));
  NAND3_X1  g547(.A1(new_n730), .A2(new_n548), .A3(new_n735), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G50gat), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n711), .A2(G50gat), .A3(new_n715), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n751), .A2(KEYINPUT48), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT48), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n730), .A2(new_n502), .A3(new_n735), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n751), .B1(new_n755), .B2(G50gat), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n753), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT108), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT108), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n753), .B(new_n759), .C1(new_n754), .C2(new_n756), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(G1331gat));
  NAND2_X1  g560(.A1(new_n723), .A2(new_n519), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n680), .A2(new_n260), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n762), .A2(new_n734), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n686), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n533), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n768));
  XOR2_X1   g567(.A(KEYINPUT49), .B(G64gat), .Z(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n767), .B2(new_n769), .ZN(G1333gat));
  AOI21_X1  g569(.A(new_n560), .B1(new_n764), .B2(new_n700), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n516), .A2(G71gat), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n771), .B1(new_n764), .B2(new_n772), .ZN(new_n773));
  XNOR2_X1  g572(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n773), .B(new_n774), .ZN(G1334gat));
  NAND2_X1  g574(.A1(new_n764), .A2(new_n548), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g576(.A1(new_n708), .A2(new_n260), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n762), .A2(KEYINPUT51), .A3(new_n710), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT110), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n762), .A2(new_n710), .A3(new_n779), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT51), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT110), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n724), .A2(new_n785), .A3(KEYINPUT51), .A4(new_n779), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n781), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n787), .A2(new_n575), .A3(new_n633), .A4(new_n686), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n778), .A2(new_n634), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n730), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(G85gat), .B1(new_n790), .B2(new_n685), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n788), .A2(new_n791), .ZN(G1336gat));
  AND2_X1   g591(.A1(new_n730), .A2(new_n789), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n574), .B1(new_n793), .B2(new_n533), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n794), .A2(KEYINPUT52), .ZN(new_n795));
  INV_X1    g594(.A(new_n787), .ZN(new_n796));
  INV_X1    g595(.A(new_n734), .ZN(new_n797));
  OR3_X1    g596(.A1(new_n797), .A2(G92gat), .A3(new_n510), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n795), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n798), .B1(new_n784), .B2(new_n780), .ZN(new_n800));
  OAI21_X1  g599(.A(KEYINPUT52), .B1(new_n794), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(G1337gat));
  NOR2_X1   g601(.A1(new_n516), .A2(G99gat), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n787), .A2(new_n633), .A3(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(G99gat), .B1(new_n790), .B2(new_n701), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(KEYINPUT111), .ZN(G1338gat));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n797), .A2(G106gat), .A3(new_n717), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT51), .B1(new_n724), .B2(new_n779), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n517), .B1(new_n506), .B2(KEYINPUT35), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n811), .B1(new_n721), .B2(new_n722), .ZN(new_n812));
  NOR4_X1   g611(.A1(new_n812), .A2(new_n783), .A3(new_n709), .A4(new_n778), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n809), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n725), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n812), .A2(new_n709), .A3(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT44), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n817), .B1(new_n727), .B2(new_n710), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n548), .B(new_n789), .C1(new_n816), .C2(new_n818), .ZN(new_n819));
  AOI22_X1  g618(.A1(new_n814), .A2(KEYINPUT112), .B1(new_n819), .B2(G106gat), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT112), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n821), .B(new_n809), .C1(new_n810), .C2(new_n813), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n808), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n787), .A2(new_n809), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n502), .B(new_n789), .C1(new_n816), .C2(new_n818), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT53), .B1(new_n825), .B2(G106gat), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT113), .B1(new_n823), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n814), .A2(KEYINPUT112), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n819), .A2(G106gat), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n829), .A2(new_n822), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT53), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT113), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n824), .A2(new_n826), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n828), .A2(new_n835), .ZN(G1339gat));
  NAND2_X1  g635(.A1(new_n763), .A2(new_n634), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n626), .A2(new_n615), .ZN(new_n838));
  OAI21_X1  g637(.A(KEYINPUT54), .B1(new_n629), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(KEYINPUT55), .B1(new_n839), .B2(new_n627), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n841), .B(new_n614), .C1(new_n629), .C2(new_n625), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n557), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n632), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n631), .B1(new_n627), .B2(new_n841), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n625), .A2(new_n614), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n841), .B1(new_n624), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n630), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(KEYINPUT55), .B1(new_n845), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n202), .B1(new_n241), .B2(new_n242), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n228), .A2(new_n229), .A3(new_n203), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n251), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n253), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n679), .A2(new_n676), .A3(new_n854), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n844), .A2(new_n849), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n633), .A2(new_n854), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n259), .B(new_n632), .C1(new_n840), .C2(new_n843), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n857), .B1(new_n849), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n856), .B1(new_n859), .B2(new_n709), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n837), .B1(new_n860), .B2(new_n707), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n861), .A2(new_n686), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n862), .A2(new_n510), .A3(new_n503), .ZN(new_n863));
  AOI21_X1  g662(.A(G113gat), .B1(new_n863), .B2(new_n259), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n861), .A2(new_n715), .ZN(new_n865));
  NOR4_X1   g664(.A1(new_n865), .A2(new_n516), .A3(new_n533), .A4(new_n685), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n260), .A2(new_n270), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n864), .B1(new_n866), .B2(new_n867), .ZN(G1340gat));
  AOI21_X1  g667(.A(G120gat), .B1(new_n863), .B2(new_n633), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n797), .A2(new_n271), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n869), .B1(new_n866), .B2(new_n870), .ZN(G1341gat));
  AND2_X1   g670(.A1(new_n863), .A2(new_n707), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n872), .A2(KEYINPUT114), .ZN(new_n873));
  AOI21_X1  g672(.A(G127gat), .B1(new_n872), .B2(KEYINPUT114), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n708), .A2(new_n261), .ZN(new_n875));
  AOI22_X1  g674(.A1(new_n873), .A2(new_n874), .B1(new_n866), .B2(new_n875), .ZN(G1342gat));
  AND2_X1   g675(.A1(new_n866), .A2(new_n710), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n877), .A2(new_n263), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n863), .A2(new_n263), .A3(new_n710), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n878), .B1(KEYINPUT56), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n880), .B1(KEYINPUT56), .B2(new_n879), .ZN(G1343gat));
  NOR3_X1   g680(.A1(new_n700), .A2(new_n717), .A3(new_n533), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n862), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n283), .B1(new_n883), .B2(new_n260), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n685), .A2(new_n700), .A3(new_n533), .ZN(new_n885));
  XNOR2_X1  g684(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n887), .B1(new_n845), .B2(new_n848), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n858), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n853), .B1(new_n628), .B2(new_n632), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n709), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(new_n856), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n707), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n837), .ZN(new_n894));
  OAI211_X1 g693(.A(KEYINPUT57), .B(new_n548), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(KEYINPUT57), .B1(new_n861), .B2(new_n502), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT115), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI211_X1 g697(.A(KEYINPUT115), .B(KEYINPUT57), .C1(new_n861), .C2(new_n502), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n885), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n259), .A2(G141gat), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n884), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  XOR2_X1   g701(.A(new_n902), .B(KEYINPUT58), .Z(G1344gat));
  INV_X1    g702(.A(KEYINPUT119), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n633), .B(new_n885), .C1(new_n898), .C2(new_n899), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n284), .A2(KEYINPUT59), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n861), .A2(new_n502), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(KEYINPUT57), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n885), .A2(new_n633), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n837), .A2(KEYINPUT117), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT117), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n763), .A2(new_n911), .A3(new_n634), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n891), .A2(new_n892), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n707), .B1(new_n914), .B2(KEYINPUT118), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT118), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n891), .A2(new_n916), .A3(new_n892), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n913), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT57), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n548), .A2(new_n919), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n908), .B(new_n909), .C1(new_n918), .C2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(G148gat), .ZN(new_n922));
  AOI22_X1  g721(.A1(new_n905), .A2(new_n906), .B1(new_n922), .B2(KEYINPUT59), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n883), .A2(G148gat), .A3(new_n634), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n904), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n905), .A2(new_n906), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n922), .A2(KEYINPUT59), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(new_n924), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n928), .A2(KEYINPUT119), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n925), .A2(new_n930), .ZN(G1345gat));
  OAI21_X1  g730(.A(G155gat), .B1(new_n900), .B2(new_n708), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n707), .A2(new_n641), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n883), .B2(new_n933), .ZN(G1346gat));
  NOR3_X1   g733(.A1(new_n883), .A2(G162gat), .A3(new_n709), .ZN(new_n935));
  XOR2_X1   g734(.A(new_n935), .B(KEYINPUT120), .Z(new_n936));
  OAI21_X1  g735(.A(G162gat), .B1(new_n900), .B2(new_n709), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1347gat));
  AND4_X1   g737(.A1(new_n533), .A2(new_n861), .A3(new_n503), .A4(new_n685), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n939), .A2(new_n362), .A3(new_n259), .ZN(new_n940));
  XOR2_X1   g739(.A(new_n940), .B(KEYINPUT121), .Z(new_n941));
  NAND2_X1  g740(.A1(new_n685), .A2(new_n533), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n865), .A2(new_n516), .A3(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  OAI21_X1  g743(.A(G169gat), .B1(new_n944), .B2(new_n260), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n941), .A2(new_n945), .ZN(G1348gat));
  OAI21_X1  g745(.A(G176gat), .B1(new_n944), .B2(new_n797), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n939), .A2(new_n363), .A3(new_n633), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(G1349gat));
  NAND2_X1  g748(.A1(new_n943), .A2(new_n707), .ZN(new_n950));
  AND3_X1   g749(.A1(new_n707), .A2(new_n375), .A3(new_n377), .ZN(new_n951));
  AOI22_X1  g750(.A1(new_n950), .A2(new_n411), .B1(new_n939), .B2(new_n951), .ZN(new_n952));
  XOR2_X1   g751(.A(KEYINPUT122), .B(KEYINPUT60), .Z(new_n953));
  XNOR2_X1  g752(.A(new_n952), .B(new_n953), .ZN(G1350gat));
  NAND3_X1  g753(.A1(new_n939), .A2(new_n378), .A3(new_n710), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n943), .A2(new_n710), .ZN(new_n956));
  XNOR2_X1  g755(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n956), .A2(G190gat), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n957), .B1(new_n956), .B2(G190gat), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n955), .B1(new_n958), .B2(new_n959), .ZN(G1351gat));
  NOR2_X1   g759(.A1(new_n942), .A2(new_n700), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n907), .A2(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(new_n963), .ZN(new_n964));
  OR3_X1    g763(.A1(new_n964), .A2(G197gat), .A3(new_n260), .ZN(new_n965));
  OAI211_X1 g764(.A(new_n908), .B(new_n961), .C1(new_n918), .C2(new_n920), .ZN(new_n966));
  OAI21_X1  g765(.A(KEYINPUT124), .B1(new_n966), .B2(new_n260), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(G197gat), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n966), .A2(KEYINPUT124), .A3(new_n260), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n965), .B1(new_n968), .B2(new_n969), .ZN(G1352gat));
  XNOR2_X1  g769(.A(KEYINPUT125), .B(G204gat), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n963), .A2(new_n633), .A3(new_n971), .ZN(new_n972));
  XOR2_X1   g771(.A(new_n972), .B(KEYINPUT62), .Z(new_n973));
  NOR2_X1   g772(.A1(new_n966), .A2(new_n797), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n973), .B1(new_n974), .B2(new_n971), .ZN(G1353gat));
  NAND3_X1  g774(.A1(new_n963), .A2(new_n429), .A3(new_n707), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n845), .A2(new_n848), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(new_n886), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n845), .A2(new_n848), .A3(KEYINPUT55), .ZN(new_n979));
  NAND4_X1  g778(.A1(new_n978), .A2(new_n259), .A3(new_n632), .A4(new_n979), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n710), .B1(new_n980), .B2(new_n857), .ZN(new_n981));
  OAI21_X1  g780(.A(KEYINPUT118), .B1(new_n981), .B2(new_n856), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n982), .A2(new_n708), .A3(new_n917), .ZN(new_n983));
  INV_X1    g782(.A(new_n913), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n920), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n919), .B1(new_n861), .B2(new_n502), .ZN(new_n986));
  NOR3_X1   g785(.A1(new_n985), .A2(new_n986), .A3(new_n962), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n987), .A2(new_n707), .ZN(new_n988));
  AND3_X1   g787(.A1(new_n988), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n989));
  AOI21_X1  g788(.A(KEYINPUT63), .B1(new_n988), .B2(G211gat), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n976), .B1(new_n989), .B2(new_n990), .ZN(G1354gat));
  OAI21_X1  g790(.A(new_n430), .B1(new_n964), .B2(new_n709), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n709), .A2(new_n430), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n993), .B1(new_n987), .B2(KEYINPUT126), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT126), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n966), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n992), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT127), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI211_X1 g798(.A(KEYINPUT127), .B(new_n992), .C1(new_n994), .C2(new_n996), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n999), .A2(new_n1000), .ZN(G1355gat));
endmodule


