

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591;

  XNOR2_X1 U326 ( .A(n408), .B(n407), .ZN(n429) );
  INV_X1 U327 ( .A(KEYINPUT113), .ZN(n406) );
  XNOR2_X1 U328 ( .A(n406), .B(KEYINPUT46), .ZN(n407) );
  INV_X1 U329 ( .A(KEYINPUT122), .ZN(n439) );
  XNOR2_X1 U330 ( .A(n439), .B(KEYINPUT54), .ZN(n440) );
  INV_X1 U331 ( .A(n448), .ZN(n381) );
  XNOR2_X1 U332 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U333 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U334 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U335 ( .A(n332), .B(n331), .ZN(n530) );
  XNOR2_X1 U336 ( .A(n461), .B(KEYINPUT58), .ZN(n462) );
  XNOR2_X1 U337 ( .A(n463), .B(n462), .ZN(G1351GAT) );
  INV_X1 U338 ( .A(KEYINPUT82), .ZN(n313) );
  XOR2_X1 U339 ( .A(G134GAT), .B(KEYINPUT81), .Z(n347) );
  XOR2_X1 U340 ( .A(KEYINPUT64), .B(KEYINPUT10), .Z(n295) );
  XNOR2_X1 U341 ( .A(KEYINPUT66), .B(KEYINPUT80), .ZN(n294) );
  XNOR2_X1 U342 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U343 ( .A(n347), .B(n296), .Z(n298) );
  NAND2_X1 U344 ( .A1(G232GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U345 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U346 ( .A(n299), .B(KEYINPUT9), .Z(n303) );
  XOR2_X1 U347 ( .A(G106GAT), .B(KEYINPUT75), .Z(n301) );
  XNOR2_X1 U348 ( .A(G99GAT), .B(G85GAT), .ZN(n300) );
  XNOR2_X1 U349 ( .A(n301), .B(n300), .ZN(n375) );
  XNOR2_X1 U350 ( .A(n375), .B(KEYINPUT11), .ZN(n302) );
  XOR2_X1 U351 ( .A(n303), .B(n302), .Z(n306) );
  XOR2_X1 U352 ( .A(KEYINPUT79), .B(G218GAT), .Z(n305) );
  XNOR2_X1 U353 ( .A(G50GAT), .B(G162GAT), .ZN(n304) );
  XNOR2_X1 U354 ( .A(n305), .B(n304), .ZN(n444) );
  XNOR2_X1 U355 ( .A(n306), .B(n444), .ZN(n312) );
  XOR2_X1 U356 ( .A(KEYINPUT8), .B(KEYINPUT73), .Z(n308) );
  XNOR2_X1 U357 ( .A(G43GAT), .B(G29GAT), .ZN(n307) );
  XNOR2_X1 U358 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U359 ( .A(KEYINPUT7), .B(n309), .Z(n403) );
  XNOR2_X1 U360 ( .A(G36GAT), .B(G190GAT), .ZN(n310) );
  XNOR2_X1 U361 ( .A(n310), .B(G92GAT), .ZN(n360) );
  XNOR2_X1 U362 ( .A(n403), .B(n360), .ZN(n311) );
  XNOR2_X1 U363 ( .A(n312), .B(n311), .ZN(n560) );
  XNOR2_X1 U364 ( .A(n313), .B(n560), .ZN(n431) );
  INV_X1 U365 ( .A(n431), .ZN(n477) );
  XOR2_X1 U366 ( .A(KEYINPUT91), .B(KEYINPUT65), .Z(n315) );
  XNOR2_X1 U367 ( .A(G183GAT), .B(KEYINPUT92), .ZN(n314) );
  XNOR2_X1 U368 ( .A(n315), .B(n314), .ZN(n321) );
  XOR2_X1 U369 ( .A(G120GAT), .B(G71GAT), .Z(n379) );
  XOR2_X1 U370 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n317) );
  XNOR2_X1 U371 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n316) );
  XNOR2_X1 U372 ( .A(n317), .B(n316), .ZN(n358) );
  XOR2_X1 U373 ( .A(n379), .B(n358), .Z(n319) );
  NAND2_X1 U374 ( .A1(G227GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U375 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U376 ( .A(n321), .B(n320), .ZN(n332) );
  XOR2_X1 U377 ( .A(G176GAT), .B(G190GAT), .Z(n323) );
  XNOR2_X1 U378 ( .A(G113GAT), .B(G134GAT), .ZN(n322) );
  XNOR2_X1 U379 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U380 ( .A(n324), .B(G99GAT), .Z(n326) );
  XOR2_X1 U381 ( .A(G15GAT), .B(G127GAT), .Z(n409) );
  XNOR2_X1 U382 ( .A(G43GAT), .B(n409), .ZN(n325) );
  XNOR2_X1 U383 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U384 ( .A(n327), .B(KEYINPUT20), .Z(n330) );
  XNOR2_X1 U385 ( .A(KEYINPUT89), .B(KEYINPUT0), .ZN(n328) );
  XNOR2_X1 U386 ( .A(n328), .B(KEYINPUT88), .ZN(n335) );
  XNOR2_X1 U387 ( .A(n335), .B(KEYINPUT90), .ZN(n329) );
  XNOR2_X1 U388 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U389 ( .A(G141GAT), .B(KEYINPUT3), .Z(n333) );
  XOR2_X1 U390 ( .A(KEYINPUT2), .B(n333), .Z(n443) );
  INV_X1 U391 ( .A(n443), .ZN(n334) );
  XOR2_X1 U392 ( .A(n335), .B(n334), .Z(n355) );
  XOR2_X1 U393 ( .A(G57GAT), .B(KEYINPUT5), .Z(n337) );
  XNOR2_X1 U394 ( .A(KEYINPUT6), .B(KEYINPUT4), .ZN(n336) );
  XNOR2_X1 U395 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U396 ( .A(G148GAT), .B(G155GAT), .Z(n339) );
  XNOR2_X1 U397 ( .A(G120GAT), .B(G127GAT), .ZN(n338) );
  XNOR2_X1 U398 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U399 ( .A(n341), .B(n340), .Z(n346) );
  XOR2_X1 U400 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n343) );
  NAND2_X1 U401 ( .A1(G225GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U402 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U403 ( .A(KEYINPUT97), .B(n344), .ZN(n345) );
  XNOR2_X1 U404 ( .A(n346), .B(n345), .ZN(n351) );
  XOR2_X1 U405 ( .A(KEYINPUT1), .B(G162GAT), .Z(n349) );
  XOR2_X1 U406 ( .A(G113GAT), .B(G1GAT), .Z(n389) );
  XNOR2_X1 U407 ( .A(n389), .B(n347), .ZN(n348) );
  XNOR2_X1 U408 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U409 ( .A(n351), .B(n350), .Z(n353) );
  XNOR2_X1 U410 ( .A(G29GAT), .B(G85GAT), .ZN(n352) );
  XNOR2_X1 U411 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U412 ( .A(n355), .B(n354), .ZN(n546) );
  XOR2_X1 U413 ( .A(G176GAT), .B(G64GAT), .Z(n378) );
  XOR2_X1 U414 ( .A(G211GAT), .B(KEYINPUT21), .Z(n357) );
  XNOR2_X1 U415 ( .A(G197GAT), .B(KEYINPUT94), .ZN(n356) );
  XNOR2_X1 U416 ( .A(n357), .B(n356), .ZN(n449) );
  XNOR2_X1 U417 ( .A(n358), .B(n449), .ZN(n365) );
  XOR2_X1 U418 ( .A(G204GAT), .B(KEYINPUT98), .Z(n363) );
  XNOR2_X1 U419 ( .A(G218GAT), .B(KEYINPUT99), .ZN(n359) );
  XOR2_X1 U420 ( .A(G8GAT), .B(G183GAT), .Z(n412) );
  XNOR2_X1 U421 ( .A(n359), .B(n412), .ZN(n361) );
  XNOR2_X1 U422 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U423 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U424 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U425 ( .A(n378), .B(n366), .Z(n368) );
  NAND2_X1 U426 ( .A1(G226GAT), .A2(G233GAT), .ZN(n367) );
  XOR2_X2 U427 ( .A(n368), .B(n367), .Z(n520) );
  INV_X1 U428 ( .A(n520), .ZN(n438) );
  XOR2_X1 U429 ( .A(KEYINPUT33), .B(KEYINPUT76), .Z(n370) );
  XNOR2_X1 U430 ( .A(G92GAT), .B(KEYINPUT78), .ZN(n369) );
  XOR2_X1 U431 ( .A(n370), .B(n369), .Z(n386) );
  XOR2_X1 U432 ( .A(KEYINPUT77), .B(KEYINPUT31), .Z(n372) );
  NAND2_X1 U433 ( .A1(G230GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U434 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U435 ( .A(n373), .B(KEYINPUT32), .Z(n377) );
  XNOR2_X1 U436 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n374) );
  XNOR2_X1 U437 ( .A(n374), .B(KEYINPUT74), .ZN(n413) );
  XNOR2_X1 U438 ( .A(n375), .B(n413), .ZN(n376) );
  XNOR2_X1 U439 ( .A(n377), .B(n376), .ZN(n384) );
  XNOR2_X1 U440 ( .A(n379), .B(n378), .ZN(n382) );
  XNOR2_X1 U441 ( .A(G148GAT), .B(G204GAT), .ZN(n380) );
  XNOR2_X1 U442 ( .A(n380), .B(G78GAT), .ZN(n448) );
  XNOR2_X1 U443 ( .A(n386), .B(n385), .ZN(n580) );
  XOR2_X1 U444 ( .A(n580), .B(KEYINPUT41), .Z(n554) );
  XOR2_X1 U445 ( .A(KEYINPUT72), .B(KEYINPUT30), .Z(n388) );
  XNOR2_X1 U446 ( .A(KEYINPUT69), .B(KEYINPUT29), .ZN(n387) );
  XNOR2_X1 U447 ( .A(n388), .B(n387), .ZN(n393) );
  XOR2_X1 U448 ( .A(G36GAT), .B(G50GAT), .Z(n391) );
  XNOR2_X1 U449 ( .A(n389), .B(G22GAT), .ZN(n390) );
  XNOR2_X1 U450 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U451 ( .A(n393), .B(n392), .Z(n395) );
  NAND2_X1 U452 ( .A1(G229GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U453 ( .A(n395), .B(n394), .ZN(n399) );
  XOR2_X1 U454 ( .A(G8GAT), .B(G197GAT), .Z(n397) );
  XNOR2_X1 U455 ( .A(G169GAT), .B(G141GAT), .ZN(n396) );
  XNOR2_X1 U456 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U457 ( .A(n399), .B(n398), .Z(n405) );
  XOR2_X1 U458 ( .A(KEYINPUT71), .B(G15GAT), .Z(n401) );
  XNOR2_X1 U459 ( .A(KEYINPUT70), .B(KEYINPUT68), .ZN(n400) );
  XNOR2_X1 U460 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U461 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U462 ( .A(n405), .B(n404), .Z(n549) );
  AND2_X1 U463 ( .A1(n554), .A2(n549), .ZN(n408) );
  XOR2_X1 U464 ( .A(G22GAT), .B(G155GAT), .Z(n453) );
  XOR2_X1 U465 ( .A(n453), .B(G64GAT), .Z(n411) );
  XNOR2_X1 U466 ( .A(G71GAT), .B(n409), .ZN(n410) );
  XNOR2_X1 U467 ( .A(n411), .B(n410), .ZN(n417) );
  XOR2_X1 U468 ( .A(n413), .B(n412), .Z(n415) );
  NAND2_X1 U469 ( .A1(G231GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U470 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U471 ( .A(n417), .B(n416), .Z(n419) );
  XNOR2_X1 U472 ( .A(G1GAT), .B(G211GAT), .ZN(n418) );
  XNOR2_X1 U473 ( .A(n419), .B(n418), .ZN(n427) );
  XOR2_X1 U474 ( .A(KEYINPUT86), .B(KEYINPUT84), .Z(n421) );
  XNOR2_X1 U475 ( .A(G78GAT), .B(KEYINPUT85), .ZN(n420) );
  XNOR2_X1 U476 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U477 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n423) );
  XNOR2_X1 U478 ( .A(KEYINPUT83), .B(KEYINPUT14), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U480 ( .A(n425), .B(n424), .Z(n426) );
  XOR2_X1 U481 ( .A(n427), .B(n426), .Z(n571) );
  NAND2_X1 U482 ( .A1(n571), .A2(n560), .ZN(n428) );
  OR2_X1 U483 ( .A1(n429), .A2(n428), .ZN(n430) );
  XNOR2_X1 U484 ( .A(n430), .B(KEYINPUT47), .ZN(n436) );
  XOR2_X1 U485 ( .A(KEYINPUT36), .B(n431), .Z(n588) );
  NOR2_X1 U486 ( .A1(n588), .A2(n571), .ZN(n432) );
  XNOR2_X1 U487 ( .A(KEYINPUT45), .B(n432), .ZN(n433) );
  INV_X1 U488 ( .A(n549), .ZN(n576) );
  NAND2_X1 U489 ( .A1(n433), .A2(n576), .ZN(n434) );
  NOR2_X1 U490 ( .A1(n434), .A2(n580), .ZN(n435) );
  NOR2_X1 U491 ( .A1(n436), .A2(n435), .ZN(n437) );
  XNOR2_X1 U492 ( .A(n437), .B(KEYINPUT48), .ZN(n548) );
  NOR2_X1 U493 ( .A1(n438), .A2(n548), .ZN(n441) );
  NOR2_X1 U494 ( .A1(n546), .A2(n442), .ZN(n575) );
  XOR2_X1 U495 ( .A(n444), .B(n443), .Z(n457) );
  XOR2_X1 U496 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n446) );
  NAND2_X1 U497 ( .A1(G228GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U498 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U499 ( .A(n447), .B(KEYINPUT23), .Z(n451) );
  XNOR2_X1 U500 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U501 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U502 ( .A(n452), .B(KEYINPUT93), .Z(n455) );
  XNOR2_X1 U503 ( .A(G106GAT), .B(n453), .ZN(n454) );
  XNOR2_X1 U504 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U505 ( .A(n457), .B(n456), .ZN(n470) );
  NAND2_X1 U506 ( .A1(n575), .A2(n470), .ZN(n459) );
  XOR2_X1 U507 ( .A(KEYINPUT55), .B(KEYINPUT123), .Z(n458) );
  XNOR2_X1 U508 ( .A(n459), .B(n458), .ZN(n460) );
  NAND2_X1 U509 ( .A1(n530), .A2(n460), .ZN(n570) );
  NOR2_X1 U510 ( .A1(n477), .A2(n570), .ZN(n463) );
  INV_X1 U511 ( .A(G190GAT), .ZN(n461) );
  NOR2_X1 U512 ( .A1(n576), .A2(n580), .ZN(n493) );
  XOR2_X1 U513 ( .A(n520), .B(KEYINPUT27), .Z(n468) );
  XNOR2_X1 U514 ( .A(KEYINPUT28), .B(KEYINPUT67), .ZN(n464) );
  XNOR2_X1 U515 ( .A(n464), .B(n470), .ZN(n526) );
  NOR2_X1 U516 ( .A1(n468), .A2(n526), .ZN(n465) );
  NAND2_X1 U517 ( .A1(n546), .A2(n465), .ZN(n529) );
  NOR2_X1 U518 ( .A1(n530), .A2(n529), .ZN(n476) );
  NOR2_X1 U519 ( .A1(n530), .A2(n470), .ZN(n466) );
  XOR2_X1 U520 ( .A(KEYINPUT100), .B(n466), .Z(n467) );
  XNOR2_X1 U521 ( .A(KEYINPUT26), .B(n467), .ZN(n573) );
  NOR2_X1 U522 ( .A1(n468), .A2(n573), .ZN(n545) );
  AND2_X1 U523 ( .A1(n520), .A2(n530), .ZN(n469) );
  XNOR2_X1 U524 ( .A(n469), .B(KEYINPUT101), .ZN(n471) );
  NAND2_X1 U525 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X1 U526 ( .A(KEYINPUT25), .B(n472), .ZN(n473) );
  NOR2_X1 U527 ( .A1(n545), .A2(n473), .ZN(n474) );
  NOR2_X1 U528 ( .A1(n546), .A2(n474), .ZN(n475) );
  NOR2_X1 U529 ( .A1(n476), .A2(n475), .ZN(n489) );
  XOR2_X1 U530 ( .A(KEYINPUT16), .B(KEYINPUT87), .Z(n479) );
  INV_X1 U531 ( .A(n571), .ZN(n585) );
  NAND2_X1 U532 ( .A1(n585), .A2(n477), .ZN(n478) );
  XNOR2_X1 U533 ( .A(n479), .B(n478), .ZN(n480) );
  NOR2_X1 U534 ( .A1(n489), .A2(n480), .ZN(n507) );
  AND2_X1 U535 ( .A1(n493), .A2(n507), .ZN(n486) );
  NAND2_X1 U536 ( .A1(n486), .A2(n546), .ZN(n481) );
  XNOR2_X1 U537 ( .A(n481), .B(KEYINPUT34), .ZN(n482) );
  XNOR2_X1 U538 ( .A(G1GAT), .B(n482), .ZN(G1324GAT) );
  NAND2_X1 U539 ( .A1(n520), .A2(n486), .ZN(n483) );
  XNOR2_X1 U540 ( .A(n483), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U541 ( .A(G15GAT), .B(KEYINPUT35), .Z(n485) );
  NAND2_X1 U542 ( .A1(n486), .A2(n530), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n485), .B(n484), .ZN(G1326GAT) );
  NAND2_X1 U544 ( .A1(n526), .A2(n486), .ZN(n487) );
  XNOR2_X1 U545 ( .A(n487), .B(KEYINPUT102), .ZN(n488) );
  XNOR2_X1 U546 ( .A(G22GAT), .B(n488), .ZN(G1327GAT) );
  XOR2_X1 U547 ( .A(G29GAT), .B(KEYINPUT39), .Z(n497) );
  NOR2_X1 U548 ( .A1(n489), .A2(n585), .ZN(n490) );
  XNOR2_X1 U549 ( .A(n490), .B(KEYINPUT103), .ZN(n491) );
  NOR2_X1 U550 ( .A1(n588), .A2(n491), .ZN(n492) );
  XOR2_X1 U551 ( .A(KEYINPUT37), .B(n492), .Z(n518) );
  NAND2_X1 U552 ( .A1(n518), .A2(n493), .ZN(n495) );
  XOR2_X1 U553 ( .A(KEYINPUT38), .B(KEYINPUT104), .Z(n494) );
  XNOR2_X1 U554 ( .A(n495), .B(n494), .ZN(n503) );
  NAND2_X1 U555 ( .A1(n503), .A2(n546), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n497), .B(n496), .ZN(G1328GAT) );
  NAND2_X1 U557 ( .A1(n503), .A2(n520), .ZN(n498) );
  XNOR2_X1 U558 ( .A(G36GAT), .B(n498), .ZN(G1329GAT) );
  XNOR2_X1 U559 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n502) );
  XOR2_X1 U560 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n500) );
  NAND2_X1 U561 ( .A1(n503), .A2(n530), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U563 ( .A(n502), .B(n501), .ZN(G1330GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n505) );
  NAND2_X1 U565 ( .A1(n503), .A2(n526), .ZN(n504) );
  XNOR2_X1 U566 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U567 ( .A(G50GAT), .B(n506), .ZN(G1331GAT) );
  INV_X1 U568 ( .A(n554), .ZN(n564) );
  NOR2_X1 U569 ( .A1(n549), .A2(n564), .ZN(n517) );
  AND2_X1 U570 ( .A1(n517), .A2(n507), .ZN(n513) );
  NAND2_X1 U571 ( .A1(n546), .A2(n513), .ZN(n508) );
  XNOR2_X1 U572 ( .A(KEYINPUT42), .B(n508), .ZN(n509) );
  XNOR2_X1 U573 ( .A(G57GAT), .B(n509), .ZN(G1332GAT) );
  XOR2_X1 U574 ( .A(G64GAT), .B(KEYINPUT109), .Z(n511) );
  NAND2_X1 U575 ( .A1(n513), .A2(n520), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(G1333GAT) );
  NAND2_X1 U577 ( .A1(n513), .A2(n530), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n512), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n515) );
  NAND2_X1 U580 ( .A1(n513), .A2(n526), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U582 ( .A(G78GAT), .B(n516), .ZN(G1335GAT) );
  AND2_X1 U583 ( .A1(n518), .A2(n517), .ZN(n525) );
  NAND2_X1 U584 ( .A1(n525), .A2(n546), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n519), .B(G85GAT), .ZN(G1336GAT) );
  XOR2_X1 U586 ( .A(G92GAT), .B(KEYINPUT111), .Z(n522) );
  NAND2_X1 U587 ( .A1(n525), .A2(n520), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n522), .B(n521), .ZN(G1337GAT) );
  NAND2_X1 U589 ( .A1(n525), .A2(n530), .ZN(n523) );
  XNOR2_X1 U590 ( .A(n523), .B(KEYINPUT112), .ZN(n524) );
  XNOR2_X1 U591 ( .A(G99GAT), .B(n524), .ZN(G1338GAT) );
  NAND2_X1 U592 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n527), .B(KEYINPUT44), .ZN(n528) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  XOR2_X1 U595 ( .A(G113GAT), .B(KEYINPUT115), .Z(n534) );
  NOR2_X1 U596 ( .A1(n548), .A2(n529), .ZN(n531) );
  NAND2_X1 U597 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U598 ( .A(KEYINPUT114), .B(n532), .Z(n541) );
  NAND2_X1 U599 ( .A1(n541), .A2(n549), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(G1340GAT) );
  XOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT49), .Z(n536) );
  NAND2_X1 U602 ( .A1(n554), .A2(n541), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n536), .B(n535), .ZN(G1341GAT) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(KEYINPUT116), .ZN(n540) );
  XOR2_X1 U605 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n538) );
  NAND2_X1 U606 ( .A1(n541), .A2(n585), .ZN(n537) );
  XNOR2_X1 U607 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U608 ( .A(n540), .B(n539), .ZN(G1342GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n543) );
  NAND2_X1 U610 ( .A1(n431), .A2(n541), .ZN(n542) );
  XNOR2_X1 U611 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U612 ( .A(G134GAT), .B(n544), .ZN(G1343GAT) );
  NAND2_X1 U613 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n558) );
  NAND2_X1 U615 ( .A1(n549), .A2(n558), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n550), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n552) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U620 ( .A(KEYINPUT119), .B(n553), .Z(n556) );
  NAND2_X1 U621 ( .A1(n558), .A2(n554), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1345GAT) );
  NAND2_X1 U623 ( .A1(n585), .A2(n558), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n557), .B(G155GAT), .ZN(G1346GAT) );
  INV_X1 U625 ( .A(n558), .ZN(n559) );
  NOR2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n562) );
  XNOR2_X1 U627 ( .A(G162GAT), .B(KEYINPUT121), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1347GAT) );
  NOR2_X1 U629 ( .A1(n576), .A2(n570), .ZN(n563) );
  XOR2_X1 U630 ( .A(G169GAT), .B(n563), .Z(G1348GAT) );
  NOR2_X1 U631 ( .A1(n570), .A2(n564), .ZN(n569) );
  XOR2_X1 U632 ( .A(KEYINPUT57), .B(KEYINPUT125), .Z(n566) );
  XNOR2_X1 U633 ( .A(G176GAT), .B(KEYINPUT124), .ZN(n565) );
  XNOR2_X1 U634 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U635 ( .A(KEYINPUT56), .B(n567), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(G1349GAT) );
  NOR2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U638 ( .A(G183GAT), .B(n572), .Z(G1350GAT) );
  INV_X1 U639 ( .A(n573), .ZN(n574) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n587) );
  NOR2_X1 U641 ( .A1(n576), .A2(n587), .ZN(n578) );
  XNOR2_X1 U642 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(n579), .ZN(G1352GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n582) );
  INV_X1 U646 ( .A(n587), .ZN(n584) );
  NAND2_X1 U647 ( .A1(n584), .A2(n580), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U649 ( .A(G204GAT), .B(n583), .ZN(G1353GAT) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n586), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n590) );
  XNOR2_X1 U653 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

