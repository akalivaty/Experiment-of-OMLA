//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 1 1 1 0 1 1 0 0 1 0 1 0 0 1 1 0 0 1 1 1 1 1 0 1 1 0 0 0 0 0 0 0 0 1 0 1 0 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n567, new_n569, new_n570, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n624, new_n627, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1185, new_n1186;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT68), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n463), .A2(KEYINPUT3), .A3(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n465), .A2(G137), .A3(new_n466), .A4(new_n468), .ZN(new_n469));
  AOI21_X1  g044(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n469), .A2(KEYINPUT69), .A3(new_n471), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n468), .A2(new_n477), .A3(G125), .ZN(new_n478));
  INV_X1    g053(.A(G113), .ZN(new_n479));
  OAI21_X1  g054(.A(KEYINPUT66), .B1(new_n479), .B2(new_n462), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n481), .A2(G113), .A3(G2104), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n478), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  AND3_X1   g058(.A1(new_n483), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n484));
  AOI21_X1  g059(.A(KEYINPUT67), .B1(new_n483), .B2(G2105), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n476), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT70), .ZN(G160));
  AND2_X1   g063(.A1(new_n465), .A2(new_n468), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(new_n466), .ZN(new_n490));
  INV_X1    g065(.A(G136), .ZN(new_n491));
  AND2_X1   g066(.A1(G112), .A2(G2105), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n492), .B1(G100), .B2(new_n466), .ZN(new_n493));
  OAI22_X1  g068(.A1(new_n490), .A2(new_n491), .B1(new_n462), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n489), .A2(KEYINPUT71), .A3(G2105), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT71), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n465), .A2(new_n468), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(new_n466), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n494), .B1(G124), .B2(new_n499), .ZN(G162));
  AND2_X1   g075(.A1(KEYINPUT4), .A2(G138), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n465), .A2(new_n468), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(G102), .A2(G2104), .ZN(new_n503));
  AOI21_X1  g078(.A(G2105), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n465), .A2(G126), .A3(new_n468), .ZN(new_n505));
  NAND2_X1  g080(.A1(G114), .A2(G2104), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n466), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n468), .A2(new_n477), .A3(G138), .A4(new_n466), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NOR3_X1   g085(.A1(new_n504), .A2(new_n507), .A3(new_n510), .ZN(G164));
  XOR2_X1   g086(.A(KEYINPUT5), .B(G543), .Z(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT72), .A2(G651), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT72), .A2(G651), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT6), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n512), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT73), .B(G88), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n522), .B1(new_n518), .B2(new_n514), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G50), .ZN(new_n524));
  NAND2_X1  g099(.A1(G75), .A2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G62), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n512), .B2(new_n526), .ZN(new_n527));
  OR2_X1    g102(.A1(KEYINPUT72), .A2(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(new_n515), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n521), .A2(new_n524), .A3(new_n530), .ZN(G303));
  INV_X1    g106(.A(G303), .ZN(G166));
  NAND2_X1  g107(.A1(new_n519), .A2(G89), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n523), .A2(G51), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n537));
  OR2_X1    g112(.A1(KEYINPUT5), .A2(G543), .ZN(new_n538));
  NAND2_X1  g113(.A1(KEYINPUT5), .A2(G543), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AND2_X1   g115(.A1(G63), .A2(G651), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n536), .A2(new_n537), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n533), .A2(new_n534), .A3(new_n542), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(KEYINPUT74), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(KEYINPUT74), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(G168));
  XNOR2_X1  g121(.A(KEYINPUT75), .B(G90), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n519), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n523), .A2(G52), .ZN(new_n549));
  NAND2_X1  g124(.A1(G77), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G64), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n512), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(new_n529), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n548), .A2(new_n549), .A3(new_n553), .ZN(G301));
  INV_X1    g129(.A(G301), .ZN(G171));
  XOR2_X1   g130(.A(KEYINPUT77), .B(G81), .Z(new_n556));
  NAND2_X1  g131(.A1(new_n519), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g132(.A(KEYINPUT76), .B(G43), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n523), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(G68), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G56), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n512), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(new_n529), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n557), .A2(new_n559), .A3(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  AND3_X1   g141(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G36), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n567), .A2(new_n570), .ZN(G188));
  NAND2_X1  g146(.A1(new_n523), .A2(G53), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT9), .ZN(new_n573));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  XNOR2_X1  g149(.A(KEYINPUT78), .B(G65), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n512), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n519), .A2(G91), .B1(new_n576), .B2(G651), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n573), .A2(new_n577), .ZN(G299));
  XOR2_X1   g153(.A(new_n543), .B(KEYINPUT74), .Z(G286));
  NAND2_X1  g154(.A1(new_n523), .A2(G49), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n518), .A2(new_n514), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n581), .A2(G87), .A3(new_n540), .ZN(new_n582));
  INV_X1    g157(.A(G651), .ZN(new_n583));
  INV_X1    g158(.A(G74), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n583), .B1(new_n512), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(new_n586));
  AND4_X1   g161(.A1(KEYINPUT79), .A2(new_n580), .A3(new_n582), .A4(new_n586), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n585), .B1(new_n523), .B2(G49), .ZN(new_n588));
  AOI21_X1  g163(.A(KEYINPUT79), .B1(new_n588), .B2(new_n582), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n587), .A2(new_n589), .ZN(G288));
  INV_X1    g165(.A(KEYINPUT6), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n591), .B1(new_n528), .B2(new_n515), .ZN(new_n592));
  OAI211_X1 g167(.A(G48), .B(G543), .C1(new_n592), .C2(new_n513), .ZN(new_n593));
  OAI211_X1 g168(.A(G86), .B(new_n540), .C1(new_n592), .C2(new_n513), .ZN(new_n594));
  INV_X1    g169(.A(G61), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n595), .B1(new_n538), .B2(new_n539), .ZN(new_n596));
  AND2_X1   g171(.A1(G73), .A2(G543), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n529), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n593), .A2(new_n594), .A3(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT80), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n599), .B(new_n600), .ZN(G305));
  NAND2_X1  g176(.A1(G72), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G60), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n512), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(new_n529), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT81), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n519), .A2(G85), .B1(new_n523), .B2(G47), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(G290));
  XNOR2_X1  g183(.A(KEYINPUT82), .B(KEYINPUT10), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n581), .A2(new_n540), .ZN(new_n611));
  INV_X1    g186(.A(G92), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(G79), .A2(G543), .ZN(new_n614));
  INV_X1    g189(.A(G66), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n512), .B2(new_n615), .ZN(new_n616));
  AOI22_X1  g191(.A1(G54), .A2(new_n523), .B1(new_n616), .B2(G651), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n519), .A2(G92), .A3(new_n609), .ZN(new_n618));
  AND3_X1   g193(.A1(new_n613), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(new_n620));
  MUX2_X1   g195(.A(new_n620), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g196(.A(new_n620), .B(G301), .S(G868), .Z(G321));
  NAND2_X1  g197(.A1(G286), .A2(G868), .ZN(new_n623));
  AND2_X1   g198(.A1(new_n573), .A2(new_n577), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(G868), .B2(new_n624), .ZN(G297));
  OAI21_X1  g200(.A(new_n623), .B1(G868), .B2(new_n624), .ZN(G280));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n619), .B1(new_n627), .B2(G860), .ZN(G148));
  NAND2_X1  g203(.A1(new_n619), .A2(new_n627), .ZN(new_n629));
  MUX2_X1   g204(.A(new_n564), .B(new_n629), .S(G868), .Z(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g206(.A1(new_n468), .A2(new_n477), .ZN(new_n632));
  AOI211_X1 g207(.A(G2105), .B(new_n632), .C1(new_n463), .C2(new_n464), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT12), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT13), .ZN(new_n635));
  XOR2_X1   g210(.A(KEYINPUT83), .B(G2100), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n499), .A2(G123), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT84), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n497), .A2(G2105), .ZN(new_n640));
  MUX2_X1   g215(.A(G99), .B(G111), .S(G2105), .Z(new_n641));
  AOI22_X1  g216(.A1(new_n640), .A2(G135), .B1(G2104), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(G2096), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n643), .A2(G2096), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n637), .A2(new_n646), .A3(new_n647), .ZN(G156));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XOR2_X1   g225(.A(G2443), .B(G2446), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G1341), .B(G1348), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(KEYINPUT14), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT15), .B(G2435), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT85), .B(G2438), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2427), .B(G2430), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n655), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n660), .B1(new_n658), .B2(new_n659), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n654), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n654), .A2(new_n661), .ZN(new_n663));
  AND3_X1   g238(.A1(new_n662), .A2(G14), .A3(new_n663), .ZN(G401));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2072), .B(G2078), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT87), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n668), .B(KEYINPUT17), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(new_n667), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n669), .A2(new_n670), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n671), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT88), .ZN(new_n676));
  OR3_X1    g251(.A1(new_n672), .A2(new_n667), .A3(new_n666), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n665), .A2(new_n667), .A3(new_n668), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT86), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT18), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n676), .A2(new_n677), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(new_n645), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(G2100), .ZN(G227));
  XOR2_X1   g258(.A(G1961), .B(G1966), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT89), .ZN(new_n685));
  XOR2_X1   g260(.A(G1956), .B(G2474), .Z(new_n686));
  OR2_X1    g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1971), .B(G1976), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT19), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n685), .A2(new_n686), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n691), .A2(new_n689), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT90), .B(KEYINPUT20), .Z(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n690), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n687), .A2(new_n689), .A3(new_n691), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n695), .B(new_n696), .C1(new_n692), .C2(new_n694), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1981), .B(G1986), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT91), .ZN(new_n701));
  XOR2_X1   g276(.A(G1991), .B(G1996), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n699), .B(new_n703), .ZN(G229));
  OR2_X1    g279(.A1(G16), .A2(G24), .ZN(new_n705));
  INV_X1    g280(.A(G16), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(G290), .B2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(G1986), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT96), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(new_n707), .B2(new_n708), .ZN(new_n711));
  MUX2_X1   g286(.A(G6), .B(G305), .S(G16), .Z(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT32), .B(G1981), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n588), .A2(new_n582), .ZN(new_n715));
  MUX2_X1   g290(.A(G23), .B(new_n715), .S(G16), .Z(new_n716));
  XOR2_X1   g291(.A(KEYINPUT33), .B(G1976), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(G16), .A2(G22), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G166), .B2(G16), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(G1971), .ZN(new_n721));
  NOR3_X1   g296(.A1(new_n714), .A2(new_n718), .A3(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT34), .ZN(new_n723));
  AOI211_X1 g298(.A(new_n709), .B(new_n711), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(G25), .A2(G29), .ZN(new_n725));
  MUX2_X1   g300(.A(G95), .B(G107), .S(G2105), .Z(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G2104), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT93), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n489), .A2(G131), .A3(new_n466), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(KEYINPUT92), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT92), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n640), .A2(new_n731), .A3(G131), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n728), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT94), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n499), .A2(G119), .ZN(new_n735));
  AND3_X1   g310(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n734), .B1(new_n733), .B2(new_n735), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n725), .B1(new_n738), .B2(G29), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT95), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT35), .B(G1991), .Z(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n724), .B(new_n742), .C1(new_n723), .C2(new_n722), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT36), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(new_n744), .ZN(new_n746));
  NOR2_X1   g321(.A1(G16), .A2(G19), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n565), .B2(G16), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT97), .Z(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G1341), .ZN(new_n750));
  INV_X1    g325(.A(G29), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G32), .ZN(new_n752));
  NAND3_X1  g327(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT26), .Z(new_n754));
  INV_X1    g329(.A(G141), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n754), .B1(new_n490), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n470), .A2(G105), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT101), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(G129), .ZN(new_n760));
  INV_X1    g335(.A(new_n499), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n752), .B1(new_n763), .B2(new_n751), .ZN(new_n764));
  XOR2_X1   g339(.A(KEYINPUT27), .B(G1996), .Z(new_n765));
  NOR2_X1   g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n766), .A2(KEYINPUT102), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(KEYINPUT102), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n750), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT31), .B(G11), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT30), .B(G28), .Z(new_n771));
  NOR2_X1   g346(.A1(G171), .A2(new_n706), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G5), .B2(new_n706), .ZN(new_n773));
  INV_X1    g348(.A(G1961), .ZN(new_n774));
  OAI221_X1 g349(.A(new_n770), .B1(G29), .B2(new_n771), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n774), .B2(new_n773), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n751), .A2(G33), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT25), .Z(new_n779));
  AND2_X1   g354(.A1(new_n468), .A2(new_n477), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n780), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n779), .B1(new_n781), .B2(new_n466), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G139), .B2(new_n640), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT100), .Z(new_n784));
  OAI21_X1  g359(.A(new_n777), .B1(new_n784), .B2(new_n751), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G2072), .ZN(new_n786));
  NOR2_X1   g361(.A1(G27), .A2(G29), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G164), .B2(G29), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G2078), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  AOI22_X1  g365(.A1(new_n644), .A2(G29), .B1(new_n764), .B2(new_n765), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n769), .A2(new_n776), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(G29), .A2(G35), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G162), .B2(G29), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT29), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G2090), .ZN(new_n796));
  NAND2_X1  g371(.A1(G168), .A2(G16), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G16), .B2(G21), .ZN(new_n798));
  INV_X1    g373(.A(G1966), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT103), .ZN(new_n801));
  NAND2_X1  g376(.A1(G160), .A2(G29), .ZN(new_n802));
  AND2_X1   g377(.A1(KEYINPUT24), .A2(G34), .ZN(new_n803));
  NOR2_X1   g378(.A1(KEYINPUT24), .A2(G34), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n751), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G2084), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n796), .A2(new_n801), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n706), .A2(G20), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT104), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT23), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(G299), .B2(G16), .ZN(new_n812));
  INV_X1    g387(.A(G1956), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(new_n798), .B2(new_n799), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n751), .A2(G26), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT28), .Z(new_n817));
  NAND2_X1  g392(.A1(new_n466), .A2(G104), .ZN(new_n818));
  NAND2_X1  g393(.A1(G116), .A2(G2105), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n462), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT98), .ZN(new_n821));
  INV_X1    g396(.A(G140), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n821), .B1(new_n490), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n640), .A2(KEYINPUT98), .A3(G140), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n820), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AND3_X1   g400(.A1(new_n499), .A2(KEYINPUT99), .A3(G128), .ZN(new_n826));
  AOI21_X1  g401(.A(KEYINPUT99), .B1(new_n499), .B2(G128), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n817), .B1(new_n828), .B2(G29), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(G2067), .ZN(new_n830));
  NOR2_X1   g405(.A1(G4), .A2(G16), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(new_n619), .B2(G16), .ZN(new_n832));
  INV_X1    g407(.A(G1348), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n815), .A2(new_n830), .A3(new_n834), .ZN(new_n835));
  NOR3_X1   g410(.A1(new_n792), .A2(new_n808), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n745), .A2(new_n746), .A3(new_n836), .ZN(G150));
  INV_X1    g412(.A(G150), .ZN(G311));
  NAND2_X1  g413(.A1(new_n519), .A2(G93), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n523), .A2(G55), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n516), .A2(new_n517), .ZN(new_n841));
  AOI22_X1  g416(.A1(new_n540), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n839), .B(new_n840), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(KEYINPUT105), .B(G860), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT37), .Z(new_n847));
  XNOR2_X1  g422(.A(new_n565), .B(new_n843), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT38), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n620), .A2(new_n627), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  AND2_X1   g427(.A1(new_n852), .A2(KEYINPUT39), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n844), .B1(new_n852), .B2(KEYINPUT39), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n847), .B1(new_n853), .B2(new_n854), .ZN(G145));
  INV_X1    g430(.A(KEYINPUT108), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n828), .B(G164), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT106), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n859), .B1(new_n736), .B2(new_n737), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n733), .A2(new_n735), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(KEYINPUT94), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n862), .A2(KEYINPUT106), .A3(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(G142), .ZN(new_n865));
  AND2_X1   g440(.A1(G118), .A2(G2105), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n866), .B1(G106), .B2(new_n466), .ZN(new_n867));
  OAI22_X1  g442(.A1(new_n490), .A2(new_n865), .B1(new_n462), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n868), .B1(G130), .B2(new_n499), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n634), .ZN(new_n870));
  AND3_X1   g445(.A1(new_n860), .A2(new_n864), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n870), .B1(new_n860), .B2(new_n864), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n858), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n870), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n736), .A2(new_n737), .A3(new_n859), .ZN(new_n875));
  AOI21_X1  g450(.A(KEYINPUT106), .B1(new_n862), .B2(new_n863), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n860), .A2(new_n864), .A3(new_n870), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n877), .A2(new_n878), .A3(new_n857), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n873), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n784), .B(new_n762), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(G160), .B(G162), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n644), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT107), .ZN(new_n885));
  INV_X1    g460(.A(new_n881), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n873), .A2(new_n879), .A3(new_n886), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n882), .A2(new_n884), .A3(new_n885), .A4(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(G37), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(KEYINPUT107), .B1(new_n880), .B2(new_n881), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n884), .B1(new_n891), .B2(new_n887), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n856), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n882), .A2(new_n885), .A3(new_n887), .ZN(new_n894));
  INV_X1    g469(.A(new_n884), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n896), .A2(KEYINPUT108), .A3(new_n889), .A4(new_n888), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n893), .A2(KEYINPUT40), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT40), .B1(new_n893), .B2(new_n897), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(G395));
  NOR2_X1   g475(.A1(new_n843), .A2(G868), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n629), .B(KEYINPUT109), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(new_n848), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n624), .A2(new_n620), .ZN(new_n904));
  NAND2_X1  g479(.A1(G299), .A2(new_n619), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT41), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT110), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(G299), .A2(KEYINPUT110), .A3(new_n619), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n910), .A2(KEYINPUT41), .A3(new_n911), .A4(new_n904), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n903), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n910), .A2(new_n911), .A3(new_n904), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n903), .A2(new_n916), .ZN(new_n917));
  OR3_X1    g492(.A1(new_n914), .A2(new_n917), .A3(KEYINPUT42), .ZN(new_n918));
  OAI21_X1  g493(.A(KEYINPUT42), .B1(new_n914), .B2(new_n917), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(G290), .B(new_n715), .ZN(new_n921));
  XNOR2_X1  g496(.A(G305), .B(G166), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n921), .B(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n920), .B(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n901), .B1(new_n925), .B2(G868), .ZN(G295));
  AOI21_X1  g501(.A(new_n901), .B1(new_n925), .B2(G868), .ZN(G331));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT111), .ZN(new_n929));
  INV_X1    g504(.A(new_n848), .ZN(new_n930));
  NOR2_X1   g505(.A1(G168), .A2(G171), .ZN(new_n931));
  AOI21_X1  g506(.A(G301), .B1(new_n544), .B2(new_n545), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(G286), .A2(G301), .ZN(new_n934));
  INV_X1    g509(.A(new_n932), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n934), .A2(new_n935), .A3(new_n848), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n913), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n933), .A2(new_n936), .A3(new_n915), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n929), .B1(new_n940), .B2(new_n924), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n938), .A2(new_n939), .ZN(new_n942));
  NOR3_X1   g517(.A1(new_n942), .A2(KEYINPUT111), .A3(new_n923), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n907), .B1(new_n933), .B2(new_n936), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n945), .A2(new_n906), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n923), .B1(new_n945), .B2(new_n915), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT112), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  OR2_X1    g523(.A1(new_n945), .A2(new_n915), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT112), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n945), .A2(new_n906), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n949), .A2(new_n950), .A3(new_n923), .A4(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n948), .A2(new_n952), .A3(new_n889), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n928), .B1(new_n944), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n955));
  AOI21_X1  g530(.A(G37), .B1(new_n942), .B2(new_n923), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n956), .B(KEYINPUT43), .C1(new_n941), .C2(new_n943), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n954), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT113), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT113), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n954), .A2(new_n960), .A3(new_n957), .A4(new_n955), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT43), .B1(new_n944), .B2(new_n953), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n956), .B(new_n928), .C1(new_n941), .C2(new_n943), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n962), .A2(KEYINPUT44), .A3(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n959), .A2(new_n961), .A3(new_n964), .ZN(G397));
  INV_X1    g540(.A(KEYINPUT127), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT115), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n828), .A2(G2067), .ZN(new_n968));
  INV_X1    g543(.A(G2067), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n969), .B(new_n825), .C1(new_n826), .C2(new_n827), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT45), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n972), .B1(G164), .B2(G1384), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n483), .A2(G2105), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT67), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n483), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n978), .A2(G40), .A3(new_n474), .A4(new_n475), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n973), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n971), .A2(KEYINPUT114), .A3(new_n980), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n762), .B(G1996), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n980), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT114), .B1(new_n971), .B2(new_n980), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n967), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n985), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n987), .A2(KEYINPUT115), .A3(new_n981), .A4(new_n983), .ZN(new_n988));
  AND2_X1   g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n738), .A2(new_n741), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n738), .A2(new_n741), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n980), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(G290), .A2(G1986), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n708), .B1(new_n606), .B2(new_n607), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n980), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n989), .A2(new_n992), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(G303), .A2(G8), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n997), .B(KEYINPUT55), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n502), .A2(new_n503), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(new_n466), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n505), .A2(new_n506), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(G2105), .ZN(new_n1002));
  INV_X1    g577(.A(new_n510), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1000), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G1384), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1004), .A2(KEYINPUT45), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT116), .ZN(new_n1007));
  INV_X1    g582(.A(G40), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n476), .A2(new_n486), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n510), .B1(new_n1001), .B2(G2105), .ZN(new_n1010));
  AOI21_X1  g585(.A(G1384), .B1(new_n1010), .B2(new_n1000), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT116), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1011), .A2(new_n1012), .A3(KEYINPUT45), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1007), .A2(new_n1009), .A3(new_n973), .A4(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G1971), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT50), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1016), .B1(G164), .B2(G1384), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1004), .A2(KEYINPUT50), .A3(new_n1005), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n979), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  XOR2_X1   g594(.A(KEYINPUT117), .B(G2090), .Z(new_n1020));
  AOI22_X1  g595(.A1(new_n1014), .A2(new_n1015), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G8), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n998), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n998), .ZN(new_n1024));
  NOR4_X1   g599(.A1(G164), .A2(KEYINPUT116), .A3(new_n972), .A4(G1384), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1012), .B1(new_n1011), .B2(KEYINPUT45), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1011), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n979), .B1(new_n1028), .B2(new_n972), .ZN(new_n1029));
  AOI21_X1  g604(.A(G1971), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  AND2_X1   g605(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1031));
  OAI211_X1 g606(.A(G8), .B(new_n1024), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1022), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1033));
  INV_X1    g608(.A(G1976), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT52), .B1(G288), .B2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n588), .A2(G1976), .A3(new_n582), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n1036), .B(KEYINPUT118), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1033), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n599), .A2(G1981), .ZN(new_n1039));
  INV_X1    g614(.A(G1981), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n593), .A2(new_n594), .A3(new_n1040), .A4(new_n598), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1039), .A2(KEYINPUT49), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT119), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1039), .A2(KEYINPUT119), .A3(KEYINPUT49), .A4(new_n1041), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT49), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1033), .A2(new_n1046), .A3(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(G8), .B1(new_n1028), .B2(new_n979), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n1052));
  XNOR2_X1  g627(.A(new_n1036), .B(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT52), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  AND3_X1   g629(.A1(new_n1038), .A2(new_n1050), .A3(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1009), .A2(new_n973), .A3(new_n1006), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n799), .ZN(new_n1057));
  XNOR2_X1  g632(.A(KEYINPUT120), .B(G2084), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT50), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1059));
  AOI211_X1 g634(.A(new_n1016), .B(G1384), .C1(new_n1010), .C2(new_n1000), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1009), .B(new_n1058), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1061));
  AOI211_X1 g636(.A(new_n1022), .B(G286), .C1(new_n1057), .C2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1023), .A2(new_n1032), .A3(new_n1055), .A4(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT63), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1011), .A2(KEYINPUT45), .ZN(new_n1066));
  AOI211_X1 g641(.A(new_n972), .B(G1384), .C1(new_n1010), .C2(new_n1000), .ZN(new_n1067));
  NOR3_X1   g642(.A1(new_n1066), .A2(new_n1067), .A3(new_n979), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1061), .B1(new_n1068), .B2(G1966), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1069), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1022), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1070), .B1(new_n1024), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT121), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1055), .B(new_n1075), .C1(new_n1073), .C2(new_n1024), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1075), .B1(new_n1023), .B2(new_n1055), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1065), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n544), .A2(G8), .A3(new_n545), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT125), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n1082), .A2(KEYINPUT51), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1019), .A2(new_n1058), .B1(new_n1056), .B2(new_n799), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1080), .B(new_n1083), .C1(new_n1084), .C2(new_n1022), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1082), .A2(KEYINPUT51), .ZN(new_n1086));
  OAI211_X1 g661(.A(G8), .B(new_n1086), .C1(new_n1069), .C2(G286), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1069), .A2(G8), .A3(G286), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1085), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT62), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n1023), .A2(new_n1032), .A3(new_n1055), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1092), .B1(new_n1014), .B2(G2078), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1092), .A2(G2078), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1009), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1095));
  AOI22_X1  g670(.A1(new_n1068), .A2(new_n1094), .B1(new_n1095), .B2(new_n774), .ZN(new_n1096));
  AOI21_X1  g671(.A(G301), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT62), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1085), .A2(new_n1087), .A3(new_n1098), .A4(new_n1088), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1090), .A2(new_n1091), .A3(new_n1097), .A4(new_n1099), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1050), .B(new_n1034), .C1(new_n589), .C2(new_n587), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1051), .B1(new_n1101), .B2(new_n1041), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1032), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1102), .B1(new_n1103), .B2(new_n1055), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1079), .A2(new_n1100), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT122), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1106), .B1(new_n1019), .B2(G1956), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1095), .A2(KEYINPUT122), .A3(new_n813), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT56), .B(G2072), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1029), .A2(new_n1007), .A3(new_n1013), .A4(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1107), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n624), .B(KEYINPUT57), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1112), .A2(new_n1107), .A3(new_n1110), .A4(new_n1108), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT61), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1028), .A2(new_n979), .ZN(new_n1119));
  XNOR2_X1  g694(.A(KEYINPUT58), .B(G1341), .ZN(new_n1120));
  OAI22_X1  g695(.A1(new_n1014), .A2(G1996), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT124), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1121), .A2(new_n1122), .A3(new_n565), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT59), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT59), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1121), .A2(new_n1122), .A3(new_n1125), .A4(new_n565), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n487), .A2(G40), .A3(new_n969), .A4(new_n1011), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT123), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1009), .A2(KEYINPUT123), .A3(new_n969), .A4(new_n1011), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1019), .A2(G1348), .ZN(new_n1133));
  OR2_X1    g708(.A1(new_n620), .A2(KEYINPUT60), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n619), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1095), .A2(new_n833), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1137), .A2(new_n620), .A3(new_n1130), .A4(new_n1131), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1135), .B1(new_n1139), .B2(KEYINPUT60), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1114), .A2(KEYINPUT61), .A3(new_n1115), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1118), .A2(new_n1127), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1115), .B(new_n619), .C1(new_n1133), .C2(new_n1132), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n1143), .A2(new_n1114), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT54), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n974), .A2(G40), .A3(new_n1094), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n1066), .A2(new_n476), .A3(new_n1147), .ZN(new_n1148));
  AOI22_X1  g723(.A1(new_n1027), .A2(new_n1148), .B1(new_n1095), .B2(new_n774), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1149), .A2(new_n1093), .A3(G301), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1146), .B1(new_n1150), .B2(new_n1097), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1093), .A2(new_n1096), .A3(G301), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1149), .A2(new_n1093), .ZN(new_n1153));
  OAI211_X1 g728(.A(KEYINPUT54), .B(new_n1152), .C1(new_n1153), .C2(G301), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1091), .A2(new_n1151), .A3(new_n1154), .A4(new_n1089), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1145), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n996), .B1(new_n1105), .B2(new_n1157), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n973), .A2(G1996), .A3(new_n979), .ZN(new_n1159));
  XOR2_X1   g734(.A(new_n1159), .B(KEYINPUT46), .Z(new_n1160));
  OAI21_X1  g735(.A(new_n980), .B1(new_n971), .B2(new_n762), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT47), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n980), .A2(new_n993), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1164), .B(KEYINPUT48), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n989), .A2(new_n992), .A3(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n986), .A2(new_n988), .A3(new_n990), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT126), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1167), .A2(new_n1168), .A3(new_n970), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n980), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1168), .B1(new_n1167), .B2(new_n970), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1163), .B(new_n1166), .C1(new_n1170), .C2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n966), .B1(new_n1158), .B2(new_n1172), .ZN(new_n1173));
  AND2_X1   g748(.A1(new_n989), .A2(new_n992), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1155), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1079), .A2(new_n1100), .A3(new_n1104), .ZN(new_n1176));
  OAI211_X1 g751(.A(new_n1174), .B(new_n995), .C1(new_n1175), .C2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1166), .A2(new_n1163), .ZN(new_n1178));
  AND2_X1   g753(.A1(new_n1169), .A2(new_n980), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1171), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1178), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1177), .A2(new_n1181), .A3(KEYINPUT127), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1173), .A2(new_n1182), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g758(.A1(new_n893), .A2(new_n897), .ZN(new_n1185));
  NOR4_X1   g759(.A1(G229), .A2(G227), .A3(new_n459), .A4(G401), .ZN(new_n1186));
  AND4_X1   g760(.A1(new_n1185), .A2(new_n954), .A3(new_n957), .A4(new_n1186), .ZN(G308));
  NAND4_X1  g761(.A1(new_n1185), .A2(new_n954), .A3(new_n957), .A4(new_n1186), .ZN(G225));
endmodule


