//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 1 1 1 1 1 1 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0 1 1 0 0 1 0 0 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n587,
    new_n588, new_n589, new_n590, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  AND2_X1   g001(.A1(new_n187), .A2(G952), .ZN(new_n188));
  NAND2_X1  g002(.A1(G234), .A2(G237), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT21), .B(G898), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G953), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n189), .A2(G902), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n190), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  XOR2_X1   g008(.A(new_n194), .B(KEYINPUT94), .Z(new_n195));
  OAI21_X1  g009(.A(G214), .B1(G237), .B2(G902), .ZN(new_n196));
  OAI21_X1  g010(.A(G210), .B1(G237), .B2(G902), .ZN(new_n197));
  INV_X1    g011(.A(G104), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT3), .B1(new_n198), .B2(G107), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n200));
  INV_X1    g014(.A(G107), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(G104), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(G107), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n199), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT79), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT79), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n199), .A2(new_n202), .A3(new_n206), .A4(new_n203), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(G101), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT80), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G101), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n199), .A2(new_n202), .A3(new_n211), .A4(new_n203), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n205), .A2(KEYINPUT80), .A3(G101), .A4(new_n207), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n210), .A2(KEYINPUT4), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT81), .ZN(new_n215));
  OR3_X1    g029(.A1(new_n208), .A2(new_n215), .A3(KEYINPUT4), .ZN(new_n216));
  XNOR2_X1  g030(.A(G116), .B(G119), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT2), .B(G113), .ZN(new_n218));
  XNOR2_X1  g032(.A(new_n217), .B(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n215), .B1(new_n208), .B2(KEYINPUT4), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n214), .A2(new_n216), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G113), .ZN(new_n223));
  XOR2_X1   g037(.A(KEYINPUT86), .B(KEYINPUT5), .Z(new_n224));
  INV_X1    g038(.A(G116), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n225), .A2(G119), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n223), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n217), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n227), .B1(new_n228), .B2(new_n224), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n228), .A2(new_n218), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n201), .A2(G104), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n198), .A2(G107), .ZN(new_n233));
  OAI21_X1  g047(.A(G101), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n229), .A2(new_n231), .A3(new_n212), .A4(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n222), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(G110), .B(G122), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n222), .A2(new_n237), .A3(new_n235), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n239), .A2(KEYINPUT6), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT6), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n236), .A2(new_n242), .A3(new_n238), .ZN(new_n243));
  XNOR2_X1  g057(.A(G143), .B(G146), .ZN(new_n244));
  NAND2_X1  g058(.A1(KEYINPUT0), .A2(G128), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XOR2_X1   g060(.A(KEYINPUT0), .B(G128), .Z(new_n247));
  OAI21_X1  g061(.A(new_n246), .B1(new_n244), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G125), .ZN(new_n249));
  INV_X1    g063(.A(G128), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n250), .A2(KEYINPUT1), .ZN(new_n251));
  INV_X1    g065(.A(G146), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G143), .ZN(new_n253));
  INV_X1    g067(.A(G143), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G146), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n251), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n250), .A2(new_n252), .A3(G143), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n254), .B(G146), .C1(new_n250), .C2(KEYINPUT1), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G125), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n249), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n187), .A2(G224), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n262), .B(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n241), .A2(new_n243), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT87), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT87), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n241), .A2(new_n267), .A3(new_n243), .A4(new_n264), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n212), .A2(new_n234), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n229), .A2(new_n231), .A3(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n237), .B(KEYINPUT8), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n217), .A2(KEYINPUT5), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n230), .B1(new_n227), .B2(new_n273), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n271), .B(new_n272), .C1(new_n270), .C2(new_n274), .ZN(new_n275));
  AND4_X1   g089(.A1(KEYINPUT7), .A2(new_n249), .A3(new_n263), .A4(new_n261), .ZN(new_n276));
  AOI22_X1  g090(.A1(new_n249), .A2(new_n261), .B1(KEYINPUT7), .B2(new_n263), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT88), .ZN(new_n279));
  OR2_X1    g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n279), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n281), .A3(new_n240), .ZN(new_n282));
  INV_X1    g096(.A(G902), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n197), .B1(new_n269), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n197), .ZN(new_n287));
  AOI211_X1 g101(.A(new_n287), .B(new_n284), .C1(new_n266), .C2(new_n268), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n195), .B(new_n196), .C1(new_n286), .C2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n291));
  INV_X1    g105(.A(G134), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G137), .ZN(new_n293));
  INV_X1    g107(.A(G137), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G134), .ZN(new_n295));
  AND3_X1   g109(.A1(new_n293), .A2(new_n295), .A3(KEYINPUT64), .ZN(new_n296));
  OAI21_X1  g110(.A(G131), .B1(new_n295), .B2(KEYINPUT64), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT65), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT11), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n299), .B1(new_n292), .B2(G137), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n294), .A2(KEYINPUT11), .A3(G134), .ZN(new_n301));
  INV_X1    g115(.A(G131), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n300), .A2(new_n301), .A3(new_n302), .A4(new_n293), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n292), .A2(G137), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT64), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n302), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT65), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n293), .A2(new_n295), .A3(KEYINPUT64), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n298), .A2(new_n303), .A3(new_n259), .A4(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n300), .A2(new_n293), .A3(new_n301), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G131), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n303), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n248), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n315), .A2(KEYINPUT30), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT30), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n317), .B1(new_n310), .B2(new_n314), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n220), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n310), .A2(new_n314), .A3(new_n219), .ZN(new_n320));
  NOR2_X1   g134(.A1(G237), .A2(G953), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G210), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT67), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n322), .B(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n324), .B(KEYINPUT68), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT26), .B(G101), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n326), .B(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n325), .B(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n319), .A2(new_n320), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(KEYINPUT31), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT31), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n319), .A2(new_n329), .A3(new_n332), .A4(new_n320), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT70), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n315), .A2(KEYINPUT69), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT69), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n310), .A2(new_n314), .A3(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n336), .A2(new_n219), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT28), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n320), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n219), .B1(new_n310), .B2(new_n314), .ZN(new_n343));
  OAI21_X1  g157(.A(KEYINPUT28), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  AOI211_X1 g158(.A(new_n335), .B(new_n329), .C1(new_n341), .C2(new_n344), .ZN(new_n345));
  AND3_X1   g159(.A1(new_n310), .A2(new_n314), .A3(new_n337), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n337), .B1(new_n310), .B2(new_n314), .ZN(new_n347));
  NOR3_X1   g161(.A1(new_n346), .A2(new_n347), .A3(new_n220), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n344), .B1(new_n348), .B2(KEYINPUT28), .ZN(new_n349));
  INV_X1    g163(.A(new_n329), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT70), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NOR3_X1   g165(.A1(new_n334), .A2(new_n345), .A3(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(G472), .A2(G902), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n291), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n315), .A2(new_n220), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n340), .B1(new_n356), .B2(new_n320), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n357), .B1(new_n340), .B2(new_n339), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n335), .B1(new_n358), .B2(new_n329), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n349), .A2(KEYINPUT70), .A3(new_n350), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n359), .A2(new_n331), .A3(new_n333), .A4(new_n360), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n361), .A2(KEYINPUT32), .A3(new_n353), .ZN(new_n362));
  AOI21_X1  g176(.A(KEYINPUT32), .B1(new_n361), .B2(new_n353), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n355), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n361), .A2(new_n353), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(new_n291), .A3(KEYINPUT32), .ZN(new_n366));
  INV_X1    g180(.A(new_n341), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT72), .B1(new_n342), .B2(new_n343), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n368), .B1(KEYINPUT72), .B2(new_n342), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n367), .B1(new_n369), .B2(KEYINPUT28), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n370), .A2(KEYINPUT29), .A3(new_n329), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n283), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n319), .A2(new_n320), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n350), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n349), .A2(new_n329), .ZN(new_n375));
  AOI21_X1  g189(.A(KEYINPUT29), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(G472), .B1(new_n372), .B2(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n364), .A2(new_n366), .A3(new_n377), .ZN(new_n378));
  XOR2_X1   g192(.A(KEYINPUT73), .B(G217), .Z(new_n379));
  INV_X1    g193(.A(G234), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n379), .B1(new_n380), .B2(G902), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT23), .ZN(new_n382));
  INV_X1    g196(.A(G119), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n382), .B1(new_n383), .B2(G128), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(G128), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n250), .A2(KEYINPUT23), .A3(G119), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  OR2_X1    g201(.A1(new_n387), .A2(KEYINPUT75), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(KEYINPUT75), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n389), .A3(G110), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT76), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT16), .ZN(new_n393));
  NOR3_X1   g207(.A1(new_n260), .A2(KEYINPUT77), .A3(G140), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G140), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G125), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n260), .A2(G140), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(new_n398), .A3(KEYINPUT77), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n393), .B1(new_n395), .B2(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n397), .A2(KEYINPUT16), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n252), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n401), .ZN(new_n403));
  XNOR2_X1  g217(.A(G125), .B(G140), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n394), .B1(new_n404), .B2(KEYINPUT77), .ZN(new_n405));
  OAI211_X1 g219(.A(G146), .B(new_n403), .C1(new_n405), .C2(new_n393), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n402), .A2(new_n406), .ZN(new_n407));
  XOR2_X1   g221(.A(KEYINPUT24), .B(G110), .Z(new_n408));
  XNOR2_X1  g222(.A(new_n408), .B(KEYINPUT74), .ZN(new_n409));
  XNOR2_X1  g223(.A(G119), .B(G128), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n388), .A2(new_n389), .A3(KEYINPUT76), .A4(G110), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n392), .A2(new_n407), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(KEYINPUT78), .B(G110), .ZN(new_n414));
  OAI22_X1  g228(.A1(new_n409), .A2(new_n410), .B1(new_n387), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n404), .A2(new_n252), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(new_n406), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(KEYINPUT22), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n420), .B(G137), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n413), .A2(new_n417), .A3(new_n421), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(new_n283), .A3(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT25), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n423), .A2(KEYINPUT25), .A3(new_n283), .A4(new_n424), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n381), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n381), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n425), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(G469), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n270), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n259), .A2(new_n212), .A3(new_n234), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n313), .ZN(new_n439));
  XOR2_X1   g253(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n440));
  NOR3_X1   g254(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n435), .A2(new_n436), .A3(KEYINPUT83), .ZN(new_n442));
  AOI21_X1  g256(.A(KEYINPUT83), .B1(new_n435), .B2(new_n436), .ZN(new_n443));
  NOR3_X1   g257(.A1(new_n442), .A2(new_n443), .A3(new_n439), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT84), .B1(new_n444), .B2(KEYINPUT12), .ZN(new_n445));
  INV_X1    g259(.A(new_n443), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n435), .A2(new_n436), .A3(KEYINPUT83), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(new_n313), .A3(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT84), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT12), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n441), .B1(new_n445), .B2(new_n451), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n214), .A2(new_n216), .A3(new_n248), .A4(new_n221), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n436), .B(KEYINPUT10), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n453), .A2(new_n439), .A3(new_n454), .ZN(new_n455));
  XOR2_X1   g269(.A(G110), .B(G140), .Z(new_n456));
  AND2_X1   g270(.A1(new_n187), .A2(G227), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n456), .B(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n452), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n439), .B1(new_n453), .B2(new_n454), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n458), .B1(new_n462), .B2(new_n455), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n433), .B(new_n283), .C1(new_n460), .C2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT85), .ZN(new_n465));
  INV_X1    g279(.A(new_n455), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n466), .A2(new_n461), .ZN(new_n467));
  OAI22_X1  g281(.A1(new_n467), .A2(new_n458), .B1(new_n452), .B2(new_n459), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT85), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n468), .A2(new_n469), .A3(new_n433), .A4(new_n283), .ZN(new_n470));
  INV_X1    g284(.A(new_n441), .ZN(new_n471));
  NOR3_X1   g285(.A1(new_n444), .A2(KEYINPUT84), .A3(KEYINPUT12), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n449), .B1(new_n448), .B2(new_n450), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n458), .B1(new_n474), .B2(new_n455), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n459), .A2(new_n461), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n283), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AOI22_X1  g291(.A1(new_n465), .A2(new_n470), .B1(G469), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G221), .ZN(new_n479));
  XOR2_X1   g293(.A(KEYINPUT9), .B(G234), .Z(new_n480));
  AOI21_X1  g294(.A(new_n479), .B1(new_n480), .B2(new_n283), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT93), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n321), .A2(G143), .A3(G214), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(G143), .B1(new_n321), .B2(G214), .ZN(new_n485));
  OAI211_X1 g299(.A(KEYINPUT17), .B(G131), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT92), .ZN(new_n487));
  INV_X1    g301(.A(G237), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n488), .A2(new_n187), .A3(G214), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n254), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n483), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT92), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n491), .A2(new_n492), .A3(KEYINPUT17), .A4(G131), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n487), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n482), .B1(new_n494), .B2(new_n407), .ZN(new_n495));
  OR3_X1    g309(.A1(new_n491), .A2(KEYINPUT90), .A3(G131), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT17), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n491), .A2(G131), .ZN(new_n498));
  OAI21_X1  g312(.A(KEYINPUT90), .B1(new_n491), .B2(G131), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n496), .A2(new_n497), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n487), .A2(new_n493), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n501), .A2(KEYINPUT93), .A3(new_n402), .A4(new_n406), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n495), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(G113), .B(G122), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(new_n198), .ZN(new_n505));
  INV_X1    g319(.A(new_n498), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n405), .A2(G146), .ZN(new_n507));
  AOI22_X1  g321(.A1(new_n506), .A2(KEYINPUT18), .B1(new_n507), .B2(new_n416), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT18), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n490), .B(new_n483), .C1(new_n509), .C2(new_n302), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(KEYINPUT89), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n503), .A2(new_n505), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n505), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT19), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n404), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n395), .A2(new_n399), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n516), .B1(new_n517), .B2(new_n515), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n518), .A2(G146), .ZN(new_n519));
  INV_X1    g333(.A(new_n406), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n496), .A2(new_n498), .A3(new_n499), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n512), .ZN(new_n524));
  OAI211_X1 g338(.A(KEYINPUT91), .B(new_n514), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT91), .ZN(new_n526));
  AOI22_X1  g340(.A1(new_n521), .A2(new_n522), .B1(new_n508), .B2(new_n511), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n526), .B1(new_n527), .B2(new_n505), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n513), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(G475), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(new_n530), .A3(new_n283), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT20), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n513), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n505), .B1(new_n503), .B2(new_n512), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n283), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(G475), .ZN(new_n537));
  XNOR2_X1  g351(.A(G128), .B(G143), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(new_n292), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n225), .A2(KEYINPUT14), .A3(G122), .ZN(new_n540));
  XNOR2_X1  g354(.A(G116), .B(G122), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  OAI211_X1 g356(.A(G107), .B(new_n540), .C1(new_n542), .C2(KEYINPUT14), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n539), .B(new_n543), .C1(G107), .C2(new_n542), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n538), .A2(KEYINPUT13), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n254), .A2(G128), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n545), .B(G134), .C1(KEYINPUT13), .C2(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n541), .B(new_n201), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n538), .A2(new_n292), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n544), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n379), .A2(new_n480), .A3(new_n187), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n551), .A2(new_n552), .ZN(new_n554));
  OR2_X1    g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n283), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT15), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(G478), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n556), .B(new_n558), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n529), .A2(KEYINPUT20), .A3(new_n530), .A4(new_n283), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n533), .A2(new_n537), .A3(new_n559), .A4(new_n560), .ZN(new_n561));
  NOR3_X1   g375(.A1(new_n478), .A2(new_n481), .A3(new_n561), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n290), .A2(new_n378), .A3(new_n432), .A4(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(G101), .ZN(G3));
  NAND2_X1  g378(.A1(new_n465), .A2(new_n470), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n477), .A2(G469), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n481), .ZN(new_n568));
  INV_X1    g382(.A(G472), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n569), .B1(new_n361), .B2(new_n283), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n570), .B1(new_n353), .B2(new_n361), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n567), .A2(new_n432), .A3(new_n568), .A4(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n533), .A2(new_n537), .A3(new_n560), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n554), .A2(KEYINPUT96), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n574), .A2(new_n553), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT33), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n576), .B1(new_n554), .B2(KEYINPUT96), .ZN(new_n577));
  XOR2_X1   g391(.A(KEYINPUT95), .B(KEYINPUT33), .Z(new_n578));
  AOI22_X1  g392(.A1(new_n575), .A2(new_n577), .B1(new_n555), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n579), .A2(G478), .A3(new_n283), .ZN(new_n580));
  INV_X1    g394(.A(new_n556), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n580), .B1(G478), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n573), .A2(new_n582), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n572), .A2(new_n289), .A3(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(KEYINPUT34), .B(G104), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n584), .B(new_n585), .ZN(G6));
  NOR2_X1   g400(.A1(new_n573), .A2(new_n559), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n572), .A2(new_n289), .A3(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(KEYINPUT35), .B(G107), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n589), .B(new_n590), .ZN(G9));
  INV_X1    g405(.A(KEYINPUT99), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n430), .A2(G902), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n418), .A2(KEYINPUT97), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT97), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n413), .A2(new_n596), .A3(new_n417), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n598), .B1(KEYINPUT36), .B2(new_n422), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n422), .A2(KEYINPUT36), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n595), .A2(new_n600), .A3(new_n597), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n594), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n429), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT98), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(KEYINPUT98), .B1(new_n602), .B2(new_n429), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(G472), .B1(new_n352), .B2(G902), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n365), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n592), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n606), .A2(new_n607), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n612), .A2(KEYINPUT99), .A3(new_n571), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n290), .A2(new_n562), .A3(new_n611), .A4(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(KEYINPUT100), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT37), .B(G110), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G12));
  AOI21_X1  g431(.A(new_n481), .B1(new_n565), .B2(new_n566), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n378), .A2(new_n618), .ZN(new_n619));
  OR2_X1    g433(.A1(new_n187), .A2(G900), .ZN(new_n620));
  OR3_X1    g434(.A1(new_n620), .A2(new_n193), .A3(KEYINPUT101), .ZN(new_n621));
  OAI21_X1  g435(.A(KEYINPUT101), .B1(new_n620), .B2(new_n193), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n621), .A2(new_n190), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n573), .A2(new_n559), .A3(new_n624), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n625), .B(new_n196), .C1(new_n286), .C2(new_n288), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n619), .A2(KEYINPUT102), .A3(new_n612), .A4(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT102), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n378), .A2(new_n618), .A3(new_n612), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n629), .B1(new_n630), .B2(new_n626), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G128), .ZN(G30));
  NAND2_X1  g447(.A1(new_n269), .A2(new_n285), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n287), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n269), .A2(new_n197), .A3(new_n285), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT103), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT38), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n373), .A2(new_n350), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n283), .B1(new_n369), .B2(new_n329), .ZN(new_n641));
  OAI21_X1  g455(.A(G472), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n364), .A2(new_n366), .A3(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n644), .A2(new_n196), .A3(new_n608), .ZN(new_n645));
  INV_X1    g459(.A(new_n559), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n573), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n623), .B(KEYINPUT39), .Z(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n618), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT40), .ZN(new_n652));
  NOR4_X1   g466(.A1(new_n639), .A2(new_n645), .A3(new_n648), .A4(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(new_n254), .ZN(G45));
  INV_X1    g468(.A(new_n196), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n655), .B1(new_n635), .B2(new_n636), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT104), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n573), .A2(new_n582), .A3(new_n623), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n656), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n196), .B1(new_n286), .B2(new_n288), .ZN(new_n661));
  OAI21_X1  g475(.A(KEYINPUT104), .B1(new_n661), .B2(new_n658), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n630), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(new_n252), .ZN(G48));
  INV_X1    g478(.A(new_n583), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n290), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n468), .A2(new_n283), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(G469), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n565), .A2(new_n568), .A3(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n670), .A2(new_n378), .A3(new_n432), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n666), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT41), .B(G113), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G15));
  NOR3_X1   g488(.A1(new_n671), .A2(new_n289), .A3(new_n588), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(new_n225), .ZN(G18));
  NAND3_X1  g490(.A1(new_n656), .A2(new_n195), .A3(new_n670), .ZN(new_n677));
  INV_X1    g491(.A(new_n561), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n378), .A2(new_n678), .A3(new_n612), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(new_n383), .ZN(G21));
  NAND4_X1  g495(.A1(new_n637), .A2(KEYINPUT105), .A3(new_n196), .A4(new_n647), .ZN(new_n682));
  OAI211_X1 g496(.A(new_n647), .B(new_n196), .C1(new_n286), .C2(new_n288), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT105), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  OAI211_X1 g500(.A(new_n331), .B(new_n333), .C1(new_n370), .C2(new_n329), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n570), .B1(new_n353), .B2(new_n687), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n688), .A2(new_n432), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n686), .A2(new_n195), .A3(new_n670), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G122), .ZN(G24));
  AND2_X1   g505(.A1(new_n612), .A2(new_n688), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n692), .A2(new_n659), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n693), .A2(new_n656), .A3(new_n670), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G125), .ZN(G27));
  INV_X1    g509(.A(KEYINPUT107), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n618), .A2(KEYINPUT106), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT106), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n698), .B1(new_n478), .B2(new_n481), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n286), .A2(new_n288), .A3(new_n655), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n697), .A2(new_n699), .A3(new_n700), .A4(new_n659), .ZN(new_n701));
  INV_X1    g515(.A(new_n363), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n361), .A2(KEYINPUT32), .A3(new_n353), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n377), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n704), .A2(KEYINPUT42), .A3(new_n432), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n696), .B1(new_n701), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n618), .A2(KEYINPUT106), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n478), .A2(new_n698), .A3(new_n481), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n635), .A2(new_n196), .A3(new_n636), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n711), .A2(new_n658), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n710), .A2(KEYINPUT107), .A3(new_n712), .A4(new_n705), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n710), .A2(new_n378), .A3(new_n432), .A4(new_n712), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT42), .ZN(new_n715));
  AOI22_X1  g529(.A1(new_n707), .A2(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(new_n302), .ZN(G33));
  NAND2_X1  g531(.A1(new_n378), .A2(new_n432), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(new_n711), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n710), .A3(new_n625), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(KEYINPUT108), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(new_n292), .ZN(G36));
  NOR2_X1   g536(.A1(new_n475), .A2(new_n476), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(G469), .ZN(new_n726));
  NAND2_X1  g540(.A1(G469), .A2(G902), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT46), .ZN(new_n729));
  AOI22_X1  g543(.A1(new_n728), .A2(new_n729), .B1(new_n470), .B2(new_n465), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n726), .A2(KEYINPUT46), .A3(new_n727), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n481), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n732), .A2(new_n650), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT43), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n734), .B1(new_n573), .B2(KEYINPUT109), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n582), .A2(new_n537), .A3(new_n533), .A4(new_n560), .ZN(new_n736));
  XOR2_X1   g550(.A(new_n735), .B(new_n736), .Z(new_n737));
  NAND3_X1  g551(.A1(new_n737), .A2(new_n610), .A3(new_n612), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT44), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n711), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n733), .B(new_n740), .C1(new_n739), .C2(new_n738), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G137), .ZN(G39));
  XNOR2_X1  g556(.A(new_n732), .B(KEYINPUT47), .ZN(new_n743));
  NOR4_X1   g557(.A1(new_n711), .A2(new_n378), .A3(new_n432), .A4(new_n658), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(KEYINPUT110), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G140), .ZN(G42));
  NAND2_X1  g561(.A1(new_n565), .A2(new_n668), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n748), .A2(new_n568), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n700), .B1(new_n743), .B2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n190), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n737), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n689), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n711), .A2(new_n669), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n754), .B1(new_n692), .B2(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n755), .A2(new_n432), .A3(new_n751), .A4(new_n643), .ZN(new_n758));
  OR3_X1    g572(.A1(new_n758), .A2(new_n573), .A3(new_n582), .ZN(new_n759));
  INV_X1    g573(.A(new_n753), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n760), .A2(new_n639), .A3(new_n655), .A4(new_n670), .ZN(new_n761));
  XOR2_X1   g575(.A(new_n761), .B(KEYINPUT50), .Z(new_n762));
  NAND3_X1  g576(.A1(new_n757), .A2(new_n759), .A3(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n757), .A2(KEYINPUT51), .A3(new_n759), .A4(new_n762), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n704), .A2(new_n432), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n756), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(KEYINPUT48), .ZN(new_n769));
  AND4_X1   g583(.A1(new_n188), .A2(new_n765), .A3(new_n766), .A4(new_n769), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n758), .A2(new_n583), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT117), .ZN(new_n772));
  INV_X1    g586(.A(new_n663), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n603), .A2(new_n604), .ZN(new_n774));
  NOR4_X1   g588(.A1(new_n478), .A2(new_n481), .A3(new_n774), .A4(new_n624), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n643), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n618), .A2(new_n604), .A3(new_n603), .A4(new_n623), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(KEYINPUT114), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n686), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n632), .A2(new_n773), .A3(new_n780), .A4(new_n694), .ZN(new_n781));
  XOR2_X1   g595(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n663), .B1(new_n631), .B2(new_n628), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n785), .A2(KEYINPUT52), .A3(new_n694), .A4(new_n780), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n656), .A2(KEYINPUT112), .A3(new_n195), .A4(new_n587), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT112), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n789), .B1(new_n289), .B2(new_n588), .ZN(new_n790));
  INV_X1    g604(.A(new_n432), .ZN(new_n791));
  NOR4_X1   g605(.A1(new_n478), .A2(new_n610), .A3(new_n791), .A4(new_n481), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n788), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n793), .A2(new_n614), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n792), .A2(new_n290), .A3(new_n665), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT111), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n563), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n796), .B1(new_n563), .B2(new_n795), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n794), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI22_X1  g614(.A1(new_n666), .A2(new_n671), .B1(new_n677), .B2(new_n679), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n801), .A2(new_n675), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n690), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n720), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n693), .A2(new_n710), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n561), .A2(new_n624), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(KEYINPUT113), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n619), .A2(new_n612), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n711), .B1(new_n806), .B2(new_n809), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n716), .A2(new_n805), .A3(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n787), .A2(new_n804), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(KEYINPUT53), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n707), .A2(new_n713), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n714), .A2(new_n715), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n810), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n816), .A2(new_n720), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n567), .A2(new_n568), .A3(new_n678), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n718), .A2(new_n289), .A3(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(KEYINPUT111), .B1(new_n820), .B2(new_n584), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(new_n797), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n822), .A2(new_n690), .A3(new_n794), .A4(new_n802), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n818), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT52), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n781), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(new_n786), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n824), .A2(new_n825), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n813), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AOI211_X1 g646(.A(KEYINPUT116), .B(KEYINPUT53), .C1(new_n824), .C2(new_n787), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n834), .B1(new_n812), .B2(new_n825), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n824), .A2(KEYINPUT53), .A3(new_n828), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n833), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n772), .B(new_n832), .C1(new_n838), .C2(new_n831), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n833), .A2(new_n835), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n831), .B1(new_n840), .B2(new_n836), .ZN(new_n841));
  INV_X1    g655(.A(new_n832), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT117), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n770), .A2(new_n771), .A3(new_n839), .A4(new_n843), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n753), .A2(new_n661), .A3(new_n669), .ZN(new_n845));
  OAI22_X1  g659(.A1(new_n844), .A2(new_n845), .B1(G952), .B2(G953), .ZN(new_n846));
  XOR2_X1   g660(.A(new_n748), .B(KEYINPUT49), .Z(new_n847));
  NOR4_X1   g661(.A1(new_n644), .A2(new_n655), .A3(new_n481), .A4(new_n736), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n639), .A2(new_n432), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n846), .A2(new_n849), .ZN(G75));
  NOR2_X1   g664(.A1(new_n830), .A2(new_n283), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT56), .B1(new_n851), .B2(G210), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n241), .A2(new_n243), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(new_n264), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(KEYINPUT55), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n852), .B(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n187), .A2(G952), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n856), .A2(new_n857), .ZN(G51));
  INV_X1    g672(.A(new_n830), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(KEYINPUT54), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n832), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n727), .A2(KEYINPUT57), .ZN(new_n862));
  OR2_X1    g676(.A1(new_n727), .A2(KEYINPUT57), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(new_n468), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n851), .A2(G469), .A3(new_n725), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n857), .B1(new_n865), .B2(new_n866), .ZN(G54));
  NAND3_X1  g681(.A1(new_n851), .A2(KEYINPUT58), .A3(G475), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n868), .B(new_n529), .Z(new_n869));
  NOR2_X1   g683(.A1(new_n869), .A2(new_n857), .ZN(G60));
  XNOR2_X1  g684(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n871));
  NAND2_X1  g685(.A1(G478), .A2(G902), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n871), .B(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n873), .B1(new_n860), .B2(new_n832), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n857), .B1(new_n874), .B2(new_n579), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n873), .B1(new_n843), .B2(new_n839), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n875), .B1(new_n876), .B2(new_n579), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT119), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT119), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n879), .B(new_n875), .C1(new_n876), .C2(new_n579), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n878), .A2(new_n880), .ZN(G63));
  XOR2_X1   g695(.A(KEYINPUT120), .B(KEYINPUT60), .Z(new_n882));
  NAND2_X1  g696(.A1(G217), .A2(G902), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n882), .B(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n859), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n423), .A2(new_n424), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n857), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n599), .A2(new_n601), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n887), .B1(new_n888), .B2(new_n885), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n889), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g704(.A(new_n192), .B1(G224), .B2(new_n187), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT121), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n892), .B1(new_n804), .B2(G953), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n853), .B1(G898), .B2(new_n187), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n893), .B(new_n894), .ZN(G69));
  AND2_X1   g709(.A1(new_n746), .A2(new_n741), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n733), .A2(new_n686), .A3(new_n767), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n785), .A2(new_n694), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n898), .A2(new_n716), .A3(new_n805), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n896), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT125), .Z(new_n901));
  OAI21_X1  g715(.A(new_n620), .B1(new_n901), .B2(G953), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n316), .A2(new_n318), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(new_n518), .Z(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n653), .A2(new_n898), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT122), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT62), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n907), .B(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n908), .A2(new_n909), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n665), .A2(new_n587), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n651), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n915), .B(new_n719), .C1(new_n913), .C2(new_n914), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n911), .A2(new_n912), .A3(new_n896), .A4(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n187), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n904), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n906), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n187), .B1(G227), .B2(G900), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT124), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n920), .B(new_n922), .ZN(G72));
  NAND2_X1  g737(.A1(new_n901), .A2(new_n804), .ZN(new_n924));
  XNOR2_X1  g738(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n569), .A2(new_n283), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n374), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n927), .B1(new_n917), .B2(new_n823), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n929), .A2(new_n640), .ZN(new_n930));
  INV_X1    g744(.A(new_n640), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n931), .A2(new_n374), .A3(new_n927), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT127), .Z(new_n933));
  NOR2_X1   g747(.A1(new_n838), .A2(new_n933), .ZN(new_n934));
  NOR4_X1   g748(.A1(new_n928), .A2(new_n930), .A3(new_n857), .A4(new_n934), .ZN(G57));
endmodule


