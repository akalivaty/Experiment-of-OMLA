//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 1 1 1 1 1 1 0 1 0 1 0 1 1 1 0 0 0 1 1 0 0 0 1 1 0 0 0 0 0 1 1 1 1 0 1 0 1 0 0 1 1 1 0 1 0 1 0 0 1 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:07 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n554, new_n556, new_n557, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n603, new_n605,
    new_n606, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1187;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT65), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT67), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND4_X1  g039(.A1(new_n461), .A2(new_n463), .A3(G137), .A4(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G101), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n461), .A2(new_n463), .A3(G125), .ZN(new_n469));
  OR2_X1    g044(.A1(new_n469), .A2(KEYINPUT68), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n469), .A2(KEYINPUT68), .B1(G113), .B2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n468), .B1(new_n472), .B2(G2105), .ZN(G160));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n474));
  AND3_X1   g049(.A1(new_n461), .A2(new_n463), .A3(new_n464), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G136), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n475), .A2(KEYINPUT69), .A3(G136), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n478), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  AND3_X1   g057(.A1(new_n461), .A2(new_n463), .A3(G2105), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT70), .ZN(new_n484));
  OR2_X1    g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n483), .A2(new_n484), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n482), .B1(G124), .B2(new_n487), .ZN(G162));
  NAND4_X1  g063(.A1(new_n461), .A2(new_n463), .A3(G138), .A4(new_n464), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT71), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n475), .A2(KEYINPUT72), .A3(new_n493), .A4(G138), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT72), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n495), .B1(new_n489), .B2(KEYINPUT4), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n489), .A2(KEYINPUT71), .A3(KEYINPUT4), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n492), .A2(new_n494), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n483), .A2(G126), .ZN(new_n499));
  OR2_X1    g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n500), .B(G2104), .C1(G114), .C2(new_n464), .ZN(new_n501));
  AND2_X1   g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT6), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G651), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n506), .A2(new_n508), .A3(new_n510), .A4(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n510), .A2(new_n512), .A3(G62), .ZN(new_n515));
  NAND2_X1  g090(.A1(G75), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n514), .A2(G88), .B1(new_n517), .B2(G651), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n506), .A2(new_n508), .A3(G50), .A4(G543), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT73), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT6), .B(G651), .ZN(new_n522));
  NAND4_X1  g097(.A1(new_n522), .A2(KEYINPUT73), .A3(G50), .A4(G543), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n518), .A2(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  NAND2_X1  g101(.A1(new_n522), .A2(G543), .ZN(new_n527));
  INV_X1    g102(.A(G51), .ZN(new_n528));
  INV_X1    g103(.A(G89), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n527), .A2(new_n528), .B1(new_n513), .B2(new_n529), .ZN(new_n530));
  XNOR2_X1  g105(.A(KEYINPUT5), .B(G543), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n531), .A2(G63), .A3(G651), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT7), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(new_n534), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n532), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n530), .A2(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  AOI22_X1  g114(.A1(new_n531), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n505), .ZN(new_n541));
  XOR2_X1   g116(.A(KEYINPUT74), .B(G52), .Z(new_n542));
  XOR2_X1   g117(.A(KEYINPUT75), .B(G90), .Z(new_n543));
  OAI22_X1  g118(.A1(new_n527), .A2(new_n542), .B1(new_n513), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n541), .A2(new_n544), .ZN(G171));
  AOI22_X1  g120(.A1(new_n531), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n546), .A2(new_n505), .ZN(new_n547));
  INV_X1    g122(.A(G43), .ZN(new_n548));
  INV_X1    g123(.A(G81), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n527), .A2(new_n548), .B1(new_n513), .B2(new_n549), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  AND3_X1   g128(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G36), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n554), .A2(new_n557), .ZN(G188));
  INV_X1    g133(.A(new_n527), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G53), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT9), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(new_n531), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n565), .A2(G651), .B1(G91), .B2(new_n514), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n561), .A2(new_n566), .ZN(G299));
  INV_X1    g142(.A(G171), .ZN(G301));
  OAI21_X1  g143(.A(G651), .B1(new_n531), .B2(G74), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n522), .A2(new_n531), .A3(G87), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n522), .A2(G49), .A3(G543), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(G288));
  NAND3_X1  g147(.A1(new_n522), .A2(new_n531), .A3(G86), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n506), .A2(new_n508), .A3(G48), .A4(G543), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n510), .A2(new_n512), .A3(G61), .ZN(new_n575));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  AND2_X1   g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g152(.A(new_n573), .B(new_n574), .C1(new_n577), .C2(new_n505), .ZN(G305));
  NAND2_X1  g153(.A1(new_n559), .A2(G47), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n514), .A2(G85), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n531), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n579), .B(new_n580), .C1(new_n505), .C2(new_n581), .ZN(G290));
  NAND2_X1  g157(.A1(G301), .A2(G868), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n514), .A2(G92), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT10), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n584), .B(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(G79), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G66), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n563), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(G651), .B1(new_n559), .B2(G54), .ZN(new_n590));
  AND2_X1   g165(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n583), .B1(new_n591), .B2(G868), .ZN(G284));
  OAI21_X1  g167(.A(new_n583), .B1(new_n591), .B2(G868), .ZN(G321));
  INV_X1    g168(.A(KEYINPUT9), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n560), .B(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n566), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n597), .A2(G868), .ZN(new_n598));
  AND2_X1   g173(.A1(G286), .A2(G868), .ZN(new_n599));
  OAI21_X1  g174(.A(KEYINPUT76), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(KEYINPUT76), .B2(new_n599), .ZN(G297));
  XOR2_X1   g176(.A(G297), .B(KEYINPUT77), .Z(G280));
  INV_X1    g177(.A(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n591), .B1(new_n603), .B2(G860), .ZN(G148));
  NAND2_X1  g179(.A1(new_n591), .A2(new_n603), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(G868), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G868), .B2(new_n552), .ZN(G323));
  XNOR2_X1  g182(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g183(.A1(new_n487), .A2(G123), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n475), .A2(G135), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT79), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n464), .A2(G111), .ZN(new_n613));
  OAI21_X1  g188(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n614));
  OAI211_X1 g189(.A(new_n609), .B(new_n612), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(G2096), .Z(new_n616));
  AND2_X1   g191(.A1(new_n461), .A2(new_n463), .ZN(new_n617));
  INV_X1    g192(.A(new_n467), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT78), .ZN(new_n622));
  INV_X1    g197(.A(G2100), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OR3_X1    g199(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n622), .A2(new_n623), .ZN(new_n626));
  NAND4_X1  g201(.A1(new_n616), .A2(new_n624), .A3(new_n625), .A4(new_n626), .ZN(G156));
  XNOR2_X1  g202(.A(G2427), .B(G2430), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT80), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2435), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n632), .A2(KEYINPUT14), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(KEYINPUT81), .B(KEYINPUT82), .Z(new_n637));
  XOR2_X1   g212(.A(new_n636), .B(new_n637), .Z(new_n638));
  XOR2_X1   g213(.A(G2451), .B(G2454), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n640), .B(new_n641), .Z(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n636), .B(new_n637), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(new_n642), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n644), .A2(G14), .A3(new_n646), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n647), .A2(KEYINPUT83), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(KEYINPUT83), .ZN(new_n649));
  AND2_X1   g224(.A1(new_n648), .A2(new_n649), .ZN(G401));
  XNOR2_X1  g225(.A(G2084), .B(G2090), .ZN(new_n651));
  INV_X1    g226(.A(KEYINPUT84), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2067), .B(G2678), .Z(new_n654));
  XOR2_X1   g229(.A(G2072), .B(G2078), .Z(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT18), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n655), .B(KEYINPUT17), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n659), .A2(new_n653), .A3(new_n654), .ZN(new_n660));
  AND2_X1   g235(.A1(new_n654), .A2(new_n655), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n653), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n662), .A2(KEYINPUT85), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(KEYINPUT85), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n664), .B1(new_n654), .B2(new_n659), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n658), .B(new_n660), .C1(new_n663), .C2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2100), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT86), .B(G2096), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(G227));
  XNOR2_X1  g244(.A(G1971), .B(G1976), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  OR2_X1    g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n673), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n671), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n671), .A2(new_n676), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT20), .ZN(new_n679));
  OAI211_X1 g254(.A(new_n675), .B(new_n677), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(new_n679), .B2(new_n678), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(G1991), .ZN(new_n682));
  INV_X1    g257(.A(G1996), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1981), .B(G1986), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n685), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n684), .B(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n687), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n688), .A2(new_n692), .ZN(G229));
  NAND2_X1  g268(.A1(new_n475), .A2(G131), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n464), .A2(G107), .ZN(new_n695));
  OAI21_X1  g270(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n694), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(new_n487), .B2(G119), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(KEYINPUT87), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT87), .ZN(new_n700));
  INV_X1    g275(.A(G119), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(new_n485), .B2(new_n486), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n700), .B1(new_n702), .B2(new_n697), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G29), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT35), .B(G1991), .ZN(new_n706));
  INV_X1    g281(.A(G29), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G25), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n705), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n706), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n707), .B1(new_n699), .B2(new_n703), .ZN(new_n711));
  INV_X1    g286(.A(new_n708), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  MUX2_X1   g289(.A(G24), .B(G290), .S(G16), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G1986), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT34), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT88), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT32), .B(G1981), .Z(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G86), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n574), .B1(new_n513), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n505), .B1(new_n575), .B2(new_n576), .ZN(new_n725));
  OAI21_X1  g300(.A(G16), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT89), .ZN(new_n727));
  INV_X1    g302(.A(G16), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G6), .ZN(new_n729));
  AND3_X1   g304(.A1(new_n726), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n727), .B1(new_n726), .B2(new_n729), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n722), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n726), .A2(new_n729), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(KEYINPUT89), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n726), .A2(new_n727), .A3(new_n729), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n734), .A2(new_n721), .A3(new_n735), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n728), .B1(new_n518), .B2(new_n524), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n728), .A2(G22), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT90), .Z(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(G1971), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n517), .A2(G651), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n522), .A2(new_n531), .A3(G88), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n521), .A2(new_n523), .ZN(new_n746));
  OAI21_X1  g321(.A(G16), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(G1971), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n747), .A2(new_n748), .A3(new_n740), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n569), .A2(new_n570), .A3(new_n571), .A4(G16), .ZN(new_n750));
  OR2_X1    g325(.A1(G16), .A2(G23), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT33), .B(G1976), .Z(new_n752));
  AND3_X1   g327(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n752), .B1(new_n750), .B2(new_n751), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AND3_X1   g330(.A1(new_n742), .A2(new_n749), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n720), .B1(new_n737), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n732), .A2(new_n736), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n742), .A2(new_n749), .A3(new_n755), .ZN(new_n759));
  NOR3_X1   g334(.A1(new_n758), .A2(KEYINPUT88), .A3(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n719), .B1(new_n757), .B2(new_n760), .ZN(new_n761));
  NAND4_X1  g336(.A1(new_n756), .A2(new_n720), .A3(new_n736), .A4(new_n732), .ZN(new_n762));
  OAI21_X1  g337(.A(KEYINPUT88), .B1(new_n758), .B2(new_n759), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n762), .A2(new_n763), .A3(KEYINPUT34), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n718), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT91), .ZN(new_n766));
  OAI21_X1  g341(.A(KEYINPUT36), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n716), .B1(new_n709), .B2(new_n713), .ZN(new_n768));
  AND3_X1   g343(.A1(new_n762), .A2(new_n763), .A3(KEYINPUT34), .ZN(new_n769));
  AOI21_X1  g344(.A(KEYINPUT34), .B1(new_n762), .B2(new_n763), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n771), .A2(KEYINPUT91), .ZN(new_n772));
  OAI21_X1  g347(.A(KEYINPUT92), .B1(new_n767), .B2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT36), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n771), .B2(KEYINPUT91), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT92), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n765), .A2(new_n766), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n774), .B(new_n768), .C1(new_n769), .C2(new_n770), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT93), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n773), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n728), .A2(G19), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n552), .B2(new_n728), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1341), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n728), .A2(G21), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G168), .B2(new_n728), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(G1966), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT31), .B(G11), .Z(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT97), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT30), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n790), .A2(G28), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n707), .B1(new_n790), .B2(G28), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n787), .B(new_n789), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n784), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(G171), .A2(G16), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G5), .B2(G16), .ZN(new_n796));
  INV_X1    g371(.A(G1961), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT98), .ZN(new_n799));
  NOR2_X1   g374(.A1(G29), .A2(G32), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n475), .A2(G141), .ZN(new_n801));
  NAND3_X1  g376(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT26), .Z(new_n803));
  NAND2_X1  g378(.A1(new_n618), .A2(G105), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n801), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n487), .B2(G129), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n800), .B1(new_n806), .B2(G29), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT27), .B(G1996), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  OAI22_X1  g384(.A1(new_n786), .A2(G1966), .B1(new_n615), .B2(new_n707), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(new_n797), .B2(new_n796), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n794), .A2(new_n799), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n728), .A2(G4), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n586), .A2(new_n590), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n813), .B1(new_n814), .B2(G16), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G1348), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT24), .ZN(new_n817));
  INV_X1    g392(.A(G34), .ZN(new_n818));
  AOI21_X1  g393(.A(G29), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(new_n817), .B2(new_n818), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G160), .B2(new_n707), .ZN(new_n821));
  INV_X1    g396(.A(G2084), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n617), .A2(G127), .ZN(new_n824));
  NAND2_X1  g399(.A1(G115), .A2(G2104), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(G2105), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n475), .A2(G139), .ZN(new_n828));
  INV_X1    g403(.A(G103), .ZN(new_n829));
  OAI21_X1  g404(.A(KEYINPUT25), .B1(new_n467), .B2(new_n829), .ZN(new_n830));
  OR3_X1    g405(.A1(new_n467), .A2(KEYINPUT25), .A3(new_n829), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n827), .A2(new_n828), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(G29), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n707), .A2(G33), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(KEYINPUT95), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT95), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n833), .A2(new_n837), .A3(new_n834), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(G2072), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n816), .B(new_n823), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n812), .A2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(G2090), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n707), .A2(G35), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(G162), .B2(new_n707), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n845), .A2(KEYINPUT29), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(KEYINPUT29), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n843), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT99), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n846), .A2(new_n843), .A3(new_n847), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n707), .A2(G27), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(G164), .B2(new_n707), .ZN(new_n852));
  INV_X1    g427(.A(G2078), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(G2067), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT28), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n475), .A2(G140), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT94), .ZN(new_n859));
  NOR3_X1   g434(.A1(new_n859), .A2(G104), .A3(G2105), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n859), .B1(G104), .B2(G2105), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n861), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n858), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n863), .B1(new_n487), .B2(G128), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n864), .A2(new_n707), .ZN(new_n865));
  INV_X1    g440(.A(G26), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n866), .A2(G29), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n857), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n867), .A2(KEYINPUT28), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n856), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OR3_X1    g446(.A1(new_n869), .A2(new_n856), .A3(new_n870), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n855), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n839), .A2(new_n840), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(KEYINPUT96), .ZN(new_n875));
  INV_X1    g450(.A(G1956), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n728), .A2(G20), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(KEYINPUT23), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT23), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n879), .B1(G299), .B2(G16), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n876), .B(new_n878), .C1(new_n880), .C2(new_n877), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT96), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n839), .A2(new_n882), .A3(new_n840), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n878), .B1(new_n880), .B2(new_n877), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(G1956), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n875), .A2(new_n881), .A3(new_n883), .A4(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n842), .A2(new_n849), .A3(new_n873), .A4(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT100), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR3_X1   g465(.A1(new_n886), .A2(new_n812), .A3(new_n841), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n891), .A2(KEYINPUT100), .A3(new_n873), .A4(new_n849), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n781), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(G311));
  NAND2_X1  g470(.A1(new_n894), .A2(KEYINPUT101), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT101), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n781), .A2(new_n893), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(G150));
  XNOR2_X1  g474(.A(KEYINPUT103), .B(G55), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n559), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n514), .A2(G93), .ZN(new_n902));
  AOI22_X1  g477(.A1(new_n531), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n903));
  OAI211_X1 g478(.A(new_n901), .B(new_n902), .C1(new_n505), .C2(new_n903), .ZN(new_n904));
  XOR2_X1   g479(.A(KEYINPUT104), .B(G860), .Z(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XOR2_X1   g481(.A(new_n906), .B(KEYINPUT37), .Z(new_n907));
  NAND2_X1  g482(.A1(new_n591), .A2(G559), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT39), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT102), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(KEYINPUT38), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n551), .B(new_n904), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n905), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n915), .B1(new_n911), .B2(new_n913), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n907), .B1(new_n914), .B2(new_n916), .ZN(G145));
  XNOR2_X1  g492(.A(new_n615), .B(new_n864), .ZN(new_n918));
  XNOR2_X1  g493(.A(G162), .B(G160), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n918), .B(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n620), .B(KEYINPUT107), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(new_n832), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n704), .B(new_n503), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n487), .A2(G130), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n475), .A2(G142), .ZN(new_n927));
  OAI21_X1  g502(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT106), .ZN(new_n929));
  OR2_X1    g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n931));
  OR3_X1    g506(.A1(new_n931), .A2(new_n464), .A3(G118), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n928), .A2(new_n929), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n931), .B1(new_n464), .B2(G118), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n930), .A2(new_n932), .A3(new_n933), .A4(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n926), .A2(new_n927), .A3(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n936), .B(new_n806), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n925), .B(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n920), .A2(new_n922), .ZN(new_n939));
  OR3_X1    g514(.A1(new_n924), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(G37), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n938), .B1(new_n924), .B2(new_n939), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  XOR2_X1   g518(.A(KEYINPUT108), .B(KEYINPUT40), .Z(new_n944));
  XNOR2_X1  g519(.A(new_n943), .B(new_n944), .ZN(G395));
  XNOR2_X1  g520(.A(new_n605), .B(new_n912), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n591), .A2(G299), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n597), .A2(new_n814), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT41), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT109), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n948), .A2(new_n949), .A3(KEYINPUT41), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n950), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n956), .A2(KEYINPUT109), .A3(KEYINPUT41), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n947), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n959));
  OR2_X1    g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G288), .ZN(new_n961));
  XNOR2_X1  g536(.A(G290), .B(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(G303), .B(G305), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n962), .B(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT111), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n965), .B(KEYINPUT42), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n958), .A2(new_n959), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n946), .A2(new_n950), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n960), .A2(new_n966), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT112), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n967), .A2(new_n968), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n972), .A2(KEYINPUT112), .A3(new_n966), .A4(new_n960), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n960), .A2(new_n967), .A3(new_n968), .ZN(new_n974));
  INV_X1    g549(.A(new_n966), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n971), .A2(new_n973), .A3(new_n976), .ZN(new_n977));
  MUX2_X1   g552(.A(new_n904), .B(new_n977), .S(G868), .Z(G295));
  MUX2_X1   g553(.A(new_n904), .B(new_n977), .S(G868), .Z(G331));
  XNOR2_X1  g554(.A(G286), .B(G171), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n913), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n980), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n982), .A2(new_n912), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n956), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n981), .A2(KEYINPUT113), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT113), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n986), .B1(new_n913), .B2(new_n980), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n983), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT114), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n990), .B1(new_n950), .B2(new_n951), .ZN(new_n991));
  AOI22_X1  g566(.A1(new_n988), .A2(new_n989), .B1(new_n954), .B2(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n991), .A2(new_n954), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n984), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n964), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT115), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n955), .B(new_n957), .C1(new_n983), .C2(new_n981), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n988), .A2(new_n950), .A3(new_n989), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n998), .A2(new_n999), .A3(new_n996), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n941), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT115), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n991), .A2(new_n954), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n983), .B1(new_n985), .B2(new_n987), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n1004), .A2(new_n1005), .A3(new_n993), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1003), .B(new_n964), .C1(new_n1006), .C2(new_n984), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n997), .A2(new_n1002), .A3(new_n1007), .A4(KEYINPUT43), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT43), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n996), .B1(new_n998), .B2(new_n999), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1009), .B1(new_n1001), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT44), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n997), .A2(new_n1002), .A3(new_n1007), .A4(new_n1009), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT43), .B1(new_n1001), .B2(new_n1010), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT44), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1013), .A2(new_n1018), .ZN(G397));
  INV_X1    g594(.A(G1384), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n503), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT45), .ZN(new_n1022));
  INV_X1    g597(.A(G40), .ZN(new_n1023));
  AOI211_X1 g598(.A(new_n1023), .B(new_n468), .C1(new_n472), .C2(G2105), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1021), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g601(.A(new_n806), .B(G1996), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n864), .B(G2067), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n704), .A2(new_n706), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n699), .A2(new_n710), .A3(new_n703), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g607(.A(G290), .B(G1986), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1026), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(G1384), .B1(new_n498), .B2(new_n502), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT50), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1024), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AOI211_X1 g612(.A(KEYINPUT50), .B(G1384), .C1(new_n498), .C2(new_n502), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n876), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1035), .A2(KEYINPUT45), .ZN(new_n1041));
  XNOR2_X1  g616(.A(KEYINPUT56), .B(G2072), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1040), .A2(new_n1041), .A3(new_n1024), .A4(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT119), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT57), .B1(new_n566), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(G299), .A2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n561), .B(new_n566), .C1(new_n1044), .C2(KEYINPUT57), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1039), .A2(new_n1043), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1035), .A2(new_n1024), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1050), .A2(G2067), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1021), .A2(KEYINPUT50), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1052), .A2(new_n1024), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G1348), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1051), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n1049), .A2(new_n814), .A3(new_n1056), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1039), .A2(new_n1043), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT120), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1048), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1058), .A2(KEYINPUT120), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1057), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT60), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1065), .A2(G1348), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1064), .B1(new_n1066), .B2(new_n1051), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1056), .A2(KEYINPUT60), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1067), .A2(new_n1068), .A3(new_n591), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1056), .A2(KEYINPUT60), .A3(new_n814), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1048), .B1(new_n1039), .B2(new_n1043), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1049), .A2(new_n1071), .A3(KEYINPUT61), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n1058), .A2(KEYINPUT61), .A3(new_n1048), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1069), .B(new_n1070), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n552), .A2(KEYINPUT122), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1040), .A2(new_n683), .A3(new_n1041), .A4(new_n1024), .ZN(new_n1076));
  XOR2_X1   g651(.A(KEYINPUT58), .B(G1341), .Z(new_n1077));
  NAND2_X1  g652(.A1(new_n1050), .A2(new_n1077), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n1076), .A2(KEYINPUT121), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT121), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1075), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  OAI211_X1 g658(.A(KEYINPUT59), .B(new_n1075), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1063), .B1(new_n1074), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G8), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1024), .B1(new_n1035), .B2(KEYINPUT45), .ZN(new_n1088));
  AOI211_X1 g663(.A(new_n1022), .B(G1384), .C1(new_n498), .C2(new_n502), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n748), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1052), .A2(new_n843), .A3(new_n1024), .A4(new_n1053), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1087), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(G303), .A2(G8), .ZN(new_n1093));
  XOR2_X1   g668(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n1094));
  XNOR2_X1  g669(.A(new_n1093), .B(new_n1094), .ZN(new_n1095));
  OR2_X1    g670(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1097), .A2(KEYINPUT53), .A3(new_n853), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1040), .A2(new_n853), .A3(new_n1041), .A4(new_n1024), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1054), .A2(new_n797), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1098), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(G171), .A2(KEYINPUT125), .A3(KEYINPUT54), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(KEYINPUT54), .B2(G171), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n961), .A2(G1976), .ZN(new_n1108));
  INV_X1    g683(.A(G1976), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT52), .B1(G288), .B2(new_n1109), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1050), .A2(G8), .A3(new_n1108), .A4(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(G305), .A2(G1981), .ZN(new_n1112));
  OR3_X1    g687(.A1(new_n724), .A2(new_n725), .A3(G1981), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT49), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1112), .A2(new_n1113), .A3(KEYINPUT49), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1116), .A2(new_n1050), .A3(G8), .A4(new_n1117), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1050), .A2(G8), .A3(new_n1108), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT52), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1111), .B(new_n1118), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1121), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1098), .A2(new_n1101), .A3(new_n1102), .A4(new_n1105), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1096), .A2(new_n1107), .A3(new_n1122), .A4(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(G1966), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1052), .A2(new_n822), .A3(new_n1024), .A4(new_n1053), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1087), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(G286), .A2(G8), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n1129), .B(KEYINPUT123), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT51), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT51), .B1(G286), .B2(G8), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1132), .B1(new_n1128), .B2(KEYINPUT124), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT124), .ZN(new_n1134));
  AOI211_X1 g709(.A(new_n1134), .B(new_n1087), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1131), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1137));
  OR2_X1    g712(.A1(new_n1137), .A2(new_n1129), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1124), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1086), .A2(new_n1139), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1128), .A2(G168), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1096), .A2(new_n1122), .A3(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(KEYINPUT118), .A2(KEYINPUT63), .ZN(new_n1143));
  OR2_X1    g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1145));
  NAND2_X1  g720(.A1(KEYINPUT118), .A2(KEYINPUT63), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1050), .A2(G8), .ZN(new_n1148));
  XOR2_X1   g723(.A(new_n1148), .B(KEYINPUT117), .Z(new_n1149));
  NAND3_X1  g724(.A1(new_n1118), .A2(new_n1109), .A3(new_n961), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1149), .B1(new_n1113), .B2(new_n1150), .ZN(new_n1151));
  AND2_X1   g726(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1121), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1151), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1140), .A2(new_n1147), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT126), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1156), .B1(new_n1157), .B2(KEYINPUT62), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT62), .ZN(new_n1159));
  AOI211_X1 g734(.A(KEYINPUT126), .B(new_n1159), .C1(new_n1136), .C2(new_n1138), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1136), .A2(new_n1159), .A3(new_n1138), .ZN(new_n1161));
  AND4_X1   g736(.A1(G171), .A2(new_n1096), .A3(new_n1122), .A4(new_n1103), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n1158), .A2(new_n1160), .A3(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1034), .B1(new_n1155), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1029), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1166), .A2(new_n1031), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1167), .B1(new_n856), .B2(new_n864), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1168), .A2(new_n1025), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n1028), .A2(new_n806), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1025), .A2(G1996), .ZN(new_n1171));
  OAI22_X1  g746(.A1(new_n1170), .A2(new_n1025), .B1(KEYINPUT46), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1172), .B1(KEYINPUT46), .B2(new_n1171), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1173), .B(KEYINPUT47), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1025), .A2(G1986), .A3(G290), .ZN(new_n1175));
  XOR2_X1   g750(.A(new_n1175), .B(KEYINPUT48), .Z(new_n1176));
  NAND2_X1  g751(.A1(new_n1032), .A2(new_n1026), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1177), .B(KEYINPUT127), .ZN(new_n1178));
  AOI211_X1 g753(.A(new_n1169), .B(new_n1174), .C1(new_n1176), .C2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1165), .A2(new_n1179), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g755(.A(G319), .ZN(new_n1182));
  OR2_X1    g756(.A1(G227), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g757(.A(new_n1183), .B1(new_n648), .B2(new_n649), .ZN(new_n1184));
  NAND4_X1  g758(.A1(new_n1184), .A2(new_n943), .A3(new_n688), .A4(new_n692), .ZN(new_n1185));
  AOI21_X1  g759(.A(new_n1185), .B1(new_n1015), .B2(new_n1014), .ZN(G308));
  INV_X1    g760(.A(G229), .ZN(new_n1187));
  NAND4_X1  g761(.A1(new_n1187), .A2(new_n1016), .A3(new_n943), .A4(new_n1184), .ZN(G225));
endmodule


