//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 1 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 1 1 1 1 1 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n448, new_n450, new_n451, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n542, new_n543, new_n544, new_n545, new_n546, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n560, new_n562, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n609, new_n611, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1149, new_n1150, new_n1151, new_n1152;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT66), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT67), .B(G452), .ZN(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT68), .Z(G173));
  XNOR2_X1  g021(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT70), .ZN(G234));
  NAND2_X1  g027(.A1(new_n450), .A2(G2106), .ZN(G217));
  OR4_X1    g028(.A1(G221), .A2(G218), .A3(G219), .A4(G220), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT71), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n455), .A2(new_n457), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(new_n455), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2106), .ZN(new_n461));
  INV_X1    g036(.A(new_n457), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G567), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  AND2_X1   g040(.A1(KEYINPUT72), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT72), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(KEYINPUT3), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  AOI21_X1  g044(.A(KEYINPUT73), .B1(new_n469), .B2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  OAI211_X1 g046(.A(KEYINPUT73), .B(KEYINPUT3), .C1(new_n466), .C2(new_n467), .ZN(new_n472));
  AOI21_X1  g047(.A(G2105), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G137), .ZN(new_n474));
  NOR3_X1   g049(.A1(new_n466), .A2(new_n467), .A3(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  XOR2_X1   g053(.A(KEYINPUT3), .B(G2104), .Z(new_n479));
  INV_X1    g054(.A(G125), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G160));
  INV_X1    g059(.A(G2105), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n485), .B1(new_n471), .B2(new_n472), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT74), .ZN(new_n488));
  OR2_X1    g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G112), .C2(new_n485), .ZN(new_n490));
  XOR2_X1   g065(.A(new_n490), .B(KEYINPUT75), .Z(new_n491));
  AOI21_X1  g066(.A(new_n491), .B1(G136), .B2(new_n473), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR4_X1   g070(.A1(new_n479), .A2(KEYINPUT4), .A3(new_n495), .A4(G2105), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT72), .ZN(new_n497));
  INV_X1    g072(.A(G2104), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT72), .A2(G2104), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n469), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n470), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n472), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n503), .A2(G138), .A3(new_n485), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n496), .B1(new_n504), .B2(KEYINPUT4), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n503), .A2(G126), .A3(G2105), .ZN(new_n506));
  OAI21_X1  g081(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n507));
  INV_X1    g082(.A(G114), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(G2105), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n505), .A2(new_n511), .ZN(G164));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G543), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT6), .B(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(G543), .ZN(new_n521));
  INV_X1    g096(.A(G50), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n517), .A2(G62), .ZN(new_n525));
  NAND2_X1  g100(.A1(G75), .A2(G543), .ZN(new_n526));
  XOR2_X1   g101(.A(new_n526), .B(KEYINPUT76), .Z(new_n527));
  AOI21_X1  g102(.A(new_n524), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n523), .A2(new_n528), .ZN(G166));
  AND2_X1   g104(.A1(new_n517), .A2(new_n518), .ZN(new_n530));
  AND2_X1   g105(.A1(G63), .A2(G651), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n530), .A2(G89), .B1(new_n517), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n521), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G51), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT7), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n532), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT77), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n537), .A2(new_n538), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(G168));
  AOI22_X1  g116(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n524), .ZN(new_n543));
  INV_X1    g118(.A(G90), .ZN(new_n544));
  INV_X1    g119(.A(G52), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n519), .A2(new_n544), .B1(new_n521), .B2(new_n545), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n543), .A2(new_n546), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n514), .A2(new_n516), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G651), .ZN(new_n553));
  XOR2_X1   g128(.A(new_n553), .B(KEYINPUT78), .Z(new_n554));
  XOR2_X1   g129(.A(KEYINPUT79), .B(G43), .Z(new_n555));
  NAND2_X1  g130(.A1(new_n533), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n530), .A2(G81), .ZN(new_n557));
  AND3_X1   g132(.A1(new_n554), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  AND3_X1   g134(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G36), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  XOR2_X1   g139(.A(new_n564), .B(KEYINPUT80), .Z(G188));
  NAND2_X1  g140(.A1(new_n533), .A2(G53), .ZN(new_n566));
  XOR2_X1   g141(.A(new_n566), .B(KEYINPUT9), .Z(new_n567));
  AOI22_X1  g142(.A1(new_n517), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G91), .ZN(new_n569));
  OAI22_X1  g144(.A1(new_n568), .A2(new_n524), .B1(new_n519), .B2(new_n569), .ZN(new_n570));
  OR2_X1    g145(.A1(new_n567), .A2(new_n570), .ZN(G299));
  AND2_X1   g146(.A1(new_n539), .A2(new_n540), .ZN(G286));
  INV_X1    g147(.A(G166), .ZN(G303));
  INV_X1    g148(.A(G74), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n524), .B1(new_n550), .B2(new_n574), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT81), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n530), .A2(G87), .B1(new_n533), .B2(G49), .ZN(new_n577));
  AND2_X1   g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(G288));
  NAND2_X1  g154(.A1(new_n530), .A2(G86), .ZN(new_n580));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G61), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n550), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(G651), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n533), .A2(G48), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n580), .A2(new_n584), .A3(new_n585), .ZN(G305));
  AOI22_X1  g161(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n587), .A2(new_n524), .ZN(new_n588));
  INV_X1    g163(.A(G85), .ZN(new_n589));
  INV_X1    g164(.A(G47), .ZN(new_n590));
  OAI22_X1  g165(.A1(new_n519), .A2(new_n589), .B1(new_n521), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(G301), .A2(G868), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n517), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n595), .A2(new_n524), .ZN(new_n596));
  INV_X1    g171(.A(G92), .ZN(new_n597));
  OR3_X1    g172(.A1(new_n519), .A2(KEYINPUT10), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n533), .A2(G54), .ZN(new_n599));
  OAI21_X1  g174(.A(KEYINPUT10), .B1(new_n519), .B2(new_n597), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n596), .A2(new_n598), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  XOR2_X1   g176(.A(new_n601), .B(KEYINPUT82), .Z(new_n602));
  OAI21_X1  g177(.A(new_n594), .B1(new_n602), .B2(G868), .ZN(G284));
  OAI21_X1  g178(.A(new_n594), .B1(new_n602), .B2(G868), .ZN(G321));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(G299), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(new_n605), .B2(G168), .ZN(G297));
  OAI21_X1  g182(.A(new_n606), .B1(new_n605), .B2(G168), .ZN(G280));
  XOR2_X1   g183(.A(KEYINPUT83), .B(G559), .Z(new_n609));
  OAI21_X1  g184(.A(new_n602), .B1(G860), .B2(new_n609), .ZN(G148));
  NAND3_X1  g185(.A1(new_n554), .A2(new_n556), .A3(new_n557), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(new_n605), .ZN(new_n612));
  AND2_X1   g187(.A1(new_n602), .A2(new_n609), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(new_n605), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR4_X1   g190(.A1(new_n479), .A2(G2105), .A3(new_n467), .A4(new_n466), .ZN(new_n616));
  XOR2_X1   g191(.A(KEYINPUT84), .B(KEYINPUT12), .Z(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT13), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(G2100), .Z(new_n620));
  NAND2_X1  g195(.A1(new_n486), .A2(G123), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n473), .A2(G135), .ZN(new_n622));
  OR2_X1    g197(.A1(G99), .A2(G2105), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n623), .B(G2104), .C1(G111), .C2(new_n485), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n621), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(G2096), .Z(new_n626));
  NAND2_X1  g201(.A1(new_n620), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT85), .ZN(G156));
  XNOR2_X1  g203(.A(G2427), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2430), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT15), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n631), .A2(G2435), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(G2435), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n632), .A2(KEYINPUT14), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2451), .B(G2454), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT16), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n634), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2443), .B(G2446), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G1341), .B(G1348), .Z(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(G14), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n639), .A2(new_n641), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT86), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n639), .A2(KEYINPUT86), .A3(new_n641), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n644), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT87), .Z(G401));
  XOR2_X1   g225(.A(G2072), .B(G2078), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT17), .ZN(new_n652));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  XOR2_X1   g228(.A(G2067), .B(G2678), .Z(new_n654));
  NAND3_X1  g229(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT88), .ZN(new_n656));
  INV_X1    g231(.A(new_n653), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n651), .A2(new_n654), .ZN(new_n658));
  OAI211_X1 g233(.A(new_n657), .B(new_n658), .C1(new_n652), .C2(new_n654), .ZN(new_n659));
  NOR3_X1   g234(.A1(new_n657), .A2(new_n651), .A3(new_n654), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT18), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n656), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2096), .B(G2100), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(G227));
  XOR2_X1   g240(.A(G1971), .B(G1976), .Z(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G1956), .B(G2474), .Z(new_n669));
  XOR2_X1   g244(.A(G1961), .B(G1966), .Z(new_n670));
  AND2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT20), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n669), .A2(new_n670), .ZN(new_n674));
  AOI22_X1  g249(.A1(new_n672), .A2(new_n673), .B1(new_n668), .B2(new_n674), .ZN(new_n675));
  OR3_X1    g250(.A1(new_n668), .A2(new_n671), .A3(new_n674), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n675), .B(new_n676), .C1(new_n673), .C2(new_n672), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1991), .B(G1996), .ZN(new_n680));
  INV_X1    g255(.A(G1981), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(G1986), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n679), .B(new_n683), .ZN(G229));
  OAI21_X1  g259(.A(KEYINPUT98), .B1(G5), .B2(G16), .ZN(new_n685));
  OR3_X1    g260(.A1(KEYINPUT98), .A2(G5), .A3(G16), .ZN(new_n686));
  INV_X1    g261(.A(G16), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n685), .B(new_n686), .C1(G301), .C2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(G1961), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OR2_X1    g265(.A1(G29), .A2(G32), .ZN(new_n691));
  NAND3_X1  g266(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT26), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(new_n473), .B2(G141), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n486), .A2(G129), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n475), .A2(G105), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n691), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT27), .B(G1996), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n690), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G2084), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT90), .B(G29), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT24), .B(G34), .Z(new_n704));
  OAI22_X1  g279(.A1(new_n483), .A2(new_n698), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n701), .B1(new_n702), .B2(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT100), .Z(new_n707));
  NOR2_X1   g282(.A1(new_n705), .A2(new_n702), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(G168), .A2(G16), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n710), .B(KEYINPUT96), .C1(G16), .C2(G21), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(KEYINPUT96), .B2(new_n710), .ZN(new_n712));
  INV_X1    g287(.A(G1966), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n699), .A2(new_n700), .ZN(new_n715));
  INV_X1    g290(.A(new_n703), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G27), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G164), .B2(new_n716), .ZN(new_n718));
  INV_X1    g293(.A(G2078), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND4_X1  g295(.A1(new_n709), .A2(new_n714), .A3(new_n715), .A4(new_n720), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n687), .A2(KEYINPUT23), .A3(G20), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT23), .ZN(new_n723));
  INV_X1    g298(.A(G20), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(G16), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n567), .A2(new_n570), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n722), .B(new_n725), .C1(new_n726), .C2(new_n687), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G1956), .ZN(new_n728));
  NOR2_X1   g303(.A1(G16), .A2(G19), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n558), .B2(G16), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n728), .B1(G1341), .B2(new_n730), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT31), .B(G11), .ZN(new_n732));
  NAND2_X1  g307(.A1(G115), .A2(G2104), .ZN(new_n733));
  INV_X1    g308(.A(G127), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n733), .B1(new_n479), .B2(new_n734), .ZN(new_n735));
  AOI22_X1  g310(.A1(new_n473), .A2(G139), .B1(G2105), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n485), .A2(G103), .A3(G2104), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT25), .Z(new_n738));
  NAND2_X1  g313(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  MUX2_X1   g314(.A(G33), .B(new_n739), .S(G29), .Z(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(G2072), .Z(new_n741));
  INV_X1    g316(.A(new_n625), .ZN(new_n742));
  INV_X1    g317(.A(G28), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n743), .A2(KEYINPUT30), .ZN(new_n744));
  AOI21_X1  g319(.A(G29), .B1(new_n743), .B2(KEYINPUT30), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT97), .Z(new_n746));
  AOI22_X1  g321(.A1(new_n742), .A2(new_n703), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  NAND4_X1  g322(.A1(new_n731), .A2(new_n732), .A3(new_n741), .A4(new_n747), .ZN(new_n748));
  AOI22_X1  g323(.A1(G128), .A2(new_n486), .B1(new_n473), .B2(G140), .ZN(new_n749));
  OR2_X1    g324(.A1(G104), .A2(G2105), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n750), .B(G2104), .C1(G116), .C2(new_n485), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT94), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(G29), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n716), .A2(G26), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT95), .B(KEYINPUT28), .Z(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G2067), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n716), .A2(G35), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G162), .B2(new_n716), .ZN(new_n761));
  MUX2_X1   g336(.A(new_n760), .B(new_n761), .S(KEYINPUT101), .Z(new_n762));
  XOR2_X1   g337(.A(KEYINPUT29), .B(G2090), .Z(new_n763));
  XOR2_X1   g338(.A(new_n762), .B(new_n763), .Z(new_n764));
  NOR4_X1   g339(.A1(new_n721), .A2(new_n748), .A3(new_n759), .A4(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n688), .A2(new_n689), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT99), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n730), .A2(G1341), .ZN(new_n768));
  NOR2_X1   g343(.A1(G4), .A2(G16), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n602), .B2(G16), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G1348), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n765), .A2(new_n767), .A3(new_n768), .A4(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n687), .A2(G23), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n578), .B2(new_n687), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT33), .Z(new_n776));
  OR2_X1    g351(.A1(new_n776), .A2(G1976), .ZN(new_n777));
  NOR2_X1   g352(.A1(G16), .A2(G22), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G166), .B2(G16), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT92), .B(G1971), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n776), .A2(G1976), .ZN(new_n782));
  NOR2_X1   g357(.A1(G6), .A2(G16), .ZN(new_n783));
  AND3_X1   g358(.A1(new_n580), .A2(new_n584), .A3(new_n585), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(G16), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT32), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(new_n681), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n777), .A2(new_n781), .A3(new_n782), .A4(new_n787), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n788), .A2(KEYINPUT34), .ZN(new_n789));
  AOI21_X1  g364(.A(KEYINPUT93), .B1(new_n788), .B2(KEYINPUT34), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n687), .A2(G24), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n592), .B2(new_n687), .ZN(new_n792));
  INV_X1    g367(.A(G1986), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n716), .A2(G25), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n486), .A2(G119), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n473), .A2(G131), .ZN(new_n797));
  OR2_X1    g372(.A1(G95), .A2(G2105), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n798), .B(G2104), .C1(G107), .C2(new_n485), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n796), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n795), .B1(new_n801), .B2(new_n716), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT91), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT35), .B(G1991), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n789), .A2(new_n790), .A3(new_n794), .A4(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT36), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n773), .A2(new_n808), .ZN(G311));
  AND2_X1   g384(.A1(new_n765), .A2(new_n772), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n810), .A2(new_n807), .A3(new_n767), .A4(new_n768), .ZN(G150));
  INV_X1    g386(.A(G93), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT102), .B(G55), .ZN(new_n813));
  OAI22_X1  g388(.A1(new_n519), .A2(new_n812), .B1(new_n521), .B2(new_n813), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT103), .Z(new_n815));
  NAND2_X1  g390(.A1(new_n517), .A2(G67), .ZN(new_n816));
  NAND2_X1  g391(.A1(G80), .A2(G543), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n524), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(G860), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT37), .Z(new_n820));
  OAI21_X1  g395(.A(new_n558), .B1(new_n818), .B2(new_n815), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n815), .A2(new_n818), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(new_n611), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT39), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n602), .A2(G559), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT38), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n825), .B(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n820), .B1(new_n828), .B2(G860), .ZN(G145));
  XNOR2_X1  g404(.A(new_n483), .B(new_n742), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(G162), .ZN(new_n831));
  INV_X1    g406(.A(new_n496), .ZN(new_n832));
  AOI211_X1 g407(.A(new_n495), .B(G2105), .C1(new_n471), .C2(new_n472), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT4), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT104), .ZN(new_n836));
  AND3_X1   g411(.A1(new_n506), .A2(new_n836), .A3(new_n510), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n836), .B1(new_n506), .B2(new_n510), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n835), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(new_n618), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n801), .B(new_n697), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n753), .B(new_n739), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n473), .A2(G142), .ZN(new_n844));
  OAI21_X1  g419(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n485), .A2(G118), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n847), .B1(G130), .B2(new_n486), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n843), .B(new_n848), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n842), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n842), .A2(new_n849), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n831), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n852), .A2(G37), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n850), .A2(new_n851), .A3(new_n831), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(KEYINPUT105), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT105), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n850), .A2(new_n851), .A3(new_n856), .A4(new_n831), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n853), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(KEYINPUT106), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT106), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n853), .A2(new_n860), .A3(new_n855), .A4(new_n857), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g438(.A(new_n613), .B(new_n824), .ZN(new_n864));
  INV_X1    g439(.A(new_n601), .ZN(new_n865));
  NAND2_X1  g440(.A1(G299), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n726), .A2(new_n601), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n864), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n868), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(KEYINPUT41), .ZN(new_n871));
  AOI21_X1  g446(.A(KEYINPUT107), .B1(new_n726), .B2(new_n601), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n872), .B1(new_n868), .B2(KEYINPUT107), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n871), .B1(new_n873), .B2(KEYINPUT41), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n869), .B1(new_n875), .B2(new_n864), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n876), .A2(KEYINPUT42), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n592), .B(G166), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(G305), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(G288), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n876), .A2(KEYINPUT42), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n877), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n880), .B1(new_n877), .B2(new_n881), .ZN(new_n883));
  OAI21_X1  g458(.A(G868), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n884), .B1(G868), .B2(new_n822), .ZN(G295));
  OAI21_X1  g460(.A(new_n884), .B1(G868), .B2(new_n822), .ZN(G331));
  NAND2_X1  g461(.A1(G168), .A2(KEYINPUT108), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n821), .A2(new_n887), .A3(new_n823), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT108), .ZN(new_n890));
  AOI21_X1  g465(.A(G171), .B1(G286), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n887), .B1(new_n821), .B2(new_n823), .ZN(new_n893));
  NOR3_X1   g468(.A1(new_n889), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n887), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n824), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n891), .B1(new_n896), .B2(new_n888), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n868), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n891), .A3(new_n888), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n892), .B1(new_n889), .B2(new_n893), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n874), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n880), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(KEYINPUT109), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n904), .A2(new_n898), .A3(new_n901), .ZN(new_n907));
  INV_X1    g482(.A(G37), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(KEYINPUT43), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT41), .ZN(new_n911));
  OR2_X1    g486(.A1(new_n873), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n870), .A2(new_n911), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n912), .A2(new_n900), .A3(new_n899), .A4(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n914), .A2(new_n898), .A3(KEYINPUT110), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n894), .A2(new_n897), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT110), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n916), .A2(new_n917), .A3(new_n913), .A4(new_n912), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n915), .A2(new_n918), .A3(new_n903), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT43), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n898), .A2(new_n880), .A3(new_n901), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n919), .A2(new_n920), .A3(new_n908), .A4(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n910), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n909), .A2(new_n920), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n919), .A2(new_n908), .A3(new_n921), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n924), .B1(new_n925), .B2(new_n920), .ZN(new_n926));
  MUX2_X1   g501(.A(new_n923), .B(new_n926), .S(KEYINPUT44), .Z(G397));
  OR2_X1    g502(.A1(new_n753), .A2(G2067), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n753), .A2(G2067), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(G1996), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n697), .B(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  OR2_X1    g508(.A1(new_n800), .A2(new_n804), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n928), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(G1384), .ZN(new_n936));
  AOI21_X1  g511(.A(KEYINPUT45), .B1(new_n839), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n474), .A2(G40), .A3(new_n482), .A4(new_n476), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n935), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT46), .ZN(new_n942));
  INV_X1    g517(.A(new_n940), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n942), .B1(new_n943), .B2(G1996), .ZN(new_n944));
  INV_X1    g519(.A(new_n930), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n940), .B1(new_n945), .B2(new_n697), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n940), .A2(KEYINPUT46), .A3(new_n931), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n944), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(KEYINPUT127), .B(KEYINPUT47), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n948), .B(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n800), .A2(new_n804), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n930), .A2(new_n932), .A3(new_n951), .A4(new_n934), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n940), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n592), .A2(new_n793), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n943), .A2(new_n954), .ZN(new_n955));
  XOR2_X1   g530(.A(new_n955), .B(KEYINPUT48), .Z(new_n956));
  AOI211_X1 g531(.A(new_n941), .B(new_n950), .C1(new_n953), .C2(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(G301), .B(KEYINPUT54), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n936), .B1(new_n505), .B2(new_n511), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT111), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT45), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n961), .B1(new_n960), .B2(new_n962), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n511), .A2(KEYINPUT104), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n506), .A2(new_n836), .A3(new_n510), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(G1384), .B1(new_n968), .B2(new_n835), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n939), .B1(new_n969), .B2(KEYINPUT45), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n965), .A2(new_n970), .A3(new_n719), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT53), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT50), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n839), .A2(new_n973), .A3(new_n936), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n939), .B1(new_n960), .B2(KEYINPUT50), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AOI22_X1  g551(.A1(new_n971), .A2(new_n972), .B1(new_n689), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n939), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n978), .B1(new_n960), .B2(new_n962), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n719), .A2(KEYINPUT53), .ZN(new_n980));
  OR3_X1    g555(.A1(new_n937), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n959), .B1(new_n977), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n713), .B1(new_n937), .B2(new_n979), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n974), .A2(new_n975), .A3(new_n702), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(G8), .ZN(new_n986));
  NAND2_X1  g561(.A1(G286), .A2(G8), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT51), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G8), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n989), .B1(new_n983), .B2(new_n984), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n991));
  INV_X1    g566(.A(new_n987), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n990), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n988), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n987), .B1(new_n983), .B2(new_n984), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n995), .B(KEYINPUT125), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n982), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n578), .A2(G1976), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n998), .B(KEYINPUT115), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n839), .A2(new_n936), .A3(new_n978), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n1001));
  AND3_X1   g576(.A1(new_n1000), .A2(new_n1001), .A3(G8), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1001), .B1(new_n1000), .B2(G8), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n999), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT52), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1000), .A2(G8), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT114), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1000), .A2(new_n1001), .A3(G8), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G1976), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT52), .B1(G288), .B2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1009), .A2(new_n999), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT118), .ZN(new_n1013));
  XNOR2_X1  g588(.A(KEYINPUT116), .B(G1981), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n580), .A2(new_n584), .A3(new_n585), .A4(new_n1015), .ZN(new_n1016));
  OAI211_X1 g591(.A(KEYINPUT117), .B(new_n1016), .C1(new_n784), .C2(new_n681), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT117), .ZN(new_n1018));
  NAND3_X1  g593(.A1(G305), .A2(new_n1018), .A3(G1981), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT49), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1017), .A2(KEYINPUT49), .A3(new_n1019), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1013), .B1(new_n1009), .B2(new_n1024), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1013), .B(new_n1024), .C1(new_n1002), .C2(new_n1003), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1005), .B(new_n1012), .C1(new_n1025), .C2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n973), .B1(new_n839), .B2(new_n936), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n973), .B(new_n936), .C1(new_n505), .C2(new_n511), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n1029), .A2(new_n939), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G2090), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n960), .A2(new_n962), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(KEYINPUT111), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n839), .A2(KEYINPUT45), .A3(new_n936), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1036), .A2(new_n978), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G1971), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n989), .B1(new_n1034), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT120), .ZN(new_n1043));
  NOR2_X1   g618(.A1(G166), .A2(new_n989), .ZN(new_n1044));
  XNOR2_X1  g619(.A(KEYINPUT112), .B(KEYINPUT55), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(KEYINPUT112), .A2(KEYINPUT55), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1047), .B1(G166), .B2(new_n989), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n1042), .A2(new_n1043), .A3(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1028), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(G1971), .B1(new_n965), .B2(new_n970), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n976), .A2(G2090), .ZN(new_n1053));
  OAI211_X1 g628(.A(G8), .B(new_n1049), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT113), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1041), .B1(G2090), .B2(new_n976), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT113), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1056), .A2(new_n1057), .A3(G8), .A4(new_n1049), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1049), .ZN(new_n1059));
  AOI22_X1  g634(.A1(new_n1033), .A2(new_n1032), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1059), .B1(new_n1060), .B2(new_n989), .ZN(new_n1061));
  AOI22_X1  g636(.A1(new_n1055), .A2(new_n1058), .B1(new_n1061), .B2(new_n1043), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1037), .A2(new_n477), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n481), .A2(KEYINPUT126), .ZN(new_n1064));
  OAI21_X1  g639(.A(G2105), .B1(new_n481), .B2(KEYINPUT126), .ZN(new_n1065));
  OAI21_X1  g640(.A(G40), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  OR3_X1    g641(.A1(new_n937), .A2(new_n980), .A3(new_n1066), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n977), .B(new_n959), .C1(new_n1063), .C2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n997), .A2(new_n1051), .A3(new_n1062), .A4(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G1348), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n976), .A2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(G2067), .B2(new_n1000), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(new_n865), .ZN(new_n1073));
  XNOR2_X1  g648(.A(KEYINPUT56), .B(G2072), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n965), .A2(new_n970), .A3(new_n1074), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n978), .B(new_n1030), .C1(new_n969), .C2(new_n973), .ZN(new_n1076));
  INV_X1    g651(.A(G1956), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT121), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1080), .B1(new_n570), .B2(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g657(.A(new_n726), .B(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1079), .A2(KEYINPUT122), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT122), .B1(new_n1079), .B2(new_n1084), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1073), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1075), .A2(new_n1078), .A3(new_n1083), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1079), .A2(new_n1084), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT61), .B1(new_n1090), .B2(new_n1088), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT60), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1071), .B(new_n601), .C1(G2067), .C2(new_n1000), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1092), .B1(new_n1073), .B2(new_n1093), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1072), .A2(KEYINPUT60), .A3(new_n601), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n1091), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT124), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1075), .A2(new_n1078), .A3(new_n1097), .A4(new_n1083), .ZN(new_n1098));
  AND2_X1   g673(.A1(new_n1098), .A2(KEYINPUT61), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1088), .A2(KEYINPUT124), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1099), .B(new_n1100), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1101));
  XOR2_X1   g676(.A(KEYINPUT58), .B(G1341), .Z(new_n1102));
  NAND2_X1  g677(.A1(new_n1000), .A2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1103), .B1(new_n1039), .B2(G1996), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT123), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  OAI211_X1 g681(.A(KEYINPUT123), .B(new_n1103), .C1(new_n1039), .C2(G1996), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n611), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  OR2_X1    g683(.A1(new_n1108), .A2(KEYINPUT59), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(KEYINPUT59), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1096), .A2(new_n1101), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1069), .B1(new_n1089), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1028), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n990), .A2(G168), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1056), .A2(G8), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1115), .B1(new_n1116), .B2(new_n1059), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1024), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n1026), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1120), .A2(KEYINPUT119), .A3(new_n1005), .A4(new_n1012), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1114), .A2(new_n1117), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT63), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1114), .A2(new_n1121), .A3(new_n1055), .A4(new_n1058), .ZN(new_n1124));
  AOI211_X1 g699(.A(G1976), .B(G288), .C1(new_n1119), .C2(new_n1026), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1016), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1009), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1123), .A2(new_n1124), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT63), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1115), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1051), .A2(new_n1062), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT62), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n986), .A2(KEYINPUT51), .A3(new_n987), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n991), .B1(new_n990), .B2(new_n992), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n996), .A2(new_n1132), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n977), .A2(new_n981), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1051), .A2(new_n1062), .A3(new_n1135), .A4(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT125), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n995), .B(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(KEYINPUT62), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(G171), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1131), .B1(new_n1137), .B2(new_n1142), .ZN(new_n1143));
  NOR3_X1   g718(.A1(new_n1112), .A2(new_n1128), .A3(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n952), .B1(G1986), .B2(G290), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n943), .B1(new_n1145), .B2(new_n954), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n957), .B1(new_n1144), .B2(new_n1146), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g722(.A(new_n464), .B1(new_n910), .B2(new_n922), .ZN(new_n1149));
  NAND2_X1  g723(.A1(new_n649), .A2(new_n664), .ZN(new_n1150));
  AOI21_X1  g724(.A(new_n1150), .B1(new_n859), .B2(new_n861), .ZN(new_n1151));
  INV_X1    g725(.A(G229), .ZN(new_n1152));
  NAND3_X1  g726(.A1(new_n1149), .A2(new_n1151), .A3(new_n1152), .ZN(G225));
  INV_X1    g727(.A(G225), .ZN(G308));
endmodule


