//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 1 1 0 0 0 1 0 0 0 1 1 0 1 1 1 0 0 0 0 0 0 0 1 1 0 0 0 1 0 0 0 0 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n441, new_n443, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n561, new_n562, new_n564,
    new_n565, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n616, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1109, new_n1110, new_n1111;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XNOR2_X1  g015(.A(KEYINPUT64), .B(G57), .ZN(new_n441));
  INV_X1    g016(.A(new_n441), .ZN(G237));
  XNOR2_X1  g017(.A(KEYINPUT65), .B(G108), .ZN(new_n443));
  INV_X1    g018(.A(new_n443), .ZN(G238));
  NAND4_X1  g019(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NAND4_X1  g029(.A1(new_n441), .A2(new_n443), .A3(G69), .A4(G120), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT66), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n454), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OAI22_X1  g035(.A1(new_n454), .A2(new_n459), .B1(new_n460), .B2(new_n456), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT67), .Z(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n472));
  NOR3_X1   g047(.A1(new_n471), .A2(new_n472), .A3(G2105), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n470), .A2(G2105), .B1(G101), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT69), .ZN(new_n475));
  OAI21_X1  g050(.A(KEYINPUT3), .B1(new_n471), .B2(new_n472), .ZN(new_n476));
  INV_X1    g051(.A(G2105), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n476), .A2(new_n477), .A3(new_n465), .ZN(new_n478));
  INV_X1    g053(.A(G137), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n475), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n465), .ZN(new_n481));
  XNOR2_X1  g056(.A(KEYINPUT68), .B(G2104), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(new_n482), .B2(KEYINPUT3), .ZN(new_n483));
  NAND4_X1  g058(.A1(new_n483), .A2(KEYINPUT69), .A3(G137), .A4(new_n477), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n474), .A2(new_n480), .A3(new_n484), .ZN(new_n485));
  XOR2_X1   g060(.A(new_n485), .B(KEYINPUT70), .Z(G160));
  NAND2_X1  g061(.A1(new_n483), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G124), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n477), .A2(G112), .ZN(new_n490));
  OAI22_X1  g065(.A1(new_n487), .A2(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n478), .A2(KEYINPUT71), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n478), .A2(KEYINPUT71), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n491), .B1(new_n496), .B2(G136), .ZN(new_n497));
  XNOR2_X1  g072(.A(new_n497), .B(KEYINPUT72), .ZN(G162));
  NAND4_X1  g073(.A1(new_n476), .A2(G126), .A3(G2105), .A4(new_n465), .ZN(new_n499));
  OR2_X1    g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n500), .B(G2104), .C1(G114), .C2(new_n477), .ZN(new_n501));
  AND3_X1   g076(.A1(new_n499), .A2(KEYINPUT73), .A3(new_n501), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n476), .A2(G138), .A3(new_n477), .A4(new_n465), .ZN(new_n503));
  INV_X1    g078(.A(G138), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT74), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT74), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT4), .ZN(new_n508));
  AOI211_X1 g083(.A(new_n504), .B(G2105), .C1(new_n506), .C2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n468), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n503), .A2(KEYINPUT4), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AOI21_X1  g086(.A(KEYINPUT73), .B1(new_n499), .B2(new_n501), .ZN(new_n512));
  NOR3_X1   g087(.A1(new_n502), .A2(new_n511), .A3(new_n512), .ZN(G164));
  XOR2_X1   g088(.A(KEYINPUT75), .B(G651), .Z(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G651), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n515), .A2(G543), .A3(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G50), .ZN(new_n520));
  INV_X1    g095(.A(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT5), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT5), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G543), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT77), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n525), .A2(new_n526), .A3(G62), .ZN(new_n527));
  NAND2_X1  g102(.A1(G75), .A2(G543), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n522), .A2(new_n524), .ZN(new_n529));
  INV_X1    g104(.A(G62), .ZN(new_n530));
  OAI21_X1  g105(.A(KEYINPUT77), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n527), .A2(new_n528), .A3(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n514), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n515), .A2(new_n525), .A3(new_n517), .ZN(new_n535));
  XNOR2_X1  g110(.A(KEYINPUT76), .B(G88), .ZN(new_n536));
  OAI211_X1 g111(.A(new_n520), .B(new_n534), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n537), .A2(KEYINPUT78), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(KEYINPUT78), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(G166));
  AND2_X1   g115(.A1(new_n519), .A2(G51), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n525), .A2(G63), .A3(G651), .ZN(new_n542));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT7), .ZN(new_n544));
  INV_X1    g119(.A(G89), .ZN(new_n545));
  OAI211_X1 g120(.A(new_n542), .B(new_n544), .C1(new_n535), .C2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n541), .A2(new_n546), .ZN(G168));
  AOI22_X1  g122(.A1(new_n525), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(new_n514), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n549), .B1(new_n519), .B2(G52), .ZN(new_n550));
  INV_X1    g125(.A(new_n535), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G90), .ZN(new_n552));
  AND2_X1   g127(.A1(new_n550), .A2(new_n552), .ZN(G171));
  NAND2_X1  g128(.A1(new_n551), .A2(G81), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n519), .A2(G43), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n525), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n556), .A2(new_n514), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n554), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  AND3_X1   g135(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G36), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT79), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n561), .A2(new_n565), .ZN(G188));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n529), .B2(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n551), .A2(G91), .B1(G651), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT9), .ZN(new_n571));
  INV_X1    g146(.A(G53), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n518), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n519), .A2(KEYINPUT9), .A3(G53), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n570), .A2(new_n573), .A3(new_n574), .ZN(G299));
  XNOR2_X1  g150(.A(G171), .B(KEYINPUT80), .ZN(G301));
  INV_X1    g151(.A(G168), .ZN(G286));
  INV_X1    g152(.A(G166), .ZN(G303));
  OAI21_X1  g153(.A(G651), .B1(new_n525), .B2(G74), .ZN(new_n579));
  INV_X1    g154(.A(G49), .ZN(new_n580));
  INV_X1    g155(.A(G87), .ZN(new_n581));
  OAI221_X1 g156(.A(new_n579), .B1(new_n518), .B2(new_n580), .C1(new_n581), .C2(new_n535), .ZN(G288));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n529), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(new_n533), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(KEYINPUT81), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n551), .A2(G86), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT82), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n519), .A2(G48), .B1(KEYINPUT81), .B2(new_n586), .ZN(new_n591));
  OAI211_X1 g166(.A(new_n590), .B(new_n591), .C1(new_n589), .C2(new_n588), .ZN(G305));
  AOI22_X1  g167(.A1(new_n525), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  XOR2_X1   g168(.A(new_n593), .B(KEYINPUT83), .Z(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(new_n533), .ZN(new_n595));
  AOI22_X1  g170(.A1(G47), .A2(new_n519), .B1(new_n551), .B2(G85), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n529), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n519), .A2(G54), .B1(G651), .B2(new_n601), .ZN(new_n602));
  XOR2_X1   g177(.A(KEYINPUT84), .B(KEYINPUT10), .Z(new_n603));
  NAND3_X1  g178(.A1(new_n551), .A2(G92), .A3(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n603), .ZN(new_n605));
  INV_X1    g180(.A(G92), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n535), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n602), .A2(new_n604), .A3(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n598), .B1(G868), .B2(new_n609), .ZN(G284));
  OAI21_X1  g185(.A(new_n598), .B1(G868), .B2(new_n609), .ZN(G321));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(G299), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(new_n612), .B2(G168), .ZN(G297));
  OAI21_X1  g189(.A(new_n613), .B1(new_n612), .B2(G168), .ZN(G280));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n609), .B1(new_n616), .B2(G860), .ZN(G148));
  NAND2_X1  g192(.A1(new_n558), .A2(new_n612), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n608), .A2(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n612), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n622), .A2(KEYINPUT85), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(KEYINPUT85), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n623), .B(new_n624), .C1(G111), .C2(new_n477), .ZN(new_n625));
  INV_X1    g200(.A(G123), .ZN(new_n626));
  INV_X1    g201(.A(G135), .ZN(new_n627));
  OAI221_X1 g202(.A(new_n625), .B1(new_n626), .B2(new_n487), .C1(new_n495), .C2(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(G2096), .Z(new_n629));
  NAND2_X1  g204(.A1(new_n510), .A2(new_n473), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT12), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2100), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n629), .A2(new_n633), .ZN(G156));
  XOR2_X1   g209(.A(KEYINPUT15), .B(G2435), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2438), .ZN(new_n636));
  XOR2_X1   g211(.A(G2427), .B(G2430), .Z(new_n637));
  OAI21_X1  g212(.A(KEYINPUT14), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT87), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n636), .A2(new_n637), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(KEYINPUT86), .B(KEYINPUT16), .Z(new_n642));
  XNOR2_X1  g217(.A(G2443), .B(G2446), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n641), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2451), .B(G2454), .Z(new_n646));
  XOR2_X1   g221(.A(G1341), .B(G1348), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n645), .B(new_n648), .Z(new_n649));
  AND2_X1   g224(.A1(new_n649), .A2(G14), .ZN(G401));
  XOR2_X1   g225(.A(G2067), .B(G2678), .Z(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2072), .B(G2078), .Z(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT18), .Z(new_n657));
  XOR2_X1   g232(.A(KEYINPUT88), .B(KEYINPUT17), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n655), .B(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n659), .B1(new_n653), .B2(new_n652), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n655), .A2(new_n651), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n654), .B1(new_n661), .B2(new_n653), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n657), .B1(new_n660), .B2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2096), .B(G2100), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(G227));
  XOR2_X1   g241(.A(G1956), .B(G2474), .Z(new_n667));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1971), .B(G1976), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT19), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n667), .A2(new_n668), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT20), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n673), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n670), .A2(new_n672), .A3(new_n674), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n677), .B(new_n678), .C1(new_n676), .C2(new_n675), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT89), .B(G1981), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n679), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G1986), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n683), .B(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(G229));
  XOR2_X1   g262(.A(KEYINPUT92), .B(KEYINPUT28), .Z(new_n688));
  INV_X1    g263(.A(G29), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G26), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n688), .B(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(G128), .ZN(new_n692));
  OAI21_X1  g267(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n477), .A2(G116), .ZN(new_n694));
  OAI22_X1  g269(.A1(new_n487), .A2(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(new_n496), .B2(G140), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n691), .B1(new_n696), .B2(new_n689), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G2067), .ZN(new_n698));
  INV_X1    g273(.A(G19), .ZN(new_n699));
  OAI21_X1  g274(.A(KEYINPUT91), .B1(new_n699), .B2(G16), .ZN(new_n700));
  OR3_X1    g275(.A1(new_n699), .A2(KEYINPUT91), .A3(G16), .ZN(new_n701));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n700), .B(new_n701), .C1(new_n559), .C2(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(G1341), .ZN(new_n704));
  NOR2_X1   g279(.A1(G29), .A2(G32), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n473), .A2(G105), .ZN(new_n706));
  NAND3_X1  g281(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT26), .Z(new_n708));
  INV_X1    g283(.A(G129), .ZN(new_n709));
  OAI211_X1 g284(.A(new_n706), .B(new_n708), .C1(new_n487), .C2(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(new_n496), .B2(G141), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n705), .B1(new_n711), .B2(G29), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT27), .B(G1996), .Z(new_n713));
  AOI211_X1 g288(.A(new_n698), .B(new_n704), .C1(new_n712), .C2(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n712), .A2(new_n713), .ZN(new_n715));
  NOR2_X1   g290(.A1(G4), .A2(G16), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(new_n609), .B2(G16), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n717), .A2(G1348), .ZN(new_n718));
  INV_X1    g293(.A(G27), .ZN(new_n719));
  NOR3_X1   g294(.A1(new_n719), .A2(KEYINPUT96), .A3(G29), .ZN(new_n720));
  INV_X1    g295(.A(new_n502), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n503), .A2(KEYINPUT4), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n509), .A2(new_n510), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n512), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n721), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n720), .B1(new_n726), .B2(G29), .ZN(new_n727));
  OAI21_X1  g302(.A(KEYINPUT96), .B1(new_n719), .B2(G29), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI211_X1 g304(.A(new_n715), .B(new_n718), .C1(G2078), .C2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(G299), .A2(G16), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n702), .A2(KEYINPUT23), .A3(G20), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT23), .ZN(new_n733));
  INV_X1    g308(.A(G20), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n733), .B1(new_n734), .B2(G16), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n731), .A2(new_n732), .A3(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G1956), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n714), .A2(new_n730), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n496), .A2(G139), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT93), .B(KEYINPUT25), .Z(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT94), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n477), .A2(G103), .A3(G2104), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n742), .B(new_n743), .Z(new_n744));
  AOI22_X1  g319(.A1(new_n510), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n745));
  OAI211_X1 g320(.A(new_n740), .B(new_n744), .C1(new_n477), .C2(new_n745), .ZN(new_n746));
  MUX2_X1   g321(.A(G33), .B(new_n746), .S(G29), .Z(new_n747));
  NOR2_X1   g322(.A1(new_n747), .A2(G2072), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n702), .A2(G5), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G171), .B2(new_n702), .ZN(new_n750));
  INV_X1    g325(.A(G1961), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n702), .A2(G21), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G168), .B2(new_n702), .ZN(new_n754));
  INV_X1    g329(.A(G1966), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n717), .A2(G1348), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT30), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n758), .A2(G28), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(G28), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n759), .A2(new_n760), .A3(new_n689), .ZN(new_n761));
  NAND4_X1  g336(.A1(new_n752), .A2(new_n756), .A3(new_n757), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n747), .A2(G2072), .ZN(new_n763));
  OAI221_X1 g338(.A(new_n763), .B1(new_n689), .B2(new_n628), .C1(G2078), .C2(new_n729), .ZN(new_n764));
  NOR4_X1   g339(.A1(new_n739), .A2(new_n748), .A3(new_n762), .A4(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(G16), .A2(G22), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G166), .B2(G16), .ZN(new_n768));
  INV_X1    g343(.A(G1971), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  MUX2_X1   g345(.A(G6), .B(G305), .S(G16), .Z(new_n771));
  XOR2_X1   g346(.A(KEYINPUT32), .B(G1981), .Z(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(KEYINPUT90), .B1(G16), .B2(G23), .ZN(new_n774));
  OR3_X1    g349(.A1(KEYINPUT90), .A2(G16), .A3(G23), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n774), .B(new_n775), .C1(G288), .C2(new_n702), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT33), .B(G1976), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n770), .A2(new_n773), .A3(new_n778), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n779), .A2(KEYINPUT34), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(KEYINPUT34), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n702), .A2(G24), .ZN(new_n782));
  INV_X1    g357(.A(G290), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(new_n702), .ZN(new_n784));
  INV_X1    g359(.A(G1986), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n689), .A2(G25), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n496), .A2(G131), .ZN(new_n788));
  INV_X1    g363(.A(G119), .ZN(new_n789));
  OAI21_X1  g364(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n477), .A2(G107), .ZN(new_n791));
  OAI22_X1  g366(.A1(new_n487), .A2(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n787), .B1(new_n793), .B2(new_n689), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT35), .B(G1991), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n794), .B(new_n796), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n780), .A2(new_n781), .A3(new_n786), .A4(new_n797), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n798), .A2(KEYINPUT36), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(KEYINPUT36), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n766), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT95), .B(KEYINPUT31), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G11), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  OR2_X1    g379(.A1(KEYINPUT24), .A2(G34), .ZN(new_n805));
  NAND2_X1  g380(.A1(KEYINPUT24), .A2(G34), .ZN(new_n806));
  AOI21_X1  g381(.A(G29), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G160), .B2(G29), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(G2084), .Z(new_n809));
  NOR2_X1   g384(.A1(G29), .A2(G35), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(G162), .B2(G29), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT29), .B(G2090), .Z(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n801), .A2(new_n804), .A3(new_n809), .A4(new_n813), .ZN(G150));
  INV_X1    g389(.A(G150), .ZN(G311));
  NAND2_X1  g390(.A1(new_n551), .A2(G93), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n519), .A2(G55), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n525), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n816), .B(new_n817), .C1(new_n514), .C2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(G860), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT37), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n559), .B(new_n819), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n609), .A2(G559), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT39), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT98), .Z(new_n829));
  INV_X1    g404(.A(G860), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(new_n826), .B2(new_n827), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n821), .B1(new_n829), .B2(new_n831), .ZN(G145));
  XNOR2_X1  g407(.A(new_n746), .B(new_n631), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n499), .A2(new_n501), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n724), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n696), .B(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n833), .B(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(G130), .ZN(new_n838));
  OAI21_X1  g413(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n477), .A2(G118), .ZN(new_n840));
  OAI22_X1  g415(.A1(new_n487), .A2(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(new_n496), .B2(G142), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n793), .B(new_n842), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n837), .B(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(G160), .B(new_n628), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(G162), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n711), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n844), .B(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(G37), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g426(.A(new_n822), .B(new_n619), .Z(new_n852));
  XNOR2_X1  g427(.A(G299), .B(new_n608), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT41), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n853), .B(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n853), .A2(KEYINPUT41), .ZN(new_n858));
  MUX2_X1   g433(.A(new_n857), .B(new_n858), .S(KEYINPUT99), .Z(new_n859));
  AOI21_X1  g434(.A(new_n855), .B1(new_n859), .B2(new_n852), .ZN(new_n860));
  XNOR2_X1  g435(.A(G166), .B(G305), .ZN(new_n861));
  XNOR2_X1  g436(.A(G290), .B(G288), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT100), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n862), .A2(new_n863), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n861), .B1(new_n866), .B2(new_n864), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n868), .B1(KEYINPUT101), .B2(KEYINPUT42), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n860), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(KEYINPUT101), .A2(KEYINPUT42), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n860), .A2(new_n869), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n871), .B1(new_n870), .B2(new_n872), .ZN(new_n874));
  OAI21_X1  g449(.A(G868), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n819), .A2(new_n612), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(G295));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n876), .ZN(G331));
  INV_X1    g453(.A(KEYINPUT43), .ZN(new_n879));
  NAND2_X1  g454(.A1(G301), .A2(G168), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n550), .A2(new_n552), .ZN(new_n881));
  NOR2_X1   g456(.A1(G168), .A2(new_n881), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n882), .A2(KEYINPUT102), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(KEYINPUT102), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n880), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(new_n822), .Z(new_n886));
  OR2_X1    g461(.A1(new_n886), .A2(new_n859), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n854), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n887), .A2(new_n868), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(new_n849), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n868), .B1(new_n887), .B2(new_n888), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n879), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n888), .B1(new_n857), .B2(new_n886), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n893), .A2(new_n867), .A3(new_n865), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n894), .A2(new_n849), .A3(new_n889), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n892), .B1(new_n879), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(KEYINPUT44), .ZN(new_n897));
  OAI21_X1  g472(.A(KEYINPUT43), .B1(new_n890), .B2(new_n891), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n898), .B1(KEYINPUT43), .B2(new_n895), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n897), .A2(new_n901), .ZN(G397));
  AOI21_X1  g477(.A(G1384), .B1(new_n724), .B2(new_n834), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n903), .A2(KEYINPUT45), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  AND4_X1   g480(.A1(G40), .A2(new_n474), .A3(new_n480), .A4(new_n484), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n793), .A2(new_n796), .ZN(new_n910));
  NOR3_X1   g485(.A1(new_n788), .A2(new_n795), .A3(new_n792), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n909), .B1(new_n913), .B2(KEYINPUT105), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n914), .B1(KEYINPUT105), .B2(new_n913), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n696), .B(G2067), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n711), .B(G1996), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n909), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(KEYINPUT104), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n915), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n908), .A2(new_n785), .A3(new_n783), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n908), .A2(G1986), .A3(G290), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  XOR2_X1   g498(.A(new_n923), .B(KEYINPUT103), .Z(new_n924));
  NOR2_X1   g499(.A1(new_n920), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(G1384), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n726), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT45), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n907), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n903), .A2(KEYINPUT45), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n931), .B(KEYINPUT106), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n932), .A2(G1971), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT50), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n906), .B1(new_n903), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT114), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n726), .A2(new_n934), .A3(new_n926), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n906), .B(KEYINPUT114), .C1(new_n903), .C2(new_n934), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n940), .A2(G2090), .ZN(new_n941));
  OAI21_X1  g516(.A(G8), .B1(new_n933), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(G303), .A2(G8), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT55), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT107), .B1(new_n943), .B2(new_n944), .ZN(new_n946));
  OR3_X1    g521(.A1(new_n943), .A2(KEYINPUT107), .A3(new_n944), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n942), .A2(new_n945), .A3(new_n946), .A4(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G8), .ZN(new_n949));
  XOR2_X1   g524(.A(new_n931), .B(KEYINPUT106), .Z(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n769), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n907), .B1(new_n927), .B2(KEYINPUT50), .ZN(new_n952));
  INV_X1    g527(.A(new_n903), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n952), .B1(KEYINPUT50), .B2(new_n953), .ZN(new_n954));
  OR2_X1    g529(.A1(new_n954), .A2(G2090), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n949), .B1(new_n951), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n947), .A2(new_n945), .A3(new_n946), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n906), .A2(new_n903), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n960), .A2(new_n949), .ZN(new_n961));
  XNOR2_X1  g536(.A(KEYINPUT108), .B(G1976), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n961), .A2(G288), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT52), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT109), .ZN(new_n966));
  INV_X1    g541(.A(G1976), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n961), .B(new_n966), .C1(new_n967), .C2(G288), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n965), .B(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n519), .A2(G48), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n588), .A2(new_n970), .A3(new_n586), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(G1981), .ZN(new_n972));
  OAI211_X1 g547(.A(KEYINPUT110), .B(new_n972), .C1(G305), .C2(G1981), .ZN(new_n973));
  OR2_X1    g548(.A1(new_n972), .A2(KEYINPUT110), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT49), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT49), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n973), .A2(new_n977), .A3(new_n974), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n976), .A2(new_n978), .A3(new_n961), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT111), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n976), .A2(new_n981), .A3(new_n978), .A4(new_n961), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n969), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n948), .A2(new_n958), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G2078), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n932), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT53), .ZN(new_n987));
  AOI22_X1  g562(.A1(new_n986), .A2(new_n987), .B1(new_n751), .B2(new_n954), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n905), .A2(new_n906), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n927), .A2(new_n928), .ZN(new_n990));
  OR4_X1    g565(.A1(new_n987), .A2(new_n989), .A3(G2078), .A4(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n988), .A2(G301), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n989), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n993), .A2(KEYINPUT53), .A3(new_n985), .A4(new_n930), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n988), .A2(new_n994), .ZN(new_n995));
  OAI211_X1 g570(.A(KEYINPUT54), .B(new_n992), .C1(new_n995), .C2(new_n881), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT54), .ZN(new_n997));
  AND3_X1   g572(.A1(new_n988), .A2(G301), .A3(new_n994), .ZN(new_n998));
  AOI21_X1  g573(.A(G301), .B1(new_n988), .B2(new_n991), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n755), .B1(new_n989), .B2(new_n990), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1001), .B1(new_n954), .B2(G2084), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(G8), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT127), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT51), .ZN(new_n1005));
  OAI221_X1 g580(.A(new_n1003), .B1(new_n1004), .B2(new_n1005), .C1(new_n949), .C2(G168), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1007));
  OAI211_X1 g582(.A(G8), .B(new_n1007), .C1(new_n1002), .C2(G286), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1006), .B(new_n1008), .C1(KEYINPUT127), .C2(KEYINPUT51), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1003), .A2(G168), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n1010), .B(KEYINPUT126), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n984), .A2(new_n996), .A3(new_n1000), .A4(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g588(.A(KEYINPUT56), .B(G2072), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n929), .A2(KEYINPUT118), .A3(new_n930), .A4(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n928), .B1(G164), .B2(G1384), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1016), .A2(new_n906), .A3(new_n930), .A4(new_n1014), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1015), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n1021));
  AND3_X1   g596(.A1(new_n940), .A2(new_n1021), .A3(new_n737), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1021), .B1(new_n940), .B2(new_n737), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1020), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(G299), .A2(KEYINPUT117), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT57), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT116), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT117), .B1(G299), .B2(new_n1027), .ZN(new_n1028));
  MUX2_X1   g603(.A(new_n1026), .B(KEYINPUT57), .S(new_n1028), .Z(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1024), .A2(new_n1030), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1029), .B(new_n1020), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1031), .A2(KEYINPUT61), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G1996), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n929), .A2(KEYINPUT121), .A3(new_n1034), .A4(new_n930), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1016), .A2(new_n1034), .A3(new_n906), .A4(new_n930), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT121), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g613(.A(KEYINPUT58), .B(G1341), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1035), .B(new_n1038), .C1(new_n960), .C2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n559), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT59), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT59), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1040), .A2(new_n1043), .A3(new_n559), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  AND2_X1   g620(.A1(new_n1033), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT123), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1048));
  XNOR2_X1  g623(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1047), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  AOI211_X1 g626(.A(KEYINPUT123), .B(new_n1049), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1046), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT124), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NOR3_X1   g630(.A1(new_n959), .A2(KEYINPUT119), .A3(G2067), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n1057));
  INV_X1    g632(.A(G2067), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1057), .B1(new_n960), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G1348), .ZN(new_n1060));
  AOI211_X1 g635(.A(new_n1056), .B(new_n1059), .C1(new_n1060), .C2(new_n954), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n609), .A2(KEYINPUT125), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(KEYINPUT60), .A3(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n609), .A2(KEYINPUT125), .ZN(new_n1064));
  OR2_X1    g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1065), .B(new_n1066), .C1(KEYINPUT60), .C2(new_n1061), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1046), .B(KEYINPUT124), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1055), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1031), .B1(new_n608), .B2(new_n1061), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n1032), .ZN(new_n1071));
  XNOR2_X1  g646(.A(new_n1071), .B(KEYINPUT120), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1013), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1012), .A2(KEYINPUT62), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT62), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1009), .A2(new_n1011), .A3(new_n1075), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1074), .A2(new_n999), .A3(new_n984), .A4(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n980), .A2(new_n982), .ZN(new_n1078));
  NOR2_X1   g653(.A1(G288), .A2(G1976), .ZN(new_n1079));
  XOR2_X1   g654(.A(new_n1079), .B(KEYINPUT112), .Z(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(G1981), .B2(G305), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT113), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT113), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1081), .B(new_n1084), .C1(G1981), .C2(G305), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1083), .A2(new_n1085), .A3(new_n961), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n951), .B1(G2090), .B2(new_n940), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n957), .B1(new_n1087), .B2(G8), .ZN(new_n1088));
  OR3_X1    g663(.A1(new_n1003), .A2(KEYINPUT63), .A3(G286), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n958), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1003), .A2(G286), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n983), .B(new_n1091), .C1(new_n956), .C2(new_n957), .ZN(new_n1092));
  AOI22_X1  g667(.A1(new_n1090), .A2(new_n983), .B1(new_n1092), .B2(KEYINPUT63), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1077), .A2(new_n1086), .A3(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n925), .B1(new_n1073), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n908), .A2(new_n1034), .ZN(new_n1096));
  XOR2_X1   g671(.A(new_n1096), .B(KEYINPUT46), .Z(new_n1097));
  AOI21_X1  g672(.A(new_n909), .B1(new_n916), .B2(new_n711), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n1099), .B(KEYINPUT47), .ZN(new_n1100));
  XOR2_X1   g675(.A(new_n921), .B(KEYINPUT48), .Z(new_n1101));
  NOR2_X1   g676(.A1(new_n920), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n919), .A2(new_n911), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n696), .A2(new_n1058), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n909), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NOR3_X1   g680(.A1(new_n1100), .A2(new_n1102), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1095), .A2(new_n1106), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g682(.A(G319), .ZN(new_n1109));
  NOR3_X1   g683(.A1(G401), .A2(new_n1109), .A3(G227), .ZN(new_n1110));
  AND2_X1   g684(.A1(new_n850), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g685(.A1(new_n899), .A2(new_n686), .A3(new_n1111), .ZN(G225));
  INV_X1    g686(.A(G225), .ZN(G308));
endmodule


