//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 1 0 1 0 1 0 0 0 0 0 1 1 0 0 1 1 1 1 1 0 1 0 1 0 0 1 0 1 1 0 0 0 1 1 1 1 1 0 1 0 1 0 0 0 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n619, new_n620, new_n621, new_n623, new_n624,
    new_n625, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n770, new_n771,
    new_n773, new_n774, new_n775, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n832, new_n833, new_n834, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870;
  INV_X1    g000(.A(KEYINPUT92), .ZN(new_n202));
  XNOR2_X1  g001(.A(G78gat), .B(G106gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT31), .B(G50gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT29), .ZN(new_n206));
  INV_X1    g005(.A(G141gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT83), .ZN(new_n208));
  INV_X1    g007(.A(G148gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(KEYINPUT83), .A2(G148gat), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n207), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n209), .A2(G141gat), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT84), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT84), .ZN(new_n215));
  INV_X1    g014(.A(new_n213), .ZN(new_n216));
  AND2_X1   g015(.A1(KEYINPUT83), .A2(G148gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(KEYINPUT83), .A2(G148gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n215), .B(new_n216), .C1(new_n219), .C2(new_n207), .ZN(new_n220));
  AND2_X1   g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT85), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT2), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n224), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G155gat), .ZN(new_n227));
  INV_X1    g026(.A(G162gat), .ZN(new_n228));
  OAI211_X1 g027(.A(KEYINPUT85), .B(KEYINPUT2), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n223), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n214), .A2(new_n220), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT86), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT86), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n214), .A2(new_n230), .A3(new_n220), .A4(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n209), .A2(G141gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n216), .A2(new_n237), .ZN(new_n238));
  AOI211_X1 g037(.A(new_n221), .B(new_n222), .C1(new_n238), .C2(new_n225), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n235), .A2(new_n236), .A3(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n241), .A2(KEYINPUT87), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT87), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n239), .B1(new_n232), .B2(new_n234), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n243), .B1(new_n244), .B2(new_n236), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n206), .B1(new_n242), .B2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G211gat), .B(G218gat), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT76), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(G211gat), .ZN(new_n250));
  INV_X1    g049(.A(G218gat), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g051(.A1(G197gat), .A2(G204gat), .ZN(new_n253));
  AND2_X1   g052(.A1(G197gat), .A2(G204gat), .ZN(new_n254));
  OAI22_X1  g053(.A1(new_n252), .A2(KEYINPUT22), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n249), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n256), .A2(KEYINPUT77), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n249), .A2(new_n255), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n246), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n258), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n206), .B1(new_n261), .B2(new_n256), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n244), .B1(new_n236), .B2(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n263), .B1(G228gat), .B2(G233gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n260), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n236), .B1(new_n259), .B2(KEYINPUT29), .ZN(new_n266));
  INV_X1    g065(.A(new_n244), .ZN(new_n267));
  AOI22_X1  g066(.A1(new_n246), .A2(new_n259), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(G228gat), .A2(G233gat), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n265), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(G22gat), .ZN(new_n271));
  INV_X1    g070(.A(G22gat), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n265), .B(new_n272), .C1(new_n268), .C2(new_n269), .ZN(new_n273));
  AOI211_X1 g072(.A(new_n202), .B(new_n205), .C1(new_n271), .C2(new_n273), .ZN(new_n274));
  AND3_X1   g073(.A1(new_n271), .A2(new_n202), .A3(new_n273), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n202), .B1(new_n271), .B2(new_n273), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n274), .B1(new_n277), .B2(new_n205), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT34), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT70), .ZN(new_n280));
  INV_X1    g079(.A(G190gat), .ZN(new_n281));
  AND2_X1   g080(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n283));
  OAI211_X1 g082(.A(KEYINPUT28), .B(new_n281), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT68), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT27), .B(G183gat), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT68), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n286), .A2(new_n287), .A3(KEYINPUT28), .A4(new_n281), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G183gat), .ZN(new_n290));
  OAI21_X1  g089(.A(KEYINPUT27), .B1(new_n290), .B2(KEYINPUT66), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT66), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT27), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n292), .A2(new_n293), .A3(G183gat), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n291), .A2(new_n294), .A3(new_n281), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT67), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT28), .ZN(new_n297));
  AND3_X1   g096(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n296), .B1(new_n295), .B2(new_n297), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n289), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G183gat), .A2(G190gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(G169gat), .A2(G176gat), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT64), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT26), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n304), .A2(new_n305), .A3(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n300), .A2(new_n301), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT24), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n311), .A2(G183gat), .A3(G190gat), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT23), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n306), .B(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT25), .B1(new_n316), .B2(new_n301), .ZN(new_n317));
  AND3_X1   g116(.A1(new_n314), .A2(new_n317), .A3(new_n304), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT65), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n301), .A2(new_n319), .A3(new_n311), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n320), .B1(G183gat), .B2(G190gat), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n311), .B1(new_n301), .B2(new_n319), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n314), .B(new_n304), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n312), .A2(new_n318), .B1(new_n323), .B2(KEYINPUT25), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n310), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(G120gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(G113gat), .ZN(new_n327));
  INV_X1    g126(.A(G113gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(G120gat), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT1), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(G127gat), .ZN(new_n331));
  OR2_X1    g130(.A1(new_n331), .A2(KEYINPUT69), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  AOI211_X1 g132(.A(KEYINPUT1), .B(G127gat), .C1(new_n327), .C2(new_n329), .ZN(new_n334));
  OAI21_X1  g133(.A(G134gat), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n330), .A2(new_n331), .ZN(new_n336));
  INV_X1    g135(.A(G134gat), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n336), .B(new_n337), .C1(new_n330), .C2(new_n332), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n280), .B1(new_n325), .B2(new_n340), .ZN(new_n341));
  AOI211_X1 g140(.A(KEYINPUT70), .B(new_n339), .C1(new_n310), .C2(new_n324), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n310), .A2(new_n339), .A3(new_n324), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NOR3_X1   g143(.A1(new_n341), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(G227gat), .A2(G233gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT73), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n279), .B1(new_n348), .B2(KEYINPUT74), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT74), .ZN(new_n350));
  AOI211_X1 g149(.A(new_n350), .B(KEYINPUT34), .C1(new_n347), .C2(KEYINPUT73), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(KEYINPUT32), .B1(new_n345), .B2(new_n346), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n325), .A2(new_n340), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT70), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n325), .A2(new_n280), .A3(new_n340), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(new_n343), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n346), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT33), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT71), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n353), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT33), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n360), .B(new_n362), .C1(new_n345), .C2(new_n346), .ZN(new_n363));
  XNOR2_X1  g162(.A(G15gat), .B(G43gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(G71gat), .B(G99gat), .ZN(new_n365));
  XOR2_X1   g164(.A(new_n364), .B(new_n365), .Z(new_n366));
  NAND2_X1  g165(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  OR2_X1    g166(.A1(new_n361), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n366), .ZN(new_n369));
  OAI221_X1 g168(.A(KEYINPUT32), .B1(new_n362), .B2(new_n369), .C1(new_n345), .C2(new_n346), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n347), .A2(new_n350), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n352), .A2(new_n368), .A3(new_n370), .A4(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n370), .B1(new_n361), .B2(new_n367), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT72), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n348), .A2(KEYINPUT74), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT34), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n348), .A2(KEYINPUT74), .A3(new_n279), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n376), .A2(new_n371), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT72), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n379), .B(new_n370), .C1(new_n361), .C2(new_n367), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n374), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(KEYINPUT75), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT75), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n374), .A2(new_n378), .A3(new_n383), .A4(new_n380), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n278), .A2(new_n372), .A3(new_n382), .A4(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n340), .B1(new_n244), .B2(new_n236), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n241), .A2(KEYINPUT87), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n244), .A2(new_n243), .A3(new_n236), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT4), .ZN(new_n390));
  AND4_X1   g189(.A1(new_n390), .A2(new_n235), .A3(new_n240), .A4(new_n339), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n390), .B1(new_n244), .B2(new_n339), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(G225gat), .A2(G233gat), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NOR3_X1   g194(.A1(new_n389), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n244), .B(new_n339), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n395), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT5), .ZN(new_n399));
  OAI21_X1  g198(.A(KEYINPUT88), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT5), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n386), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n403), .B1(new_n242), .B2(new_n245), .ZN(new_n404));
  OR2_X1    g203(.A1(new_n391), .A2(new_n392), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(new_n405), .A3(new_n394), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT88), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n401), .B1(new_n397), .B2(new_n395), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n400), .A2(new_n402), .A3(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(KEYINPUT89), .B(KEYINPUT0), .ZN(new_n411));
  XNOR2_X1  g210(.A(G57gat), .B(G85gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(G1gat), .B(G29gat), .ZN(new_n414));
  XOR2_X1   g213(.A(new_n413), .B(new_n414), .Z(new_n415));
  NAND2_X1  g214(.A1(new_n410), .A2(new_n415), .ZN(new_n416));
  XOR2_X1   g215(.A(KEYINPUT90), .B(KEYINPUT6), .Z(new_n417));
  INV_X1    g216(.A(new_n415), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n400), .A2(new_n409), .A3(new_n418), .A4(new_n402), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n416), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT91), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OR2_X1    g221(.A1(new_n416), .A2(new_n417), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n416), .A2(KEYINPUT91), .A3(new_n417), .A4(new_n419), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT82), .B(G36gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT81), .B(G8gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(G64gat), .B(G92gat), .ZN(new_n429));
  XOR2_X1   g228(.A(new_n428), .B(new_n429), .Z(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n325), .A2(KEYINPUT78), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT78), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n310), .A2(new_n433), .A3(new_n324), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT29), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(G226gat), .A2(G233gat), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT79), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n434), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n433), .B1(new_n310), .B2(new_n324), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n206), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT79), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n441), .A2(new_n442), .A3(new_n436), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n325), .A2(new_n437), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n438), .A2(new_n443), .A3(new_n259), .A4(new_n444), .ZN(new_n445));
  NOR3_X1   g244(.A1(new_n439), .A2(new_n436), .A3(new_n440), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n437), .A2(KEYINPUT29), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n446), .B1(new_n325), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n259), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AND3_X1   g249(.A1(new_n445), .A2(new_n450), .A3(KEYINPUT80), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT80), .B1(new_n445), .B2(new_n450), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n431), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n431), .B1(new_n445), .B2(new_n450), .ZN(new_n454));
  OR2_X1    g253(.A1(new_n454), .A2(KEYINPUT30), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(KEYINPUT30), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n453), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n425), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(KEYINPUT35), .B1(new_n385), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n378), .A2(new_n373), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n372), .A2(new_n461), .ZN(new_n462));
  XOR2_X1   g261(.A(KEYINPUT95), .B(KEYINPUT35), .Z(new_n463));
  AOI21_X1  g262(.A(new_n463), .B1(new_n423), .B2(new_n420), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n278), .A2(new_n462), .A3(new_n458), .A4(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT36), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n372), .A2(new_n461), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n382), .A2(new_n372), .A3(new_n384), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n468), .B1(new_n469), .B2(KEYINPUT36), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n277), .A2(new_n205), .ZN(new_n471));
  INV_X1    g270(.A(new_n274), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n459), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n397), .A2(new_n395), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT93), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT93), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n404), .A2(new_n405), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n477), .B1(new_n478), .B2(new_n395), .ZN(new_n479));
  OAI211_X1 g278(.A(KEYINPUT39), .B(new_n476), .C1(new_n479), .C2(new_n475), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT39), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n478), .A2(new_n481), .A3(new_n395), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n480), .A2(new_n418), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT40), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(KEYINPUT94), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(KEYINPUT94), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n480), .A2(new_n418), .A3(new_n486), .A4(new_n482), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n457), .A2(new_n416), .A3(new_n485), .A4(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT38), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT37), .B1(new_n451), .B2(new_n452), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n445), .A2(new_n450), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT37), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n489), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n438), .A2(new_n443), .A3(new_n444), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n492), .B1(new_n495), .B2(new_n449), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n496), .B1(new_n449), .B2(new_n448), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n497), .A2(new_n489), .A3(new_n431), .A4(new_n493), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n430), .B1(new_n491), .B2(KEYINPUT38), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n423), .A2(new_n498), .A3(new_n420), .A4(new_n499), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n278), .B(new_n488), .C1(new_n494), .C2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n470), .A2(new_n474), .A3(new_n501), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n466), .A2(KEYINPUT96), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT96), .B1(new_n466), .B2(new_n502), .ZN(new_n504));
  OR2_X1    g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(G8gat), .ZN(new_n506));
  XOR2_X1   g305(.A(G15gat), .B(G22gat), .Z(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  OR2_X1    g307(.A1(new_n508), .A2(G1gat), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT98), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT16), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n508), .B1(new_n512), .B2(G1gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  OR2_X1    g313(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n511), .A2(new_n514), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT21), .ZN(new_n517));
  XNOR2_X1  g316(.A(G57gat), .B(G64gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n518), .B(KEYINPUT99), .ZN(new_n519));
  NAND2_X1  g318(.A1(G71gat), .A2(G78gat), .ZN(new_n520));
  OR2_X1    g319(.A1(G71gat), .A2(G78gat), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT9), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n520), .B(new_n521), .C1(new_n518), .C2(new_n522), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n515), .B(new_n516), .C1(new_n517), .C2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(new_n290), .ZN(new_n528));
  NAND2_X1  g327(.A1(G231gat), .A2(G233gat), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n528), .B(new_n529), .Z(new_n530));
  XOR2_X1   g329(.A(G127gat), .B(G155gat), .Z(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(KEYINPUT20), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n530), .B(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n526), .A2(new_n517), .ZN(new_n534));
  XNOR2_X1  g333(.A(KEYINPUT100), .B(KEYINPUT19), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(new_n250), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n534), .B(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n533), .B(new_n537), .ZN(new_n538));
  XOR2_X1   g337(.A(G190gat), .B(G218gat), .Z(new_n539));
  NOR2_X1   g338(.A1(new_n539), .A2(KEYINPUT101), .ZN(new_n540));
  OR3_X1    g339(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n541));
  OAI21_X1  g340(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n541), .A2(new_n542), .B1(G29gat), .B2(G36gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(G43gat), .B(G50gat), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n543), .B1(KEYINPUT15), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(KEYINPUT15), .ZN(new_n546));
  XOR2_X1   g345(.A(new_n545), .B(new_n546), .Z(new_n547));
  NAND2_X1  g346(.A1(G85gat), .A2(G92gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT7), .ZN(new_n549));
  NAND2_X1  g348(.A1(G99gat), .A2(G106gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT8), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n549), .B(new_n551), .C1(G85gat), .C2(G92gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(G99gat), .B(G106gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n540), .B1(new_n547), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT41), .ZN(new_n556));
  NAND2_X1  g355(.A1(G232gat), .A2(G233gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n547), .B(KEYINPUT17), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  OAI221_X1 g358(.A(new_n555), .B1(new_n556), .B2(new_n557), .C1(new_n559), .C2(new_n554), .ZN(new_n560));
  XNOR2_X1  g359(.A(G134gat), .B(G162gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n539), .A2(KEYINPUT101), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n557), .A2(new_n556), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n562), .B(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n538), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n505), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n515), .A2(new_n516), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n559), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n571), .B1(new_n570), .B2(new_n547), .ZN(new_n572));
  NAND2_X1  g371(.A1(G229gat), .A2(G233gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT18), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n570), .B(new_n547), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n573), .B(KEYINPUT13), .Z(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(KEYINPUT97), .B(KEYINPUT11), .ZN(new_n580));
  XNOR2_X1  g379(.A(G169gat), .B(G197gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G113gat), .B(G141gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n584), .B(KEYINPUT12), .Z(new_n585));
  OR2_X1    g384(.A1(new_n579), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n579), .A2(new_n585), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n554), .B(new_n526), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT10), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n554), .A2(KEYINPUT10), .A3(new_n524), .A4(new_n525), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G230gat), .A2(G233gat), .ZN(new_n595));
  AND2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n590), .A2(new_n595), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G120gat), .B(G148gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(G176gat), .B(G204gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT102), .B1(new_n598), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n603), .B1(new_n598), .B2(new_n602), .ZN(new_n604));
  OAI211_X1 g403(.A(KEYINPUT102), .B(new_n601), .C1(new_n596), .C2(new_n597), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n589), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n569), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n425), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g412(.A1(new_n609), .A2(new_n458), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n614), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n615), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n616), .B(KEYINPUT42), .Z(new_n617));
  OAI21_X1  g416(.A(new_n617), .B1(new_n506), .B2(new_n614), .ZN(G1325gat));
  INV_X1    g417(.A(new_n470), .ZN(new_n619));
  AND3_X1   g418(.A1(new_n610), .A2(G15gat), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(G15gat), .B1(new_n610), .B2(new_n462), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(G1326gat));
  NOR2_X1   g421(.A1(new_n609), .A2(new_n278), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(new_n272), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT103), .B(KEYINPUT43), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(G1327gat));
  INV_X1    g425(.A(new_n538), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n608), .A2(new_n627), .ZN(new_n628));
  NOR3_X1   g427(.A1(new_n505), .A2(new_n567), .A3(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NOR3_X1   g429(.A1(new_n630), .A2(G29gat), .A3(new_n425), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n631), .B(KEYINPUT104), .Z(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT45), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT108), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT107), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n502), .A2(KEYINPUT105), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT105), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n470), .A2(new_n474), .A3(new_n637), .A4(new_n501), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n636), .A2(new_n466), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT106), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n636), .A2(new_n466), .A3(KEYINPUT106), .A4(new_n638), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n567), .A2(KEYINPUT44), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n635), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n644), .ZN(new_n646));
  AOI211_X1 g445(.A(KEYINPUT107), .B(new_n646), .C1(new_n641), .C2(new_n642), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT44), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n503), .A2(new_n504), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n648), .B1(new_n649), .B2(new_n566), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n645), .A2(new_n647), .A3(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n634), .B1(new_n651), .B2(new_n628), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n643), .A2(new_n644), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(KEYINPUT107), .ZN(new_n654));
  INV_X1    g453(.A(new_n650), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n643), .A2(new_n635), .A3(new_n644), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n628), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n657), .A2(KEYINPUT108), .A3(new_n658), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n652), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(G29gat), .B1(new_n660), .B2(new_n425), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n633), .A2(new_n661), .ZN(G1328gat));
  OAI21_X1  g461(.A(G36gat), .B1(new_n660), .B2(new_n458), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n630), .A2(G36gat), .A3(new_n458), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT46), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n665), .ZN(G1329gat));
  INV_X1    g465(.A(new_n462), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n630), .A2(G43gat), .A3(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n657), .A2(new_n619), .A3(new_n658), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n668), .B1(new_n669), .B2(G43gat), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(KEYINPUT47), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n660), .A2(new_n470), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n668), .B1(new_n672), .B2(G43gat), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n671), .B1(new_n673), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g473(.A(G50gat), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n629), .A2(new_n675), .A3(new_n473), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n651), .A2(new_n278), .A3(new_n628), .ZN(new_n677));
  OAI211_X1 g476(.A(KEYINPUT48), .B(new_n676), .C1(new_n677), .C2(new_n675), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n278), .B1(new_n652), .B2(new_n659), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n676), .B1(new_n679), .B2(new_n675), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT109), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT48), .ZN(new_n682));
  AND3_X1   g481(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n681), .B1(new_n680), .B2(new_n682), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n678), .B1(new_n683), .B2(new_n684), .ZN(G1331gat));
  NOR2_X1   g484(.A1(new_n568), .A2(new_n588), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n643), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n607), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n611), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(G57gat), .ZN(G1332gat));
  AOI211_X1 g490(.A(new_n458), .B(new_n688), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n692));
  NOR2_X1   g491(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1333gat));
  OAI21_X1  g493(.A(G71gat), .B1(new_n688), .B2(new_n470), .ZN(new_n695));
  OR2_X1    g494(.A1(new_n667), .A2(G71gat), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n695), .B1(new_n688), .B2(new_n696), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n697), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g497(.A1(new_n689), .A2(new_n473), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g499(.A1(new_n588), .A2(new_n538), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n657), .A2(new_n607), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n702), .A2(G85gat), .A3(new_n611), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n639), .A2(new_n566), .A3(new_n701), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT51), .ZN(new_n705));
  OR2_X1    g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n705), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n706), .A2(KEYINPUT110), .A3(new_n707), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n707), .A2(KEYINPUT110), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n708), .A2(new_n607), .A3(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n710), .A2(new_n425), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n703), .B1(G85gat), .B2(new_n711), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n712), .B(KEYINPUT111), .Z(G1336gat));
  NAND2_X1  g512(.A1(new_n702), .A2(new_n457), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(G92gat), .ZN(new_n715));
  INV_X1    g514(.A(new_n710), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n458), .A2(G92gat), .ZN(new_n717));
  AOI21_X1  g516(.A(KEYINPUT52), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n704), .A2(KEYINPUT112), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(new_n705), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n721), .A2(new_n606), .ZN(new_n722));
  AOI22_X1  g521(.A1(new_n714), .A2(G92gat), .B1(new_n717), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT52), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n719), .B1(new_n723), .B2(new_n724), .ZN(G1337gat));
  XOR2_X1   g524(.A(KEYINPUT113), .B(G99gat), .Z(new_n726));
  NOR3_X1   g525(.A1(new_n710), .A2(new_n667), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n702), .A2(new_n619), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n727), .B1(new_n728), .B2(new_n726), .ZN(new_n729));
  XOR2_X1   g528(.A(new_n729), .B(KEYINPUT114), .Z(G1338gat));
  NAND2_X1  g529(.A1(new_n702), .A2(new_n473), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(G106gat), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n278), .A2(G106gat), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT53), .ZN(new_n734));
  AOI22_X1  g533(.A1(new_n716), .A2(new_n733), .B1(KEYINPUT115), .B2(new_n734), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n732), .B(new_n735), .C1(KEYINPUT115), .C2(new_n734), .ZN(new_n736));
  AOI22_X1  g535(.A1(new_n731), .A2(G106gat), .B1(new_n722), .B2(new_n733), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n736), .B1(new_n737), .B2(new_n734), .ZN(G1339gat));
  INV_X1    g537(.A(KEYINPUT54), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n602), .B1(new_n596), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(KEYINPUT54), .B1(new_n594), .B2(new_n595), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n596), .B2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT55), .ZN(new_n743));
  OR2_X1    g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n598), .A2(new_n602), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT116), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n742), .A2(new_n743), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n588), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n572), .A2(new_n573), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n576), .A2(new_n577), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n584), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n586), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n607), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n566), .B1(new_n751), .B2(new_n756), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n750), .A2(new_n566), .A3(new_n755), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n627), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n686), .A2(new_n606), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n761), .A2(new_n425), .A3(new_n385), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n762), .A2(new_n458), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n763), .A2(new_n328), .A3(new_n588), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n761), .A2(new_n425), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n765), .A2(new_n462), .A3(new_n458), .A4(new_n278), .ZN(new_n766));
  OAI21_X1  g565(.A(G113gat), .B1(new_n766), .B2(new_n589), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n764), .A2(new_n767), .ZN(G1340gat));
  OAI21_X1  g567(.A(G120gat), .B1(new_n766), .B2(new_n606), .ZN(new_n769));
  XOR2_X1   g568(.A(new_n769), .B(KEYINPUT117), .Z(new_n770));
  NAND3_X1  g569(.A1(new_n763), .A2(new_n326), .A3(new_n607), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(G1341gat));
  NOR3_X1   g571(.A1(new_n766), .A2(new_n331), .A3(new_n627), .ZN(new_n773));
  XOR2_X1   g572(.A(new_n773), .B(KEYINPUT118), .Z(new_n774));
  AOI21_X1  g573(.A(G127gat), .B1(new_n763), .B2(new_n538), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n774), .A2(new_n775), .ZN(G1342gat));
  NOR2_X1   g575(.A1(new_n567), .A2(new_n457), .ZN(new_n777));
  XNOR2_X1  g576(.A(KEYINPUT69), .B(G134gat), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n762), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  XOR2_X1   g578(.A(new_n779), .B(KEYINPUT56), .Z(new_n780));
  OAI21_X1  g579(.A(G134gat), .B1(new_n766), .B2(new_n567), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(G1343gat));
  AOI21_X1  g581(.A(new_n278), .B1(new_n759), .B2(new_n760), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n619), .A2(new_n425), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n458), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n207), .B1(new_n787), .B2(new_n589), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT119), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT57), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n783), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n588), .A2(new_n745), .A3(new_n749), .A4(new_n744), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n566), .B1(new_n756), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n627), .B1(new_n758), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n278), .B1(new_n794), .B2(new_n760), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n791), .B(new_n786), .C1(new_n790), .C2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n588), .A2(G141gat), .ZN(new_n797));
  OAI221_X1 g596(.A(new_n788), .B1(new_n789), .B2(KEYINPUT58), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n789), .A2(KEYINPUT58), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n798), .B(new_n799), .ZN(G1344gat));
  INV_X1    g599(.A(KEYINPUT59), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n801), .B(new_n219), .C1(new_n796), .C2(new_n606), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n783), .A2(KEYINPUT57), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n795), .A2(KEYINPUT57), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n607), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n209), .B1(new_n806), .B2(new_n786), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n802), .B1(new_n807), .B2(new_n801), .ZN(new_n808));
  OR3_X1    g607(.A1(new_n787), .A2(new_n219), .A3(new_n606), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT120), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n810), .B(new_n811), .ZN(G1345gat));
  OAI21_X1  g611(.A(new_n227), .B1(new_n787), .B2(new_n627), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n538), .A2(G155gat), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n796), .B2(new_n814), .ZN(new_n815));
  XOR2_X1   g614(.A(new_n815), .B(KEYINPUT121), .Z(G1346gat));
  NAND4_X1  g615(.A1(new_n783), .A2(new_n228), .A3(new_n777), .A4(new_n784), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n796), .A2(new_n567), .ZN(new_n818));
  XOR2_X1   g617(.A(new_n818), .B(KEYINPUT122), .Z(new_n819));
  OAI21_X1  g618(.A(new_n817), .B1(new_n819), .B2(new_n228), .ZN(G1347gat));
  NOR2_X1   g619(.A1(new_n611), .A2(new_n458), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  OR4_X1    g621(.A1(new_n667), .A2(new_n761), .A3(new_n473), .A4(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(G169gat), .B1(new_n823), .B2(new_n589), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n385), .A2(new_n458), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n825), .A2(KEYINPUT123), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n825), .A2(KEYINPUT123), .ZN(new_n827));
  NOR4_X1   g626(.A1(new_n761), .A2(new_n611), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(G169gat), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n828), .A2(new_n829), .A3(new_n588), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n824), .A2(new_n830), .ZN(G1348gat));
  INV_X1    g630(.A(G176gat), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n823), .A2(new_n832), .A3(new_n606), .ZN(new_n833));
  AOI21_X1  g632(.A(G176gat), .B1(new_n828), .B2(new_n607), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n833), .A2(new_n834), .ZN(G1349gat));
  NOR2_X1   g634(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n836));
  OAI21_X1  g635(.A(G183gat), .B1(new_n823), .B2(new_n627), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n828), .A2(new_n286), .A3(new_n538), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n840));
  XOR2_X1   g639(.A(new_n839), .B(new_n840), .Z(G1350gat));
  INV_X1    g640(.A(KEYINPUT61), .ZN(new_n842));
  OAI221_X1 g641(.A(G190gat), .B1(KEYINPUT125), .B2(new_n842), .C1(new_n823), .C2(new_n567), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(KEYINPUT125), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n828), .A2(new_n281), .A3(new_n566), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(G1351gat));
  NOR2_X1   g646(.A1(new_n619), .A2(new_n822), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n783), .A2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(G197gat), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n849), .A2(new_n850), .A3(new_n588), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n803), .A2(new_n804), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n852), .A2(new_n848), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n853), .A2(new_n588), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n851), .B1(new_n854), .B2(new_n850), .ZN(G1352gat));
  XNOR2_X1  g654(.A(KEYINPUT126), .B(G204gat), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n849), .A2(new_n607), .A3(new_n856), .ZN(new_n857));
  XOR2_X1   g656(.A(new_n857), .B(KEYINPUT62), .Z(new_n858));
  NOR3_X1   g657(.A1(new_n805), .A2(new_n619), .A3(new_n822), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n858), .B1(new_n859), .B2(new_n856), .ZN(G1353gat));
  NAND2_X1  g659(.A1(new_n853), .A2(new_n538), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(G211gat), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n862), .A2(KEYINPUT127), .A3(KEYINPUT63), .ZN(new_n863));
  OR2_X1    g662(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n864));
  NAND2_X1  g663(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n861), .A2(G211gat), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n849), .A2(new_n250), .A3(new_n538), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n863), .A2(new_n866), .A3(new_n867), .ZN(G1354gat));
  AOI21_X1  g667(.A(G218gat), .B1(new_n849), .B2(new_n566), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n567), .A2(new_n251), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n869), .B1(new_n853), .B2(new_n870), .ZN(G1355gat));
endmodule


