

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746;

  INV_X1 U376 ( .A(n591), .ZN(n681) );
  NOR2_X1 U377 ( .A1(G953), .A2(G237), .ZN(n516) );
  XNOR2_X1 U378 ( .A(G119), .B(G113), .ZN(n479) );
  AND2_X1 U379 ( .A1(n363), .A2(n617), .ZN(n395) );
  XNOR2_X1 U380 ( .A(KEYINPUT38), .B(n609), .ZN(n676) );
  INV_X1 U381 ( .A(G953), .ZN(n370) );
  AND2_X2 U382 ( .A1(n414), .A2(n413), .ZN(n406) );
  AND2_X4 U383 ( .A1(n395), .A2(n656), .ZN(n715) );
  XNOR2_X2 U384 ( .A(n616), .B(KEYINPUT73), .ZN(n656) );
  XNOR2_X2 U385 ( .A(n499), .B(n410), .ZN(n704) );
  NOR2_X1 U386 ( .A1(n660), .A2(n527), .ZN(n528) );
  NOR2_X1 U387 ( .A1(n545), .A2(n418), .ZN(n372) );
  NAND2_X1 U388 ( .A1(n399), .A2(n400), .ZN(n601) );
  XNOR2_X1 U389 ( .A(n542), .B(KEYINPUT32), .ZN(n744) );
  XNOR2_X1 U390 ( .A(n372), .B(n371), .ZN(n632) );
  NOR2_X1 U391 ( .A1(n679), .A2(n682), .ZN(n571) );
  XNOR2_X1 U392 ( .A(n577), .B(KEYINPUT1), .ZN(n660) );
  XNOR2_X1 U393 ( .A(n512), .B(n511), .ZN(n664) );
  XNOR2_X1 U394 ( .A(n398), .B(n354), .ZN(n549) );
  OR2_X1 U395 ( .A1(n711), .A2(G902), .ZN(n398) );
  XNOR2_X1 U396 ( .A(n711), .B(n710), .ZN(n712) );
  XNOR2_X1 U397 ( .A(n733), .B(G146), .ZN(n525) );
  XNOR2_X1 U398 ( .A(n494), .B(n403), .ZN(n733) );
  XNOR2_X1 U399 ( .A(n493), .B(G134), .ZN(n403) );
  XNOR2_X1 U400 ( .A(n402), .B(G146), .ZN(n484) );
  XNOR2_X1 U401 ( .A(n487), .B(KEYINPUT4), .ZN(n494) );
  INV_X1 U402 ( .A(n373), .ZN(n480) );
  XOR2_X1 U403 ( .A(KEYINPUT12), .B(KEYINPUT101), .Z(n456) );
  XNOR2_X1 U404 ( .A(G101), .B(KEYINPUT3), .ZN(n373) );
  INV_X1 U405 ( .A(G125), .ZN(n402) );
  NOR2_X1 U406 ( .A1(n743), .A2(KEYINPUT65), .ZN(n385) );
  XNOR2_X1 U407 ( .A(n484), .B(n453), .ZN(n458) );
  XNOR2_X1 U408 ( .A(KEYINPUT10), .B(G140), .ZN(n453) );
  INV_X1 U409 ( .A(n572), .ZN(n397) );
  OR2_X2 U410 ( .A1(n621), .A2(G902), .ZN(n430) );
  XNOR2_X1 U411 ( .A(G122), .B(G104), .ZN(n483) );
  INV_X1 U412 ( .A(KEYINPUT81), .ZN(n379) );
  INV_X1 U413 ( .A(KEYINPUT0), .ZN(n428) );
  AND2_X1 U414 ( .A1(n377), .A2(n358), .ZN(n399) );
  XNOR2_X1 U415 ( .A(n600), .B(n599), .ZN(n400) );
  XNOR2_X1 U416 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n579) );
  INV_X1 U417 ( .A(KEYINPUT48), .ZN(n441) );
  NOR2_X1 U418 ( .A1(n601), .A2(n441), .ZN(n438) );
  AND2_X1 U419 ( .A1(n559), .A2(n408), .ZN(n407) );
  INV_X1 U420 ( .A(KEYINPUT44), .ZN(n408) );
  XOR2_X1 U421 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n464) );
  XNOR2_X1 U422 ( .A(n501), .B(n500), .ZN(n504) );
  XNOR2_X1 U423 ( .A(G140), .B(G101), .ZN(n500) );
  XNOR2_X1 U424 ( .A(n497), .B(G107), .ZN(n498) );
  XNOR2_X1 U425 ( .A(n409), .B(G469), .ZN(n577) );
  INV_X1 U426 ( .A(n515), .ZN(n659) );
  NOR2_X1 U427 ( .A1(n664), .A2(n536), .ZN(n515) );
  XNOR2_X1 U428 ( .A(n525), .B(n526), .ZN(n621) );
  INV_X1 U429 ( .A(n483), .ZN(n401) );
  INV_X1 U430 ( .A(KEYINPUT67), .ZN(n404) );
  XNOR2_X1 U431 ( .A(n721), .B(n488), .ZN(n700) );
  XNOR2_X1 U432 ( .A(n486), .B(n382), .ZN(n488) );
  XNOR2_X1 U433 ( .A(n484), .B(n424), .ZN(n486) );
  XNOR2_X1 U434 ( .A(n494), .B(n485), .ZN(n382) );
  XNOR2_X1 U435 ( .A(n631), .B(n552), .ZN(n612) );
  XNOR2_X1 U436 ( .A(n471), .B(G478), .ZN(n553) );
  INV_X1 U437 ( .A(n659), .ZN(n419) );
  INV_X1 U438 ( .A(KEYINPUT90), .ZN(n492) );
  INV_X1 U439 ( .A(KEYINPUT65), .ZN(n534) );
  NAND2_X1 U440 ( .A1(n744), .A2(n636), .ZN(n374) );
  XOR2_X1 U441 ( .A(KEYINPUT95), .B(KEYINPUT20), .Z(n508) );
  INV_X1 U442 ( .A(KEYINPUT72), .ZN(n519) );
  XNOR2_X1 U443 ( .A(G137), .B(KEYINPUT68), .ZN(n495) );
  XNOR2_X1 U444 ( .A(n426), .B(n425), .ZN(n424) );
  XNOR2_X1 U445 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n426) );
  XNOR2_X1 U446 ( .A(KEYINPUT87), .B(KEYINPUT85), .ZN(n425) );
  NAND2_X1 U447 ( .A1(G237), .A2(G234), .ZN(n473) );
  AND2_X1 U448 ( .A1(n602), .A2(n441), .ZN(n391) );
  INV_X1 U449 ( .A(KEYINPUT45), .ZN(n411) );
  NOR2_X1 U450 ( .A1(G237), .A2(G902), .ZN(n478) );
  XNOR2_X1 U451 ( .A(G119), .B(G110), .ZN(n444) );
  XOR2_X1 U452 ( .A(KEYINPUT66), .B(KEYINPUT8), .Z(n451) );
  XOR2_X1 U453 ( .A(KEYINPUT103), .B(KEYINPUT102), .Z(n442) );
  XNOR2_X1 U454 ( .A(G122), .B(G134), .ZN(n463) );
  XOR2_X1 U455 ( .A(G902), .B(KEYINPUT15), .Z(n617) );
  INV_X1 U456 ( .A(n618), .ZN(n727) );
  XNOR2_X1 U457 ( .A(n505), .B(n498), .ZN(n410) );
  XNOR2_X1 U458 ( .A(n504), .B(n503), .ZN(n505) );
  AND2_X1 U459 ( .A1(n568), .A2(n432), .ZN(n587) );
  NOR2_X1 U460 ( .A1(n659), .A2(n396), .ZN(n432) );
  XNOR2_X1 U461 ( .A(n539), .B(KEYINPUT22), .ZN(n555) );
  XNOR2_X1 U462 ( .A(n621), .B(KEYINPUT62), .ZN(n623) );
  XNOR2_X1 U463 ( .A(n376), .B(n482), .ZN(n721) );
  XNOR2_X1 U464 ( .A(G113), .B(G143), .ZN(n454) );
  XNOR2_X1 U465 ( .A(n578), .B(KEYINPUT42), .ZN(n746) );
  INV_X1 U466 ( .A(KEYINPUT40), .ZN(n394) );
  XNOR2_X1 U467 ( .A(n368), .B(n367), .ZN(n586) );
  INV_X1 U468 ( .A(KEYINPUT36), .ZN(n367) );
  NOR2_X1 U469 ( .A1(n603), .A2(n585), .ZN(n368) );
  INV_X1 U470 ( .A(KEYINPUT35), .ZN(n532) );
  XNOR2_X1 U471 ( .A(n417), .B(n416), .ZN(n646) );
  XNOR2_X1 U472 ( .A(KEYINPUT99), .B(KEYINPUT31), .ZN(n416) );
  NAND2_X1 U473 ( .A1(n427), .A2(n355), .ZN(n417) );
  AND2_X1 U474 ( .A1(n547), .A2(n387), .ZN(n427) );
  XNOR2_X1 U475 ( .A(n594), .B(n378), .ZN(n637) );
  INV_X1 U476 ( .A(KEYINPUT77), .ZN(n378) );
  NOR2_X1 U477 ( .A1(n549), .A2(n553), .ZN(n551) );
  INV_X1 U478 ( .A(KEYINPUT98), .ZN(n371) );
  NAND2_X1 U479 ( .A1(n546), .A2(n419), .ZN(n418) );
  XNOR2_X1 U480 ( .A(n716), .B(n362), .ZN(n718) );
  XNOR2_X1 U481 ( .A(n717), .B(KEYINPUT122), .ZN(n362) );
  INV_X1 U482 ( .A(KEYINPUT56), .ZN(n383) );
  AND2_X1 U483 ( .A1(n697), .A2(n369), .ZN(n386) );
  AND2_X1 U484 ( .A1(n696), .A2(n370), .ZN(n369) );
  XOR2_X1 U485 ( .A(KEYINPUT13), .B(G475), .Z(n354) );
  NOR2_X1 U486 ( .A1(n659), .A2(n660), .ZN(n355) );
  XOR2_X1 U487 ( .A(n393), .B(n445), .Z(n356) );
  AND2_X1 U488 ( .A1(G210), .A2(n489), .ZN(n357) );
  AND2_X1 U489 ( .A1(n596), .A2(n595), .ZN(n358) );
  XOR2_X1 U490 ( .A(n743), .B(n534), .Z(n359) );
  AND2_X1 U491 ( .A1(n614), .A2(KEYINPUT2), .ZN(n360) );
  NOR2_X1 U492 ( .A1(G952), .A2(n370), .ZN(n719) );
  INV_X1 U493 ( .A(n719), .ZN(n388) );
  NAND2_X1 U494 ( .A1(n745), .A2(n746), .ZN(n580) );
  XNOR2_X1 U495 ( .A(n570), .B(n394), .ZN(n745) );
  NAND2_X1 U496 ( .A1(n365), .A2(n364), .ZN(n363) );
  XNOR2_X1 U497 ( .A(n380), .B(n379), .ZN(n615) );
  NAND2_X1 U498 ( .A1(n433), .A2(n397), .ZN(n396) );
  NOR2_X1 U499 ( .A1(n704), .A2(G902), .ZN(n409) );
  NOR2_X2 U500 ( .A1(n618), .A2(n615), .ZN(n616) );
  NAND2_X1 U501 ( .A1(n361), .A2(KEYINPUT44), .ZN(n414) );
  NAND2_X1 U502 ( .A1(n559), .A2(n385), .ZN(n361) );
  XNOR2_X1 U503 ( .A(n585), .B(n490), .ZN(n415) );
  XNOR2_X2 U504 ( .A(n412), .B(n411), .ZN(n618) );
  INV_X1 U505 ( .A(KEYINPUT2), .ZN(n364) );
  NAND2_X1 U506 ( .A1(n727), .A2(n738), .ZN(n365) );
  XNOR2_X1 U507 ( .A(n366), .B(KEYINPUT123), .ZN(G66) );
  NAND2_X1 U508 ( .A1(n389), .A2(n388), .ZN(n366) );
  INV_X1 U509 ( .A(n601), .ZN(n435) );
  NAND2_X1 U510 ( .A1(n406), .A2(n405), .ZN(n412) );
  NAND2_X1 U511 ( .A1(n618), .A2(n364), .ZN(n652) );
  XNOR2_X1 U512 ( .A(n422), .B(KEYINPUT107), .ZN(n413) );
  XNOR2_X1 U513 ( .A(n458), .B(n401), .ZN(n459) );
  NAND2_X1 U514 ( .A1(n700), .A2(n506), .ZN(n421) );
  XNOR2_X2 U515 ( .A(n374), .B(KEYINPUT83), .ZN(n559) );
  XNOR2_X1 U516 ( .A(n622), .B(n623), .ZN(n375) );
  XNOR2_X1 U517 ( .A(n420), .B(n524), .ZN(n376) );
  NOR2_X2 U518 ( .A1(n375), .A2(n719), .ZN(n626) );
  NAND2_X1 U519 ( .A1(n573), .A2(n664), .ZN(n581) );
  NOR2_X1 U520 ( .A1(n648), .A2(n640), .ZN(n377) );
  XNOR2_X1 U521 ( .A(n443), .B(n732), .ZN(n381) );
  INV_X1 U522 ( .A(n637), .ZN(n642) );
  NAND2_X1 U523 ( .A1(n637), .A2(KEYINPUT47), .ZN(n595) );
  NAND2_X1 U524 ( .A1(n436), .A2(n360), .ZN(n380) );
  XOR2_X2 U525 ( .A(G116), .B(G107), .Z(n481) );
  NAND2_X1 U526 ( .A1(n359), .A2(n407), .ZN(n405) );
  XNOR2_X1 U527 ( .A(n381), .B(n452), .ZN(n620) );
  NOR2_X2 U528 ( .A1(n531), .A2(n590), .ZN(n533) );
  XNOR2_X1 U529 ( .A(n384), .B(n383), .ZN(G51) );
  NAND2_X1 U530 ( .A1(n703), .A2(n388), .ZN(n384) );
  XNOR2_X1 U531 ( .A(n386), .B(n698), .ZN(G75) );
  BUF_X2 U532 ( .A(n669), .Z(n387) );
  XNOR2_X1 U533 ( .A(n619), .B(n390), .ZN(n389) );
  INV_X1 U534 ( .A(n620), .ZN(n390) );
  XNOR2_X1 U535 ( .A(n481), .B(n483), .ZN(n420) );
  NOR2_X2 U536 ( .A1(n555), .A2(n556), .ZN(n544) );
  NOR2_X1 U537 ( .A1(n434), .A2(n391), .ZN(n440) );
  NOR2_X1 U538 ( .A1(n620), .A2(G902), .ZN(n512) );
  XNOR2_X1 U539 ( .A(n392), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X2 U540 ( .A1(n714), .A2(n719), .ZN(n392) );
  XNOR2_X1 U541 ( .A(n444), .B(KEYINPUT94), .ZN(n393) );
  XNOR2_X1 U542 ( .A(n461), .B(n462), .ZN(n711) );
  XNOR2_X2 U543 ( .A(n404), .B(G131), .ZN(n493) );
  XNOR2_X2 U544 ( .A(G128), .B(G143), .ZN(n487) );
  NAND2_X1 U545 ( .A1(n415), .A2(n491), .ZN(n429) );
  NAND2_X1 U546 ( .A1(n593), .A2(n415), .ZN(n594) );
  NAND2_X1 U547 ( .A1(n632), .A2(n646), .ZN(n548) );
  NAND2_X1 U548 ( .A1(n439), .A2(n438), .ZN(n437) );
  NOR2_X1 U549 ( .A1(n574), .A2(n581), .ZN(n575) );
  NOR2_X1 U550 ( .A1(n435), .A2(KEYINPUT48), .ZN(n434) );
  NAND2_X1 U551 ( .A1(n588), .A2(n675), .ZN(n585) );
  XNOR2_X2 U552 ( .A(n421), .B(n357), .ZN(n588) );
  NAND2_X1 U553 ( .A1(n423), .A2(n628), .ZN(n422) );
  NAND2_X1 U554 ( .A1(n554), .A2(n591), .ZN(n423) );
  XNOR2_X2 U555 ( .A(n429), .B(n428), .ZN(n547) );
  XNOR2_X2 U556 ( .A(n430), .B(G472), .ZN(n669) );
  XNOR2_X1 U557 ( .A(n431), .B(n569), .ZN(n611) );
  NAND2_X1 U558 ( .A1(n587), .A2(n676), .ZN(n431) );
  INV_X1 U559 ( .A(n577), .ZN(n433) );
  AND2_X1 U560 ( .A1(n436), .A2(n614), .ZN(n738) );
  NAND2_X1 U561 ( .A1(n440), .A2(n437), .ZN(n436) );
  INV_X1 U562 ( .A(n602), .ZN(n439) );
  XNOR2_X1 U563 ( .A(n702), .B(n701), .ZN(n703) );
  XNOR2_X1 U564 ( .A(n580), .B(n579), .ZN(n602) );
  XNOR2_X1 U565 ( .A(n700), .B(n699), .ZN(n701) );
  XNOR2_X2 U566 ( .A(n480), .B(n479), .ZN(n524) );
  AND2_X1 U567 ( .A1(G221), .A2(n468), .ZN(n443) );
  INV_X1 U568 ( .A(KEYINPUT69), .ZN(n599) );
  XNOR2_X1 U569 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U570 ( .A(n522), .B(n521), .ZN(n523) );
  INV_X1 U571 ( .A(n502), .ZN(n503) );
  INV_X1 U572 ( .A(KEYINPUT25), .ZN(n509) );
  INV_X1 U573 ( .A(n651), .ZN(n613) );
  XNOR2_X1 U574 ( .A(n510), .B(n509), .ZN(n511) );
  NOR2_X1 U575 ( .A1(n613), .A2(n650), .ZN(n614) );
  INV_X1 U576 ( .A(KEYINPUT104), .ZN(n550) );
  XNOR2_X1 U577 ( .A(n467), .B(n466), .ZN(n470) );
  INV_X1 U578 ( .A(KEYINPUT105), .ZN(n552) );
  INV_X1 U579 ( .A(KEYINPUT63), .ZN(n624) );
  XNOR2_X1 U580 ( .A(n713), .B(n712), .ZN(n714) );
  XNOR2_X1 U581 ( .A(n624), .B(KEYINPUT84), .ZN(n625) );
  XOR2_X1 U582 ( .A(KEYINPUT23), .B(G128), .Z(n445) );
  XOR2_X1 U583 ( .A(KEYINPUT24), .B(KEYINPUT92), .Z(n447) );
  XNOR2_X1 U584 ( .A(KEYINPUT91), .B(KEYINPUT93), .ZN(n446) );
  XNOR2_X1 U585 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U586 ( .A(n448), .B(KEYINPUT75), .ZN(n449) );
  XNOR2_X1 U587 ( .A(n356), .B(n449), .ZN(n452) );
  NAND2_X1 U588 ( .A1(G234), .A2(n370), .ZN(n450) );
  XNOR2_X1 U589 ( .A(n451), .B(n450), .ZN(n468) );
  XNOR2_X1 U590 ( .A(n458), .B(n495), .ZN(n732) );
  XNOR2_X1 U591 ( .A(n454), .B(n493), .ZN(n462) );
  NAND2_X1 U592 ( .A1(n516), .A2(G214), .ZN(n455) );
  XNOR2_X1 U593 ( .A(n456), .B(n455), .ZN(n457) );
  XOR2_X1 U594 ( .A(n457), .B(KEYINPUT11), .Z(n460) );
  XNOR2_X1 U595 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U596 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U597 ( .A(n465), .B(n442), .ZN(n467) );
  XNOR2_X1 U598 ( .A(n487), .B(n481), .ZN(n466) );
  NAND2_X1 U599 ( .A1(G217), .A2(n468), .ZN(n469) );
  XNOR2_X1 U600 ( .A(n470), .B(n469), .ZN(n717) );
  NOR2_X1 U601 ( .A1(G902), .A2(n717), .ZN(n471) );
  INV_X1 U602 ( .A(n553), .ZN(n472) );
  NAND2_X1 U603 ( .A1(n549), .A2(n472), .ZN(n590) );
  XNOR2_X1 U604 ( .A(n473), .B(KEYINPUT14), .ZN(n475) );
  NAND2_X1 U605 ( .A1(G952), .A2(n475), .ZN(n690) );
  NOR2_X1 U606 ( .A1(G953), .A2(n690), .ZN(n567) );
  NOR2_X1 U607 ( .A1(G898), .A2(n370), .ZN(n474) );
  XOR2_X1 U608 ( .A(KEYINPUT88), .B(n474), .Z(n720) );
  NAND2_X1 U609 ( .A1(G902), .A2(n475), .ZN(n562) );
  NOR2_X1 U610 ( .A1(n720), .A2(n562), .ZN(n476) );
  NOR2_X1 U611 ( .A1(n567), .A2(n476), .ZN(n477) );
  XNOR2_X1 U612 ( .A(n477), .B(KEYINPUT89), .ZN(n491) );
  XNOR2_X1 U613 ( .A(KEYINPUT74), .B(KEYINPUT19), .ZN(n490) );
  XNOR2_X1 U614 ( .A(n478), .B(KEYINPUT71), .ZN(n489) );
  XOR2_X1 U615 ( .A(G110), .B(KEYINPUT86), .Z(n502) );
  XOR2_X1 U616 ( .A(KEYINPUT16), .B(n502), .Z(n482) );
  NAND2_X1 U617 ( .A1(G224), .A2(n370), .ZN(n485) );
  INV_X1 U618 ( .A(n617), .ZN(n506) );
  NAND2_X1 U619 ( .A1(G214), .A2(n489), .ZN(n675) );
  XNOR2_X1 U620 ( .A(n547), .B(n492), .ZN(n545) );
  INV_X1 U621 ( .A(n525), .ZN(n499) );
  INV_X1 U622 ( .A(n495), .ZN(n496) );
  XOR2_X1 U623 ( .A(n496), .B(G104), .Z(n497) );
  NAND2_X1 U624 ( .A1(G227), .A2(n370), .ZN(n501) );
  NAND2_X1 U625 ( .A1(G234), .A2(n506), .ZN(n507) );
  XNOR2_X1 U626 ( .A(n508), .B(n507), .ZN(n513) );
  NAND2_X1 U627 ( .A1(G217), .A2(n513), .ZN(n510) );
  NAND2_X1 U628 ( .A1(n513), .A2(G221), .ZN(n514) );
  XNOR2_X1 U629 ( .A(n514), .B(KEYINPUT21), .ZN(n663) );
  XNOR2_X1 U630 ( .A(n663), .B(KEYINPUT96), .ZN(n536) );
  XOR2_X1 U631 ( .A(KEYINPUT97), .B(KEYINPUT5), .Z(n518) );
  NAND2_X1 U632 ( .A1(G210), .A2(n516), .ZN(n517) );
  XNOR2_X1 U633 ( .A(n518), .B(n517), .ZN(n522) );
  XNOR2_X1 U634 ( .A(G137), .B(G116), .ZN(n520) );
  XNOR2_X1 U635 ( .A(n524), .B(n523), .ZN(n526) );
  XNOR2_X1 U636 ( .A(n669), .B(KEYINPUT6), .ZN(n582) );
  OR2_X1 U637 ( .A1(n659), .A2(n582), .ZN(n527) );
  XNOR2_X1 U638 ( .A(n528), .B(KEYINPUT33), .ZN(n691) );
  NOR2_X1 U639 ( .A1(n545), .A2(n691), .ZN(n530) );
  INV_X1 U640 ( .A(KEYINPUT34), .ZN(n529) );
  XNOR2_X1 U641 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X2 U642 ( .A(n533), .B(n532), .ZN(n743) );
  INV_X1 U643 ( .A(n549), .ZN(n535) );
  NAND2_X1 U644 ( .A1(n535), .A2(n553), .ZN(n679) );
  NOR2_X1 U645 ( .A1(n536), .A2(n679), .ZN(n537) );
  XNOR2_X1 U646 ( .A(KEYINPUT106), .B(n537), .ZN(n538) );
  NAND2_X1 U647 ( .A1(n538), .A2(n547), .ZN(n539) );
  INV_X1 U648 ( .A(n664), .ZN(n556) );
  XOR2_X1 U649 ( .A(KEYINPUT76), .B(n582), .Z(n540) );
  NOR2_X1 U650 ( .A1(n660), .A2(n540), .ZN(n541) );
  NAND2_X1 U651 ( .A1(n544), .A2(n541), .ZN(n542) );
  INV_X1 U652 ( .A(n660), .ZN(n606) );
  NOR2_X1 U653 ( .A1(n387), .A2(n606), .ZN(n543) );
  NAND2_X1 U654 ( .A1(n544), .A2(n543), .ZN(n636) );
  NOR2_X1 U655 ( .A1(n387), .A2(n577), .ZN(n546) );
  XNOR2_X1 U656 ( .A(n548), .B(KEYINPUT100), .ZN(n554) );
  XNOR2_X2 U657 ( .A(n551), .B(n550), .ZN(n631) );
  NAND2_X1 U658 ( .A1(n549), .A2(n553), .ZN(n644) );
  NAND2_X1 U659 ( .A1(n612), .A2(n644), .ZN(n591) );
  NOR2_X1 U660 ( .A1(n555), .A2(n606), .ZN(n558) );
  AND2_X1 U661 ( .A1(n556), .A2(n582), .ZN(n557) );
  NAND2_X1 U662 ( .A1(n558), .A2(n557), .ZN(n628) );
  XOR2_X1 U663 ( .A(KEYINPUT30), .B(KEYINPUT112), .Z(n561) );
  NAND2_X1 U664 ( .A1(n669), .A2(n675), .ZN(n560) );
  XNOR2_X1 U665 ( .A(n561), .B(n560), .ZN(n568) );
  OR2_X1 U666 ( .A1(n370), .A2(n562), .ZN(n563) );
  XNOR2_X1 U667 ( .A(KEYINPUT108), .B(n563), .ZN(n564) );
  NOR2_X1 U668 ( .A1(G900), .A2(n564), .ZN(n565) );
  XOR2_X1 U669 ( .A(KEYINPUT109), .B(n565), .Z(n566) );
  NOR2_X1 U670 ( .A1(n567), .A2(n566), .ZN(n572) );
  INV_X1 U671 ( .A(n588), .ZN(n609) );
  XOR2_X1 U672 ( .A(KEYINPUT82), .B(KEYINPUT39), .Z(n569) );
  NOR2_X1 U673 ( .A1(n611), .A2(n644), .ZN(n570) );
  NAND2_X1 U674 ( .A1(n676), .A2(n675), .ZN(n682) );
  XOR2_X1 U675 ( .A(KEYINPUT41), .B(n571), .Z(n658) );
  INV_X1 U676 ( .A(n387), .ZN(n574) );
  NOR2_X1 U677 ( .A1(n663), .A2(n572), .ZN(n573) );
  XOR2_X1 U678 ( .A(KEYINPUT28), .B(n575), .Z(n576) );
  NOR2_X1 U679 ( .A1(n577), .A2(n576), .ZN(n593) );
  NAND2_X1 U680 ( .A1(n658), .A2(n593), .ZN(n578) );
  NOR2_X1 U681 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U682 ( .A(KEYINPUT110), .B(n583), .ZN(n584) );
  INV_X1 U683 ( .A(n644), .ZN(n641) );
  NAND2_X1 U684 ( .A1(n584), .A2(n641), .ZN(n603) );
  NOR2_X1 U685 ( .A1(n660), .A2(n586), .ZN(n648) );
  NAND2_X1 U686 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U687 ( .A1(n590), .A2(n589), .ZN(n640) );
  NAND2_X1 U688 ( .A1(n681), .A2(KEYINPUT47), .ZN(n592) );
  XNOR2_X1 U689 ( .A(n592), .B(KEYINPUT78), .ZN(n596) );
  NOR2_X1 U690 ( .A1(n681), .A2(KEYINPUT47), .ZN(n597) );
  XNOR2_X1 U691 ( .A(KEYINPUT70), .B(n597), .ZN(n598) );
  NAND2_X1 U692 ( .A1(n598), .A2(n642), .ZN(n600) );
  INV_X1 U693 ( .A(n603), .ZN(n604) );
  NAND2_X1 U694 ( .A1(n604), .A2(n675), .ZN(n605) );
  NOR2_X1 U695 ( .A1(n606), .A2(n605), .ZN(n608) );
  XNOR2_X1 U696 ( .A(KEYINPUT43), .B(KEYINPUT111), .ZN(n607) );
  XNOR2_X1 U697 ( .A(n608), .B(n607), .ZN(n610) );
  NAND2_X1 U698 ( .A1(n610), .A2(n609), .ZN(n651) );
  NOR2_X1 U699 ( .A1(n612), .A2(n611), .ZN(n650) );
  NAND2_X1 U700 ( .A1(G217), .A2(n715), .ZN(n619) );
  NAND2_X1 U701 ( .A1(G472), .A2(n715), .ZN(n622) );
  XNOR2_X1 U702 ( .A(n626), .B(n625), .ZN(G57) );
  XOR2_X1 U703 ( .A(G101), .B(KEYINPUT113), .Z(n627) );
  XNOR2_X1 U704 ( .A(n628), .B(n627), .ZN(G3) );
  NOR2_X1 U705 ( .A1(n632), .A2(n644), .ZN(n629) );
  XOR2_X1 U706 ( .A(KEYINPUT114), .B(n629), .Z(n630) );
  XNOR2_X1 U707 ( .A(G104), .B(n630), .ZN(G6) );
  XNOR2_X1 U708 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n634) );
  NOR2_X1 U709 ( .A1(n631), .A2(n632), .ZN(n633) );
  XNOR2_X1 U710 ( .A(n634), .B(n633), .ZN(n635) );
  XNOR2_X1 U711 ( .A(G107), .B(n635), .ZN(G9) );
  XNOR2_X1 U712 ( .A(G110), .B(n636), .ZN(G12) );
  XOR2_X1 U713 ( .A(G128), .B(KEYINPUT29), .Z(n639) );
  OR2_X1 U714 ( .A1(n637), .A2(n631), .ZN(n638) );
  XNOR2_X1 U715 ( .A(n639), .B(n638), .ZN(G30) );
  XOR2_X1 U716 ( .A(G143), .B(n640), .Z(G45) );
  NAND2_X1 U717 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U718 ( .A(n643), .B(G146), .ZN(G48) );
  NOR2_X1 U719 ( .A1(n644), .A2(n646), .ZN(n645) );
  XOR2_X1 U720 ( .A(G113), .B(n645), .Z(G15) );
  NOR2_X1 U721 ( .A1(n631), .A2(n646), .ZN(n647) );
  XOR2_X1 U722 ( .A(G116), .B(n647), .Z(G18) );
  XNOR2_X1 U723 ( .A(G125), .B(n648), .ZN(n649) );
  XNOR2_X1 U724 ( .A(n649), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U725 ( .A(G134), .B(n650), .Z(G36) );
  XNOR2_X1 U726 ( .A(G140), .B(n651), .ZN(G42) );
  XNOR2_X1 U727 ( .A(n652), .B(KEYINPUT79), .ZN(n654) );
  NOR2_X1 U728 ( .A1(n738), .A2(KEYINPUT2), .ZN(n653) );
  NOR2_X1 U729 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U730 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U731 ( .A(n657), .B(KEYINPUT80), .ZN(n697) );
  INV_X1 U732 ( .A(n658), .ZN(n692) );
  AND2_X1 U733 ( .A1(n387), .A2(n355), .ZN(n671) );
  XOR2_X1 U734 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n662) );
  NAND2_X1 U735 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U736 ( .A(n662), .B(n661), .ZN(n667) );
  NAND2_X1 U737 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U738 ( .A(KEYINPUT49), .B(n665), .Z(n666) );
  NAND2_X1 U739 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U740 ( .A1(n387), .A2(n668), .ZN(n670) );
  NOR2_X1 U741 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U742 ( .A(n672), .B(KEYINPUT51), .Z(n673) );
  XNOR2_X1 U743 ( .A(KEYINPUT116), .B(n673), .ZN(n674) );
  NOR2_X1 U744 ( .A1(n692), .A2(n674), .ZN(n687) );
  NOR2_X1 U745 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U746 ( .A(KEYINPUT117), .B(n677), .Z(n678) );
  NOR2_X1 U747 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U748 ( .A(n680), .B(KEYINPUT118), .ZN(n684) );
  NOR2_X1 U749 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U750 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U751 ( .A1(n685), .A2(n691), .ZN(n686) );
  NOR2_X1 U752 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U753 ( .A(n688), .B(KEYINPUT52), .ZN(n689) );
  NOR2_X1 U754 ( .A1(n690), .A2(n689), .ZN(n695) );
  NOR2_X1 U755 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U756 ( .A(KEYINPUT119), .B(n693), .Z(n694) );
  NOR2_X1 U757 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U758 ( .A(KEYINPUT53), .B(KEYINPUT120), .ZN(n698) );
  NAND2_X1 U759 ( .A1(n715), .A2(G210), .ZN(n702) );
  XOR2_X1 U760 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n699) );
  XOR2_X1 U761 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n706) );
  XNOR2_X1 U762 ( .A(n704), .B(KEYINPUT121), .ZN(n705) );
  XNOR2_X1 U763 ( .A(n706), .B(n705), .ZN(n708) );
  NAND2_X1 U764 ( .A1(n715), .A2(G469), .ZN(n707) );
  XOR2_X1 U765 ( .A(n708), .B(n707), .Z(n709) );
  NOR2_X1 U766 ( .A1(n719), .A2(n709), .ZN(G54) );
  NAND2_X1 U767 ( .A1(n715), .A2(G475), .ZN(n713) );
  INV_X1 U768 ( .A(KEYINPUT59), .ZN(n710) );
  NAND2_X1 U769 ( .A1(n715), .A2(G478), .ZN(n716) );
  NOR2_X1 U770 ( .A1(n719), .A2(n718), .ZN(G63) );
  INV_X1 U771 ( .A(n720), .ZN(n722) );
  NOR2_X1 U772 ( .A1(n722), .A2(n721), .ZN(n731) );
  XOR2_X1 U773 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n724) );
  NAND2_X1 U774 ( .A1(G224), .A2(G953), .ZN(n723) );
  XNOR2_X1 U775 ( .A(n724), .B(n723), .ZN(n725) );
  XNOR2_X1 U776 ( .A(KEYINPUT124), .B(n725), .ZN(n726) );
  NAND2_X1 U777 ( .A1(G898), .A2(n726), .ZN(n729) );
  NAND2_X1 U778 ( .A1(n727), .A2(n370), .ZN(n728) );
  NAND2_X1 U779 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U780 ( .A(n731), .B(n730), .ZN(G69) );
  XOR2_X1 U781 ( .A(n733), .B(n732), .Z(n734) );
  XNOR2_X1 U782 ( .A(KEYINPUT126), .B(n734), .ZN(n739) );
  XNOR2_X1 U783 ( .A(KEYINPUT127), .B(n739), .ZN(n735) );
  XNOR2_X1 U784 ( .A(G227), .B(n735), .ZN(n736) );
  NAND2_X1 U785 ( .A1(n736), .A2(G900), .ZN(n737) );
  NAND2_X1 U786 ( .A1(n737), .A2(G953), .ZN(n742) );
  XNOR2_X1 U787 ( .A(n739), .B(n738), .ZN(n740) );
  NAND2_X1 U788 ( .A1(n740), .A2(n370), .ZN(n741) );
  NAND2_X1 U789 ( .A1(n742), .A2(n741), .ZN(G72) );
  XOR2_X1 U790 ( .A(G122), .B(n743), .Z(G24) );
  XNOR2_X1 U791 ( .A(n744), .B(G119), .ZN(G21) );
  XNOR2_X1 U792 ( .A(G131), .B(n745), .ZN(G33) );
  XNOR2_X1 U793 ( .A(G137), .B(n746), .ZN(G39) );
endmodule

