

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759;

  AND2_X2 U361 ( .A1(n476), .A2(n477), .ZN(n358) );
  NAND2_X1 U362 ( .A1(n645), .A2(n646), .ZN(n740) );
  XNOR2_X1 U363 ( .A(n481), .B(n340), .ZN(n361) );
  INV_X1 U364 ( .A(KEYINPUT44), .ZN(n340) );
  XNOR2_X1 U365 ( .A(n486), .B(G119), .ZN(n378) );
  XNOR2_X1 U366 ( .A(G116), .B(G113), .ZN(n377) );
  XNOR2_X2 U367 ( .A(n538), .B(n339), .ZN(n734) );
  XNOR2_X2 U368 ( .A(n419), .B(n484), .ZN(n339) );
  NAND2_X1 U369 ( .A1(n633), .A2(n346), .ZN(n479) );
  XNOR2_X2 U370 ( .A(n615), .B(n480), .ZN(n633) );
  NAND2_X2 U371 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X2 U372 ( .A1(n716), .A2(n548), .ZN(n550) );
  XNOR2_X2 U373 ( .A(n561), .B(n501), .ZN(n545) );
  XNOR2_X2 U374 ( .A(n500), .B(n499), .ZN(n561) );
  XNOR2_X1 U375 ( .A(n545), .B(n494), .ZN(n746) );
  NAND2_X1 U376 ( .A1(n421), .A2(n420), .ZN(n472) );
  AND2_X1 U377 ( .A1(n424), .A2(n422), .ZN(n421) );
  NAND2_X1 U378 ( .A1(n740), .A2(n465), .ZN(n402) );
  XNOR2_X1 U379 ( .A(n385), .B(n466), .ZN(n465) );
  AND2_X1 U380 ( .A1(n384), .A2(n607), .ZN(n747) );
  NOR2_X1 U381 ( .A1(n757), .A2(n759), .ZN(n578) );
  XNOR2_X1 U382 ( .A(n362), .B(n354), .ZN(n756) );
  NOR2_X1 U383 ( .A1(n637), .A2(n700), .ZN(n622) );
  NOR2_X1 U384 ( .A1(n630), .A2(n713), .ZN(n618) );
  OR2_X1 U385 ( .A1(n456), .A2(n592), .ZN(n594) );
  NAND2_X1 U386 ( .A1(n431), .A2(n429), .ZN(n688) );
  NOR2_X1 U387 ( .A1(n587), .A2(n400), .ZN(n667) );
  XNOR2_X1 U388 ( .A(n475), .B(n586), .ZN(n608) );
  XNOR2_X1 U389 ( .A(n524), .B(n523), .ZN(n697) );
  INV_X1 U390 ( .A(n498), .ZN(n500) );
  XNOR2_X1 U391 ( .A(KEYINPUT81), .B(KEYINPUT66), .ZN(n499) );
  XNOR2_X1 U392 ( .A(G128), .B(G143), .ZN(n498) );
  INV_X1 U393 ( .A(n681), .ZN(n476) );
  XNOR2_X1 U394 ( .A(n402), .B(n649), .ZN(n681) );
  XOR2_X1 U395 ( .A(KEYINPUT92), .B(n528), .Z(n684) );
  INV_X1 U396 ( .A(KEYINPUT10), .ZN(n462) );
  XNOR2_X1 U397 ( .A(n467), .B(KEYINPUT72), .ZN(n568) );
  XNOR2_X1 U398 ( .A(G131), .B(G146), .ZN(n467) );
  XNOR2_X1 U399 ( .A(KEYINPUT4), .B(KEYINPUT65), .ZN(n501) );
  OR2_X1 U400 ( .A1(n678), .A2(n606), .ZN(n367) );
  XNOR2_X1 U401 ( .A(n365), .B(n457), .ZN(n384) );
  INV_X1 U402 ( .A(KEYINPUT48), .ZN(n457) );
  AND2_X1 U403 ( .A1(n676), .A2(n597), .ZN(n598) );
  AND2_X1 U404 ( .A1(n437), .A2(n435), .ZN(n432) );
  INV_X1 U405 ( .A(KEYINPUT42), .ZN(n396) );
  NOR2_X1 U406 ( .A1(n697), .A2(n573), .ZN(n579) );
  NAND2_X1 U407 ( .A1(n697), .A2(n696), .ZN(n693) );
  OR2_X1 U408 ( .A1(n722), .A2(G902), .ZN(n418) );
  XNOR2_X1 U409 ( .A(n513), .B(n453), .ZN(n557) );
  INV_X1 U410 ( .A(KEYINPUT8), .ZN(n453) );
  NOR2_X1 U411 ( .A1(n342), .A2(n715), .ZN(n492) );
  NAND2_X1 U412 ( .A1(n413), .A2(n410), .ZN(n605) );
  NAND2_X1 U413 ( .A1(n412), .A2(n411), .ZN(n410) );
  AND2_X1 U414 ( .A1(n415), .A2(n414), .ZN(n413) );
  XNOR2_X1 U415 ( .A(n571), .B(KEYINPUT106), .ZN(n589) );
  NOR2_X1 U416 ( .A1(n595), .A2(n666), .ZN(n596) );
  XNOR2_X1 U417 ( .A(KEYINPUT41), .B(KEYINPUT117), .ZN(n577) );
  NOR2_X1 U418 ( .A1(G953), .A2(G237), .ZN(n564) );
  XNOR2_X1 U419 ( .A(G101), .B(KEYINPUT100), .ZN(n502) );
  XNOR2_X1 U420 ( .A(n373), .B(n371), .ZN(n370) );
  XNOR2_X1 U421 ( .A(n567), .B(n372), .ZN(n371) );
  XNOR2_X1 U422 ( .A(n565), .B(n562), .ZN(n373) );
  INV_X1 U423 ( .A(KEYINPUT11), .ZN(n372) );
  XNOR2_X1 U424 ( .A(n566), .B(n563), .ZN(n369) );
  XOR2_X1 U425 ( .A(KEYINPUT103), .B(KEYINPUT101), .Z(n563) );
  NOR2_X1 U426 ( .A1(n756), .A2(n482), .ZN(n364) );
  NOR2_X1 U427 ( .A1(n367), .A2(n506), .ZN(n383) );
  INV_X1 U428 ( .A(n587), .ZN(n394) );
  NAND2_X1 U429 ( .A1(n430), .A2(n341), .ZN(n429) );
  AND2_X1 U430 ( .A1(n439), .A2(n438), .ZN(n431) );
  INV_X1 U431 ( .A(n599), .ZN(n593) );
  XNOR2_X1 U432 ( .A(n522), .B(KEYINPUT25), .ZN(n523) );
  NOR2_X1 U433 ( .A1(G902), .A2(n731), .ZN(n524) );
  XNOR2_X1 U434 ( .A(n582), .B(n581), .ZN(n694) );
  INV_X1 U435 ( .A(KEYINPUT1), .ZN(n581) );
  XNOR2_X1 U436 ( .A(n518), .B(n516), .ZN(n460) );
  XNOR2_X1 U437 ( .A(KEYINPUT23), .B(KEYINPUT73), .ZN(n518) );
  XNOR2_X1 U438 ( .A(n745), .B(n464), .ZN(n461) );
  XNOR2_X1 U439 ( .A(n514), .B(n517), .ZN(n464) );
  XNOR2_X1 U440 ( .A(G128), .B(G119), .ZN(n517) );
  AND2_X1 U441 ( .A1(n740), .A2(n548), .ZN(n455) );
  XNOR2_X1 U442 ( .A(n374), .B(n507), .ZN(n538) );
  XNOR2_X1 U443 ( .A(G104), .B(n375), .ZN(n374) );
  XNOR2_X1 U444 ( .A(KEYINPUT90), .B(G101), .ZN(n375) );
  XNOR2_X1 U445 ( .A(n568), .B(n347), .ZN(n494) );
  NOR2_X1 U446 ( .A1(n427), .A2(n426), .ZN(n425) );
  INV_X1 U447 ( .A(KEYINPUT121), .ZN(n426) );
  XNOR2_X1 U448 ( .A(n600), .B(KEYINPUT110), .ZN(n601) );
  NOR2_X1 U449 ( .A1(n587), .A2(n396), .ZN(n391) );
  NAND2_X1 U450 ( .A1(n668), .A2(n469), .ZN(n600) );
  NOR2_X1 U451 ( .A1(n616), .A2(n470), .ZN(n469) );
  NAND2_X1 U452 ( .A1(n579), .A2(n584), .ZN(n470) );
  NOR2_X1 U453 ( .A1(n489), .A2(n488), .ZN(n487) );
  INV_X1 U454 ( .A(n572), .ZN(n488) );
  BUF_X1 U455 ( .A(n593), .Z(n456) );
  XNOR2_X1 U456 ( .A(n585), .B(KEYINPUT70), .ZN(n586) );
  INV_X1 U457 ( .A(KEYINPUT19), .ZN(n585) );
  XNOR2_X1 U458 ( .A(n570), .B(n569), .ZN(n366) );
  NOR2_X1 U459 ( .A1(G902), .A2(n726), .ZN(n570) );
  BUF_X1 U460 ( .A(n697), .Z(n448) );
  INV_X1 U461 ( .A(n616), .ZN(n636) );
  INV_X1 U462 ( .A(KEYINPUT64), .ZN(n454) );
  XNOR2_X1 U463 ( .A(n382), .B(n355), .ZN(n381) );
  XNOR2_X1 U464 ( .A(G122), .B(G113), .ZN(n562) );
  XNOR2_X1 U465 ( .A(G143), .B(G104), .ZN(n567) );
  NAND2_X1 U466 ( .A1(n684), .A2(KEYINPUT116), .ZN(n438) );
  XOR2_X1 U467 ( .A(KEYINPUT97), .B(KEYINPUT20), .Z(n510) );
  XOR2_X1 U468 ( .A(KEYINPUT91), .B(KEYINPUT17), .Z(n543) );
  INV_X1 U469 ( .A(KEYINPUT18), .ZN(n539) );
  XNOR2_X1 U470 ( .A(G125), .B(G146), .ZN(n540) );
  INV_X1 U471 ( .A(KEYINPUT86), .ZN(n466) );
  OR2_X1 U472 ( .A1(G902), .A2(G237), .ZN(n549) );
  NAND2_X1 U473 ( .A1(n436), .A2(n434), .ZN(n397) );
  OR2_X1 U474 ( .A1(n437), .A2(n435), .ZN(n434) );
  INV_X1 U475 ( .A(KEYINPUT38), .ZN(n450) );
  XNOR2_X1 U476 ( .A(n617), .B(n440), .ZN(n713) );
  INV_X1 U477 ( .A(KEYINPUT33), .ZN(n440) );
  NAND2_X1 U478 ( .A1(n636), .A2(n629), .ZN(n617) );
  XNOR2_X1 U479 ( .A(n529), .B(n490), .ZN(n489) );
  XNOR2_X1 U480 ( .A(n530), .B(KEYINPUT113), .ZN(n490) );
  NAND2_X1 U481 ( .A1(n700), .A2(n584), .ZN(n529) );
  XNOR2_X1 U482 ( .A(n700), .B(KEYINPUT6), .ZN(n616) );
  XNOR2_X1 U483 ( .A(n746), .B(n493), .ZN(n525) );
  XNOR2_X1 U484 ( .A(KEYINPUT104), .B(KEYINPUT9), .ZN(n553) );
  XOR2_X1 U485 ( .A(G134), .B(KEYINPUT7), .Z(n554) );
  XNOR2_X1 U486 ( .A(G107), .B(G122), .ZN(n551) );
  XOR2_X1 U487 ( .A(KEYINPUT105), .B(G116), .Z(n552) );
  XNOR2_X1 U488 ( .A(n473), .B(n368), .ZN(n726) );
  XNOR2_X1 U489 ( .A(n370), .B(n369), .ZN(n368) );
  INV_X1 U490 ( .A(n367), .ZN(n607) );
  AND2_X1 U491 ( .A1(n387), .A2(n396), .ZN(n386) );
  INV_X1 U492 ( .A(n432), .ZN(n388) );
  INV_X1 U493 ( .A(n397), .ZN(n399) );
  NAND2_X1 U494 ( .A1(n397), .A2(n396), .ZN(n395) );
  AND2_X1 U495 ( .A1(n700), .A2(n579), .ZN(n575) );
  XNOR2_X1 U496 ( .A(n401), .B(G478), .ZN(n588) );
  NOR2_X1 U497 ( .A1(n728), .A2(G902), .ZN(n401) );
  INV_X1 U498 ( .A(KEYINPUT99), .ZN(n444) );
  INV_X1 U499 ( .A(KEYINPUT0), .ZN(n480) );
  NAND2_X1 U500 ( .A1(n358), .A2(G472), .ZN(n650) );
  XNOR2_X1 U501 ( .A(n485), .B(G122), .ZN(n484) );
  INV_X1 U502 ( .A(KEYINPUT16), .ZN(n485) );
  XNOR2_X1 U503 ( .A(n519), .B(n520), .ZN(n731) );
  XNOR2_X1 U504 ( .A(n461), .B(n459), .ZN(n519) );
  XNOR2_X1 U505 ( .A(n515), .B(n460), .ZN(n459) );
  XNOR2_X1 U506 ( .A(n468), .B(n746), .ZN(n722) );
  XNOR2_X1 U507 ( .A(n449), .B(n538), .ZN(n468) );
  XNOR2_X1 U508 ( .A(n508), .B(G140), .ZN(n449) );
  NAND2_X1 U509 ( .A1(n358), .A2(G469), .ZN(n724) );
  NAND2_X1 U510 ( .A1(n358), .A2(G210), .ZN(n478) );
  NOR2_X1 U511 ( .A1(n423), .A2(G953), .ZN(n422) );
  NOR2_X1 U512 ( .A1(n492), .A2(KEYINPUT121), .ZN(n423) );
  NOR2_X1 U513 ( .A1(n604), .A2(n599), .ZN(n678) );
  NAND2_X1 U514 ( .A1(n392), .A2(n390), .ZN(n757) );
  AND2_X1 U515 ( .A1(n395), .A2(n393), .ZN(n392) );
  NAND2_X1 U516 ( .A1(n343), .A2(n399), .ZN(n390) );
  NAND2_X1 U517 ( .A1(n389), .A2(n386), .ZN(n393) );
  NAND2_X1 U518 ( .A1(n405), .A2(n403), .ZN(n759) );
  NAND2_X1 U519 ( .A1(n404), .A2(n349), .ZN(n403) );
  AND2_X1 U520 ( .A1(n406), .A2(n408), .ZN(n405) );
  NOR2_X1 U521 ( .A1(n600), .A2(n456), .ZN(n580) );
  INV_X1 U522 ( .A(n619), .ZN(n451) );
  XNOR2_X1 U523 ( .A(n628), .B(n360), .ZN(n482) );
  INV_X1 U524 ( .A(KEYINPUT32), .ZN(n360) );
  XNOR2_X1 U525 ( .A(n589), .B(KEYINPUT109), .ZN(n668) );
  BUF_X1 U526 ( .A(n608), .Z(n400) );
  INV_X1 U527 ( .A(n448), .ZN(n445) );
  INV_X1 U528 ( .A(KEYINPUT67), .ZN(n447) );
  INV_X1 U529 ( .A(n668), .ZN(n670) );
  INV_X1 U530 ( .A(n733), .ZN(n380) );
  XNOR2_X1 U531 ( .A(n482), .B(n359), .ZN(G21) );
  INV_X1 U532 ( .A(G119), .ZN(n359) );
  INV_X1 U533 ( .A(n589), .ZN(n409) );
  NOR2_X1 U534 ( .A1(n684), .A2(KEYINPUT116), .ZN(n341) );
  AND2_X1 U535 ( .A1(n712), .A2(n711), .ZN(n342) );
  AND2_X1 U536 ( .A1(n398), .A2(n391), .ZN(n343) );
  NAND2_X1 U537 ( .A1(G210), .A2(n549), .ZN(n344) );
  AND2_X1 U538 ( .A1(n640), .A2(n654), .ZN(n345) );
  XNOR2_X1 U539 ( .A(KEYINPUT107), .B(n621), .ZN(n346) );
  XOR2_X1 U540 ( .A(G137), .B(G134), .Z(n347) );
  AND2_X1 U541 ( .A1(n345), .A2(n642), .ZN(n348) );
  AND2_X1 U542 ( .A1(n409), .A2(n407), .ZN(n349) );
  XNOR2_X1 U543 ( .A(KEYINPUT115), .B(KEYINPUT40), .ZN(n350) );
  XOR2_X1 U544 ( .A(KEYINPUT39), .B(KEYINPUT74), .Z(n351) );
  XOR2_X1 U545 ( .A(n718), .B(n717), .Z(n352) );
  XOR2_X1 U546 ( .A(KEYINPUT22), .B(KEYINPUT68), .Z(n353) );
  XOR2_X1 U547 ( .A(KEYINPUT79), .B(KEYINPUT35), .Z(n354) );
  XOR2_X1 U548 ( .A(n726), .B(n497), .Z(n355) );
  OR2_X1 U549 ( .A1(n506), .A2(n505), .ZN(n356) );
  XNOR2_X1 U550 ( .A(G902), .B(KEYINPUT15), .ZN(n648) );
  XNOR2_X1 U551 ( .A(KEYINPUT71), .B(KEYINPUT60), .ZN(n357) );
  INV_X1 U552 ( .A(G953), .ZN(n739) );
  NAND2_X1 U553 ( .A1(n358), .A2(G475), .ZN(n382) );
  NAND2_X1 U554 ( .A1(n358), .A2(G478), .ZN(n727) );
  NAND2_X1 U555 ( .A1(n358), .A2(G217), .ZN(n730) );
  NAND2_X1 U556 ( .A1(n361), .A2(n345), .ZN(n644) );
  NAND2_X1 U557 ( .A1(n361), .A2(n348), .ZN(n646) );
  NAND2_X1 U558 ( .A1(n452), .A2(n451), .ZN(n362) );
  NAND2_X1 U559 ( .A1(n458), .A2(n598), .ZN(n365) );
  NAND2_X1 U560 ( .A1(n363), .A2(n356), .ZN(n477) );
  NAND2_X1 U561 ( .A1(n384), .A2(n383), .ZN(n385) );
  NAND2_X1 U562 ( .A1(n626), .A2(n694), .ZN(n637) );
  NAND2_X1 U563 ( .A1(n647), .A2(n455), .ZN(n363) );
  NAND2_X1 U564 ( .A1(n364), .A2(n483), .ZN(n481) );
  NAND2_X1 U565 ( .A1(n446), .A2(n445), .ZN(n483) );
  NAND2_X1 U566 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U567 ( .A1(n525), .A2(G902), .ZN(n527) );
  NAND2_X1 U568 ( .A1(n667), .A2(n687), .ZN(n590) );
  NAND2_X1 U569 ( .A1(n588), .A2(n366), .ZN(n571) );
  NOR2_X1 U570 ( .A1(n588), .A2(n366), .ZN(n663) );
  NOR2_X1 U571 ( .A1(n591), .A2(n366), .ZN(n620) );
  NAND2_X1 U572 ( .A1(n591), .A2(n366), .ZN(n619) );
  XNOR2_X2 U573 ( .A(n378), .B(n377), .ZN(n419) );
  XNOR2_X1 U574 ( .A(n379), .B(n357), .ZN(G60) );
  NAND2_X1 U575 ( .A1(n381), .A2(n380), .ZN(n379) );
  NAND2_X1 U576 ( .A1(n433), .A2(n432), .ZN(n398) );
  NAND2_X1 U577 ( .A1(n394), .A2(n388), .ZN(n387) );
  NAND2_X1 U578 ( .A1(n688), .A2(n394), .ZN(n389) );
  NAND2_X1 U579 ( .A1(n399), .A2(n398), .ZN(n714) );
  XNOR2_X1 U580 ( .A(n478), .B(n352), .ZN(n719) );
  XNOR2_X1 U581 ( .A(n650), .B(n651), .ZN(n652) );
  XNOR2_X1 U582 ( .A(n724), .B(n723), .ZN(n725) );
  INV_X1 U583 ( .A(n633), .ZN(n630) );
  INV_X1 U584 ( .A(n605), .ZN(n404) );
  NAND2_X1 U585 ( .A1(n605), .A2(n350), .ZN(n406) );
  INV_X1 U586 ( .A(n350), .ZN(n407) );
  NAND2_X1 U587 ( .A1(n589), .A2(n350), .ZN(n408) );
  NOR2_X1 U588 ( .A1(n683), .A2(n351), .ZN(n411) );
  INV_X1 U589 ( .A(n592), .ZN(n412) );
  NAND2_X1 U590 ( .A1(n683), .A2(n351), .ZN(n414) );
  NAND2_X1 U591 ( .A1(n592), .A2(n351), .ZN(n415) );
  XNOR2_X2 U592 ( .A(n416), .B(n444), .ZN(n632) );
  NAND2_X1 U593 ( .A1(n582), .A2(n417), .ZN(n416) );
  INV_X1 U594 ( .A(n693), .ZN(n417) );
  XNOR2_X2 U595 ( .A(n418), .B(G469), .ZN(n582) );
  XNOR2_X1 U596 ( .A(n419), .B(n504), .ZN(n493) );
  OR2_X1 U597 ( .A1(n428), .A2(KEYINPUT121), .ZN(n420) );
  NAND2_X1 U598 ( .A1(n428), .A2(n425), .ZN(n424) );
  INV_X1 U599 ( .A(n492), .ZN(n427) );
  XNOR2_X1 U600 ( .A(n682), .B(KEYINPUT83), .ZN(n428) );
  NAND2_X1 U601 ( .A1(n688), .A2(n577), .ZN(n436) );
  INV_X1 U602 ( .A(n683), .ZN(n430) );
  INV_X1 U603 ( .A(n688), .ZN(n433) );
  INV_X1 U604 ( .A(n577), .ZN(n435) );
  INV_X1 U605 ( .A(n686), .ZN(n437) );
  NAND2_X1 U606 ( .A1(n683), .A2(KEYINPUT116), .ZN(n439) );
  NOR2_X2 U607 ( .A1(n652), .A2(n733), .ZN(n443) );
  NAND2_X1 U608 ( .A1(n626), .A2(n627), .ZN(n628) );
  XNOR2_X2 U609 ( .A(n479), .B(n353), .ZN(n626) );
  INV_X2 U610 ( .A(KEYINPUT3), .ZN(n486) );
  XNOR2_X1 U611 ( .A(n441), .B(KEYINPUT124), .ZN(G54) );
  NOR2_X2 U612 ( .A1(n725), .A2(n733), .ZN(n441) );
  XNOR2_X1 U613 ( .A(n442), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U614 ( .A1(n719), .A2(n733), .ZN(n442) );
  XNOR2_X1 U615 ( .A(n443), .B(n653), .ZN(G57) );
  XNOR2_X1 U616 ( .A(n622), .B(n447), .ZN(n446) );
  XNOR2_X2 U617 ( .A(n593), .B(n450), .ZN(n683) );
  XNOR2_X1 U618 ( .A(n618), .B(KEYINPUT34), .ZN(n452) );
  NOR2_X1 U619 ( .A1(n694), .A2(n693), .ZN(n629) );
  NAND2_X1 U620 ( .A1(n557), .A2(G221), .ZN(n520) );
  XNOR2_X2 U621 ( .A(n454), .B(G953), .ZN(n749) );
  XNOR2_X1 U622 ( .A(n578), .B(KEYINPUT46), .ZN(n458) );
  XNOR2_X2 U623 ( .A(n463), .B(n462), .ZN(n745) );
  XNOR2_X2 U624 ( .A(G140), .B(G125), .ZN(n463) );
  XNOR2_X1 U625 ( .A(n472), .B(n471), .ZN(G75) );
  INV_X1 U626 ( .A(KEYINPUT53), .ZN(n471) );
  XNOR2_X1 U627 ( .A(n568), .B(n474), .ZN(n473) );
  INV_X1 U628 ( .A(n745), .ZN(n474) );
  NAND2_X1 U629 ( .A1(n599), .A2(n584), .ZN(n475) );
  XNOR2_X2 U630 ( .A(n550), .B(n344), .ZN(n599) );
  INV_X1 U631 ( .A(n483), .ZN(n661) );
  NAND2_X1 U632 ( .A1(n491), .A2(n487), .ZN(n592) );
  XNOR2_X1 U633 ( .A(n632), .B(KEYINPUT111), .ZN(n491) );
  XNOR2_X1 U634 ( .A(n722), .B(n495), .ZN(n723) );
  XOR2_X1 U635 ( .A(n721), .B(n720), .Z(n495) );
  AND2_X1 U636 ( .A1(G210), .A2(n564), .ZN(n496) );
  XNOR2_X1 U637 ( .A(KEYINPUT59), .B(KEYINPUT69), .ZN(n497) );
  INV_X1 U638 ( .A(KEYINPUT24), .ZN(n516) );
  XNOR2_X1 U639 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U640 ( .A(n503), .B(n496), .ZN(n504) );
  NOR2_X1 U641 ( .A1(n749), .A2(G952), .ZN(n733) );
  XNOR2_X1 U642 ( .A(n502), .B(KEYINPUT5), .ZN(n503) );
  XNOR2_X1 U643 ( .A(n525), .B(KEYINPUT62), .ZN(n651) );
  INV_X1 U644 ( .A(KEYINPUT2), .ZN(n506) );
  INV_X1 U645 ( .A(n648), .ZN(n548) );
  XOR2_X1 U646 ( .A(KEYINPUT84), .B(n548), .Z(n505) );
  XNOR2_X1 U647 ( .A(G107), .B(G110), .ZN(n507) );
  AND2_X1 U648 ( .A1(G227), .A2(n749), .ZN(n508) );
  XOR2_X1 U649 ( .A(KEYINPUT98), .B(KEYINPUT21), .Z(n512) );
  NAND2_X1 U650 ( .A1(G234), .A2(n648), .ZN(n509) );
  XNOR2_X1 U651 ( .A(n510), .B(n509), .ZN(n521) );
  NAND2_X1 U652 ( .A1(n521), .A2(G221), .ZN(n511) );
  XNOR2_X1 U653 ( .A(n512), .B(n511), .ZN(n696) );
  NAND2_X1 U654 ( .A1(n749), .A2(G234), .ZN(n513) );
  XOR2_X1 U655 ( .A(KEYINPUT82), .B(G137), .Z(n515) );
  XNOR2_X1 U656 ( .A(G146), .B(G110), .ZN(n514) );
  NAND2_X1 U657 ( .A1(n521), .A2(G217), .ZN(n522) );
  XOR2_X1 U658 ( .A(KEYINPUT30), .B(KEYINPUT112), .Z(n530) );
  XNOR2_X1 U659 ( .A(KEYINPUT75), .B(G472), .ZN(n526) );
  XNOR2_X2 U660 ( .A(n527), .B(n526), .ZN(n700) );
  NAND2_X1 U661 ( .A1(G214), .A2(n549), .ZN(n528) );
  INV_X1 U662 ( .A(n684), .ZN(n584) );
  NAND2_X1 U663 ( .A1(G237), .A2(G234), .ZN(n531) );
  XNOR2_X1 U664 ( .A(n531), .B(KEYINPUT14), .ZN(n534) );
  NAND2_X1 U665 ( .A1(G952), .A2(n534), .ZN(n532) );
  XNOR2_X1 U666 ( .A(KEYINPUT93), .B(n532), .ZN(n712) );
  AND2_X1 U667 ( .A1(n739), .A2(n712), .ZN(n533) );
  XOR2_X1 U668 ( .A(KEYINPUT94), .B(n533), .Z(n611) );
  NAND2_X1 U669 ( .A1(n534), .A2(G902), .ZN(n535) );
  XNOR2_X1 U670 ( .A(n535), .B(KEYINPUT95), .ZN(n609) );
  NOR2_X1 U671 ( .A1(n749), .A2(G900), .ZN(n536) );
  NAND2_X1 U672 ( .A1(n609), .A2(n536), .ZN(n537) );
  NAND2_X1 U673 ( .A1(n611), .A2(n537), .ZN(n572) );
  XNOR2_X1 U674 ( .A(n734), .B(n541), .ZN(n547) );
  NAND2_X1 U675 ( .A1(G224), .A2(n749), .ZN(n542) );
  XNOR2_X1 U676 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U677 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U678 ( .A(n547), .B(n546), .ZN(n716) );
  XNOR2_X1 U679 ( .A(n552), .B(n551), .ZN(n556) );
  XNOR2_X1 U680 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U681 ( .A(n556), .B(n555), .Z(n559) );
  NAND2_X1 U682 ( .A1(G217), .A2(n557), .ZN(n558) );
  XNOR2_X1 U683 ( .A(n558), .B(n559), .ZN(n560) );
  XNOR2_X1 U684 ( .A(n561), .B(n560), .ZN(n728) );
  XOR2_X1 U685 ( .A(KEYINPUT12), .B(KEYINPUT102), .Z(n566) );
  NAND2_X1 U686 ( .A1(n564), .A2(G214), .ZN(n565) );
  XNOR2_X1 U687 ( .A(KEYINPUT13), .B(G475), .ZN(n569) );
  NAND2_X1 U688 ( .A1(n696), .A2(n572), .ZN(n573) );
  XNOR2_X1 U689 ( .A(KEYINPUT114), .B(KEYINPUT28), .ZN(n574) );
  XNOR2_X1 U690 ( .A(n575), .B(n574), .ZN(n576) );
  NAND2_X1 U691 ( .A1(n582), .A2(n576), .ZN(n587) );
  INV_X1 U692 ( .A(n588), .ZN(n591) );
  INV_X1 U693 ( .A(n620), .ZN(n686) );
  XNOR2_X1 U694 ( .A(n580), .B(KEYINPUT36), .ZN(n583) );
  INV_X1 U695 ( .A(n694), .ZN(n602) );
  NAND2_X1 U696 ( .A1(n583), .A2(n602), .ZN(n676) );
  INV_X1 U697 ( .A(n663), .ZN(n673) );
  NAND2_X1 U698 ( .A1(n589), .A2(n673), .ZN(n687) );
  XNOR2_X1 U699 ( .A(KEYINPUT47), .B(n590), .ZN(n595) );
  NOR2_X1 U700 ( .A1(n619), .A2(n594), .ZN(n666) );
  XNOR2_X1 U701 ( .A(KEYINPUT76), .B(n596), .ZN(n597) );
  NOR2_X1 U702 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U703 ( .A(n603), .B(KEYINPUT43), .ZN(n604) );
  OR2_X1 U704 ( .A1(n673), .A2(n605), .ZN(n677) );
  INV_X1 U705 ( .A(n677), .ZN(n606) );
  XOR2_X1 U706 ( .A(KEYINPUT77), .B(n747), .Z(n647) );
  INV_X1 U707 ( .A(n608), .ZN(n614) );
  NOR2_X1 U708 ( .A1(G898), .A2(n739), .ZN(n735) );
  NAND2_X1 U709 ( .A1(n609), .A2(n735), .ZN(n610) );
  XNOR2_X1 U710 ( .A(n610), .B(KEYINPUT96), .ZN(n612) );
  NAND2_X1 U711 ( .A1(n612), .A2(n611), .ZN(n613) );
  NAND2_X1 U712 ( .A1(n620), .A2(n696), .ZN(n621) );
  NOR2_X1 U713 ( .A1(n694), .A2(n448), .ZN(n623) );
  XOR2_X1 U714 ( .A(KEYINPUT108), .B(n623), .Z(n625) );
  XNOR2_X1 U715 ( .A(n636), .B(KEYINPUT80), .ZN(n624) );
  NOR2_X1 U716 ( .A1(n625), .A2(n624), .ZN(n627) );
  NAND2_X1 U717 ( .A1(n700), .A2(n629), .ZN(n703) );
  NOR2_X1 U718 ( .A1(n630), .A2(n703), .ZN(n631) );
  XNOR2_X1 U719 ( .A(n631), .B(KEYINPUT31), .ZN(n672) );
  NOR2_X1 U720 ( .A1(n700), .A2(n632), .ZN(n634) );
  NAND2_X1 U721 ( .A1(n634), .A2(n633), .ZN(n657) );
  NAND2_X1 U722 ( .A1(n672), .A2(n657), .ZN(n635) );
  NAND2_X1 U723 ( .A1(n635), .A2(n687), .ZN(n640) );
  OR2_X1 U724 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U725 ( .A(n638), .B(KEYINPUT87), .ZN(n639) );
  NAND2_X1 U726 ( .A1(n639), .A2(n448), .ZN(n654) );
  XNOR2_X1 U727 ( .A(KEYINPUT85), .B(KEYINPUT45), .ZN(n642) );
  INV_X1 U728 ( .A(n642), .ZN(n643) );
  INV_X1 U729 ( .A(KEYINPUT78), .ZN(n649) );
  XOR2_X1 U730 ( .A(KEYINPUT63), .B(KEYINPUT88), .Z(n653) );
  XNOR2_X1 U731 ( .A(G101), .B(n654), .ZN(G3) );
  NOR2_X1 U732 ( .A1(n670), .A2(n657), .ZN(n655) );
  XOR2_X1 U733 ( .A(KEYINPUT118), .B(n655), .Z(n656) );
  XNOR2_X1 U734 ( .A(G104), .B(n656), .ZN(G6) );
  NOR2_X1 U735 ( .A1(n673), .A2(n657), .ZN(n659) );
  XNOR2_X1 U736 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n658) );
  XNOR2_X1 U737 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U738 ( .A(G107), .B(n660), .ZN(G9) );
  XNOR2_X1 U739 ( .A(G110), .B(n661), .ZN(n662) );
  XNOR2_X1 U740 ( .A(n662), .B(KEYINPUT119), .ZN(G12) );
  XOR2_X1 U741 ( .A(G128), .B(KEYINPUT29), .Z(n665) );
  NAND2_X1 U742 ( .A1(n667), .A2(n663), .ZN(n664) );
  XNOR2_X1 U743 ( .A(n665), .B(n664), .ZN(G30) );
  XOR2_X1 U744 ( .A(G143), .B(n666), .Z(G45) );
  NAND2_X1 U745 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U746 ( .A(n669), .B(G146), .ZN(G48) );
  NOR2_X1 U747 ( .A1(n670), .A2(n672), .ZN(n671) );
  XOR2_X1 U748 ( .A(G113), .B(n671), .Z(G15) );
  NOR2_X1 U749 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U750 ( .A(G116), .B(n674), .Z(G18) );
  XOR2_X1 U751 ( .A(G125), .B(KEYINPUT37), .Z(n675) );
  XNOR2_X1 U752 ( .A(n676), .B(n675), .ZN(G27) );
  XNOR2_X1 U753 ( .A(G134), .B(n677), .ZN(G36) );
  XOR2_X1 U754 ( .A(G140), .B(n678), .Z(G42) );
  AND2_X1 U755 ( .A1(n740), .A2(n747), .ZN(n679) );
  NOR2_X1 U756 ( .A1(KEYINPUT2), .A2(n679), .ZN(n680) );
  NOR2_X1 U757 ( .A1(n681), .A2(n680), .ZN(n682) );
  AND2_X1 U758 ( .A1(n683), .A2(n684), .ZN(n685) );
  NOR2_X1 U759 ( .A1(n686), .A2(n685), .ZN(n691) );
  INV_X1 U760 ( .A(n687), .ZN(n689) );
  NOR2_X1 U761 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U762 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U763 ( .A1(n713), .A2(n692), .ZN(n708) );
  NAND2_X1 U764 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U765 ( .A(n695), .B(KEYINPUT50), .ZN(n702) );
  NOR2_X1 U766 ( .A1(n448), .A2(n696), .ZN(n698) );
  XOR2_X1 U767 ( .A(KEYINPUT49), .B(n698), .Z(n699) );
  NOR2_X1 U768 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U769 ( .A1(n702), .A2(n701), .ZN(n704) );
  NAND2_X1 U770 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U771 ( .A(KEYINPUT51), .B(n705), .ZN(n706) );
  NOR2_X1 U772 ( .A1(n714), .A2(n706), .ZN(n707) );
  NOR2_X1 U773 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U774 ( .A(n709), .B(KEYINPUT52), .Z(n710) );
  XNOR2_X1 U775 ( .A(KEYINPUT120), .B(n710), .ZN(n711) );
  NOR2_X1 U776 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U777 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n718) );
  XNOR2_X1 U778 ( .A(n716), .B(KEYINPUT89), .ZN(n717) );
  XOR2_X1 U779 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n721) );
  XNOR2_X1 U780 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n720) );
  XNOR2_X1 U781 ( .A(n728), .B(n727), .ZN(n729) );
  NOR2_X1 U782 ( .A1(n733), .A2(n729), .ZN(G63) );
  XNOR2_X1 U783 ( .A(n731), .B(n730), .ZN(n732) );
  NOR2_X1 U784 ( .A1(n733), .A2(n732), .ZN(G66) );
  NOR2_X1 U785 ( .A1(n735), .A2(n734), .ZN(n744) );
  XOR2_X1 U786 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n737) );
  NAND2_X1 U787 ( .A1(G224), .A2(G953), .ZN(n736) );
  XNOR2_X1 U788 ( .A(n737), .B(n736), .ZN(n738) );
  NAND2_X1 U789 ( .A1(n738), .A2(G898), .ZN(n742) );
  NAND2_X1 U790 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U791 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U792 ( .A(n744), .B(n743), .ZN(G69) );
  XOR2_X1 U793 ( .A(n746), .B(n745), .Z(n750) );
  XNOR2_X1 U794 ( .A(n747), .B(n750), .ZN(n748) );
  NAND2_X1 U795 ( .A1(n749), .A2(n748), .ZN(n755) );
  XOR2_X1 U796 ( .A(n750), .B(G227), .Z(n751) );
  XNOR2_X1 U797 ( .A(n751), .B(KEYINPUT126), .ZN(n752) );
  NAND2_X1 U798 ( .A1(n752), .A2(G900), .ZN(n753) );
  NAND2_X1 U799 ( .A1(G953), .A2(n753), .ZN(n754) );
  NAND2_X1 U800 ( .A1(n755), .A2(n754), .ZN(G72) );
  XOR2_X1 U801 ( .A(n756), .B(G122), .Z(G24) );
  XNOR2_X1 U802 ( .A(G137), .B(KEYINPUT127), .ZN(n758) );
  XNOR2_X1 U803 ( .A(n758), .B(n757), .ZN(G39) );
  XOR2_X1 U804 ( .A(n759), .B(G131), .Z(G33) );
endmodule

