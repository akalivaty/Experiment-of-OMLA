//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 1 0 1 0 1 1 1 1 0 0 1 0 1 0 0 0 0 0 1 1 0 0 1 0 0 1 0 0 0 0 0 1 0 0 0 0 0 1 1 1 1 0 0 1 1 1 1 0 0 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n449, new_n451, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n559, new_n561, new_n562, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n631, new_n632, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n448));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  INV_X1    g025(.A(new_n449), .ZN(new_n451));
  NAND2_X1  g026(.A1(new_n451), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n451), .A2(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NAND4_X1  g031(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT67), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n458), .A2(G567), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT68), .Z(new_n462));
  AOI21_X1  g037(.A(new_n462), .B1(new_n456), .B2(G2106), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n463), .B(KEYINPUT69), .ZN(G319));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(new_n465), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G137), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n467), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n471), .A2(G125), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n472), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(KEYINPUT70), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n480));
  AOI22_X1  g055(.A1(new_n471), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n480), .B1(new_n481), .B2(new_n472), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n475), .B1(new_n479), .B2(new_n482), .ZN(G160));
  INV_X1    g058(.A(new_n473), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT71), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G112), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(new_n488), .B2(G2105), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n472), .B1(new_n469), .B2(new_n470), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n489), .B1(G124), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g067(.A(new_n492), .B(KEYINPUT72), .ZN(G162));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n494), .B1(new_n473), .B2(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n471), .A2(KEYINPUT4), .A3(G138), .A4(new_n472), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n490), .A2(G126), .ZN(new_n498));
  OR2_X1    g073(.A1(G102), .A2(G2105), .ZN(new_n499));
  XNOR2_X1  g074(.A(KEYINPUT73), .B(G114), .ZN(new_n500));
  OAI211_X1 g075(.A(G2104), .B(new_n499), .C1(new_n500), .C2(new_n472), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n496), .A2(new_n497), .A3(new_n498), .A4(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n504), .B1(new_n505), .B2(KEYINPUT74), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT74), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(KEYINPUT5), .A3(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT75), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  AND3_X1   g086(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n510), .B1(new_n509), .B2(new_n511), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G88), .ZN(new_n515));
  INV_X1    g090(.A(G62), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n516), .B1(new_n506), .B2(new_n508), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n517), .A2(KEYINPUT76), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n519), .B1(new_n517), .B2(KEYINPUT76), .ZN(new_n520));
  OAI21_X1  g095(.A(G651), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n511), .A2(G543), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G50), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n515), .A2(new_n521), .A3(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  AND2_X1   g101(.A1(G63), .A2(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n509), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  INV_X1    g105(.A(G51), .ZN(new_n531));
  OAI211_X1 g106(.A(new_n528), .B(new_n530), .C1(new_n531), .C2(new_n522), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n532), .B1(new_n514), .B2(G89), .ZN(G168));
  NAND2_X1  g108(.A1(new_n514), .A2(G90), .ZN(new_n534));
  NAND2_X1  g109(.A1(G77), .A2(G543), .ZN(new_n535));
  AND3_X1   g110(.A1(new_n507), .A2(KEYINPUT5), .A3(G543), .ZN(new_n536));
  AOI21_X1  g111(.A(G543), .B1(new_n507), .B2(KEYINPUT5), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(G64), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n535), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n540), .A2(G651), .B1(G52), .B2(new_n523), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n534), .A2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n544), .B1(new_n506), .B2(new_n508), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT77), .ZN(new_n546));
  AND2_X1   g121(.A1(G68), .A2(G543), .ZN(new_n547));
  OR3_X1    g122(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n546), .B1(new_n545), .B2(new_n547), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n548), .A2(G651), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n509), .A2(new_n511), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(KEYINPUT75), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n552), .A2(G81), .A3(new_n553), .ZN(new_n554));
  XNOR2_X1  g129(.A(KEYINPUT78), .B(G43), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n523), .A2(new_n555), .ZN(new_n556));
  AND3_X1   g131(.A1(new_n550), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n559));
  XOR2_X1   g134(.A(new_n559), .B(KEYINPUT79), .Z(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  AND2_X1   g138(.A1(KEYINPUT6), .A2(G651), .ZN(new_n564));
  NOR2_X1   g139(.A1(KEYINPUT6), .A2(G651), .ZN(new_n565));
  OAI211_X1 g140(.A(G53), .B(G543), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT80), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT9), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n566), .A2(new_n567), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n566), .A2(new_n567), .A3(KEYINPUT9), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n514), .A2(G91), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT81), .ZN(new_n573));
  AND3_X1   g148(.A1(new_n506), .A2(new_n573), .A3(new_n508), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n573), .B1(new_n506), .B2(new_n508), .ZN(new_n575));
  OAI21_X1  g150(.A(G65), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(G78), .A2(G543), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g153(.A(KEYINPUT82), .B1(new_n578), .B2(G651), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT82), .ZN(new_n580));
  INV_X1    g155(.A(G651), .ZN(new_n581));
  AOI211_X1 g156(.A(new_n580), .B(new_n581), .C1(new_n576), .C2(new_n577), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n572), .B1(new_n579), .B2(new_n582), .ZN(G299));
  INV_X1    g158(.A(G168), .ZN(G286));
  OR2_X1    g159(.A1(new_n509), .A2(G74), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n585), .A2(G651), .B1(new_n523), .B2(G49), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n552), .A2(new_n553), .ZN(new_n587));
  INV_X1    g162(.A(G87), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(G288));
  INV_X1    g164(.A(KEYINPUT83), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n514), .A2(new_n590), .A3(G86), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n552), .A2(G86), .A3(new_n553), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(KEYINPUT83), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(G73), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G61), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n538), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(G651), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n523), .A2(G48), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n594), .A2(new_n601), .ZN(G305));
  INV_X1    g177(.A(KEYINPUT84), .ZN(new_n603));
  NAND2_X1  g178(.A1(G72), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G60), .ZN(new_n605));
  OAI211_X1 g180(.A(new_n603), .B(new_n604), .C1(new_n538), .C2(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n605), .B1(new_n506), .B2(new_n508), .ZN(new_n607));
  INV_X1    g182(.A(new_n604), .ZN(new_n608));
  OAI21_X1  g183(.A(KEYINPUT84), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n606), .A2(G651), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n523), .A2(G47), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n552), .A2(G85), .A3(new_n553), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(G290));
  NAND2_X1  g188(.A1(G301), .A2(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n523), .A2(G54), .ZN(new_n615));
  NAND2_X1  g190(.A1(G79), .A2(G543), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(KEYINPUT81), .B1(new_n536), .B2(new_n537), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n506), .A2(new_n573), .A3(new_n508), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(KEYINPUT85), .B(G66), .Z(new_n621));
  AOI21_X1  g196(.A(new_n617), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n615), .B1(new_n622), .B2(new_n581), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n552), .A2(G92), .A3(new_n553), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT10), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n514), .A2(KEYINPUT10), .A3(G92), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n623), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n614), .B1(new_n628), .B2(G868), .ZN(G284));
  OAI21_X1  g204(.A(new_n614), .B1(new_n628), .B2(G868), .ZN(G321));
  NAND2_X1  g205(.A1(G286), .A2(G868), .ZN(new_n631));
  INV_X1    g206(.A(G299), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(new_n632), .B2(G868), .ZN(G297));
  OAI21_X1  g208(.A(new_n631), .B1(new_n632), .B2(G868), .ZN(G280));
  XNOR2_X1  g209(.A(KEYINPUT86), .B(G559), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n628), .B1(G860), .B2(new_n635), .ZN(G148));
  NAND3_X1  g211(.A1(new_n550), .A2(new_n554), .A3(new_n556), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n637), .A2(G868), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n628), .A2(new_n635), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT87), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n638), .B1(new_n640), .B2(G868), .ZN(G323));
  XNOR2_X1  g216(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g217(.A1(new_n471), .A2(new_n466), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT12), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT13), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n646), .A2(G2100), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n490), .A2(G123), .ZN(new_n648));
  INV_X1    g223(.A(KEYINPUT88), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n651));
  INV_X1    g226(.A(G111), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n651), .B1(new_n652), .B2(G2105), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n653), .B1(new_n484), .B2(G135), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n655), .A2(G2096), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n646), .A2(G2100), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(G2096), .ZN(new_n658));
  NAND4_X1  g233(.A1(new_n647), .A2(new_n656), .A3(new_n657), .A4(new_n658), .ZN(G156));
  XNOR2_X1  g234(.A(G2427), .B(G2438), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2430), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT15), .B(G2435), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n663), .A2(KEYINPUT14), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G1341), .B(G1348), .Z(new_n666));
  XNOR2_X1  g241(.A(G2443), .B(G2446), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n665), .B(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G2451), .B(G2454), .Z(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT89), .B(KEYINPUT16), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(G14), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n669), .A2(new_n672), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(G401));
  XOR2_X1   g251(.A(G2084), .B(G2090), .Z(new_n677));
  XOR2_X1   g252(.A(G2067), .B(G2678), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT90), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT91), .Z(new_n680));
  XOR2_X1   g255(.A(G2072), .B(G2078), .Z(new_n681));
  AOI21_X1  g256(.A(new_n677), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT92), .B(KEYINPUT17), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n681), .B(new_n683), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n682), .B1(new_n680), .B2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n677), .ZN(new_n686));
  NOR3_X1   g261(.A1(new_n679), .A2(new_n681), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT18), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n680), .A2(new_n684), .A3(new_n677), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n685), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G2096), .B(G2100), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(G227));
  XNOR2_X1  g267(.A(G1971), .B(G1976), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT19), .ZN(new_n694));
  XOR2_X1   g269(.A(G1956), .B(G2474), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT93), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1961), .B(G1966), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT94), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n694), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(new_n700), .B2(new_n699), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT20), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n696), .A2(new_n698), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n704), .A2(new_n699), .A3(new_n694), .ZN(new_n705));
  OAI211_X1 g280(.A(new_n703), .B(new_n705), .C1(new_n694), .C2(new_n704), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1991), .B(G1996), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  XNOR2_X1  g286(.A(G1981), .B(G1986), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  OR3_X1    g288(.A1(new_n710), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n710), .B2(new_n711), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n714), .A2(new_n715), .ZN(G229));
  NAND2_X1  g291(.A1(new_n514), .A2(G87), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n717), .A2(KEYINPUT95), .A3(new_n586), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(KEYINPUT95), .B1(new_n717), .B2(new_n586), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G16), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G16), .B2(G23), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT33), .B(G1976), .Z(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n600), .B1(new_n591), .B2(new_n593), .ZN(new_n727));
  INV_X1    g302(.A(G16), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G6), .B2(new_n728), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT32), .B(G1981), .Z(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n726), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n728), .A2(G22), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT96), .Z(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G303), .B2(G16), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G1971), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n731), .B2(new_n730), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n723), .A2(new_n725), .ZN(new_n739));
  NOR3_X1   g314(.A1(new_n733), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT34), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  INV_X1    g318(.A(G29), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G25), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n484), .A2(G131), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n490), .A2(G119), .ZN(new_n747));
  OR2_X1    g322(.A1(G95), .A2(G2105), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n748), .B(G2104), .C1(G107), .C2(new_n472), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n746), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n745), .B1(new_n751), .B2(new_n744), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT35), .B(G1991), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(G1986), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n728), .A2(G24), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G290), .B2(G16), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n754), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n755), .B2(new_n757), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n742), .A2(new_n743), .A3(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT36), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT99), .B(KEYINPUT28), .Z(new_n763));
  NAND2_X1  g338(.A1(new_n744), .A2(G26), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n490), .A2(G128), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n472), .A2(G116), .ZN(new_n767));
  OAI21_X1  g342(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n768));
  INV_X1    g343(.A(G140), .ZN(new_n769));
  OAI221_X1 g344(.A(new_n766), .B1(new_n767), .B2(new_n768), .C1(new_n769), .C2(new_n473), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT97), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  AND3_X1   g347(.A1(new_n772), .A2(KEYINPUT98), .A3(G29), .ZN(new_n773));
  AOI21_X1  g348(.A(KEYINPUT98), .B1(new_n772), .B2(G29), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n765), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(G2067), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n744), .A2(G32), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n484), .A2(G141), .B1(G105), .B2(new_n466), .ZN(new_n779));
  NAND3_X1  g354(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT26), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G129), .B2(new_n490), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n778), .B1(new_n784), .B2(new_n744), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT27), .B(G1996), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(G5), .A2(G16), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT103), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G301), .B2(new_n728), .ZN(new_n790));
  INV_X1    g365(.A(G1961), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT101), .B(KEYINPUT24), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G34), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n793), .A2(G29), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G160), .B2(G29), .ZN(new_n795));
  OAI22_X1  g370(.A1(new_n790), .A2(new_n791), .B1(new_n795), .B2(G2084), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT30), .B(G28), .ZN(new_n797));
  OR2_X1    g372(.A1(KEYINPUT31), .A2(G11), .ZN(new_n798));
  NAND2_X1  g373(.A1(KEYINPUT31), .A2(G11), .ZN(new_n799));
  AOI22_X1  g374(.A1(new_n797), .A2(new_n744), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n655), .B2(new_n744), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n801), .A2(KEYINPUT102), .ZN(new_n802));
  AND2_X1   g377(.A1(new_n801), .A2(KEYINPUT102), .ZN(new_n803));
  NOR4_X1   g378(.A1(new_n787), .A2(new_n796), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n728), .A2(G19), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(new_n557), .B2(new_n728), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(G1341), .Z(new_n807));
  NAND3_X1  g382(.A1(new_n777), .A2(new_n804), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n744), .A2(G27), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G164), .B2(new_n744), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G2078), .ZN(new_n811));
  OR2_X1    g386(.A1(G29), .A2(G33), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n471), .A2(G127), .ZN(new_n813));
  NAND2_X1  g388(.A1(G115), .A2(G2104), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n472), .B1(new_n815), .B2(KEYINPUT100), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(KEYINPUT100), .B2(new_n815), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT25), .ZN(new_n818));
  NAND2_X1  g393(.A1(G103), .A2(G2104), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n819), .B2(G2105), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n472), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n484), .A2(G139), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n817), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n812), .B1(new_n823), .B2(new_n744), .ZN(new_n824));
  INV_X1    g399(.A(G2072), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n728), .A2(G21), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(G168), .B2(new_n728), .ZN(new_n827));
  OAI22_X1  g402(.A1(new_n824), .A2(new_n825), .B1(G1966), .B2(new_n827), .ZN(new_n828));
  AOI211_X1 g403(.A(new_n811), .B(new_n828), .C1(new_n791), .C2(new_n790), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n827), .A2(G1966), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n824), .A2(new_n825), .B1(G2084), .B2(new_n795), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n728), .A2(G4), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n628), .B2(new_n728), .ZN(new_n833));
  INV_X1    g408(.A(G1348), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n829), .A2(new_n830), .A3(new_n831), .A4(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n808), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(G29), .A2(G35), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(G162), .B2(G29), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT29), .ZN(new_n840));
  INV_X1    g415(.A(G2090), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n728), .A2(G20), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT23), .Z(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(G299), .B2(G16), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(G1956), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n837), .A2(new_n842), .A3(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n762), .A2(new_n847), .ZN(G311));
  OR2_X1    g423(.A1(new_n762), .A2(new_n847), .ZN(G150));
  NAND2_X1  g424(.A1(new_n628), .A2(G559), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT38), .ZN(new_n851));
  NAND2_X1  g426(.A1(G80), .A2(G543), .ZN(new_n852));
  INV_X1    g427(.A(G67), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n852), .B1(new_n538), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n581), .B1(new_n854), .B2(KEYINPUT104), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(KEYINPUT104), .B2(new_n854), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n552), .A2(G93), .A3(new_n553), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT105), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n523), .A2(G55), .ZN(new_n859));
  AND3_X1   g434(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n858), .B1(new_n857), .B2(new_n859), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n856), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n862), .A2(new_n637), .ZN(new_n863));
  INV_X1    g438(.A(G93), .ZN(new_n864));
  NOR3_X1   g439(.A1(new_n512), .A2(new_n513), .A3(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n859), .ZN(new_n866));
  OAI21_X1  g441(.A(KEYINPUT105), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n557), .B1(new_n869), .B2(new_n856), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n863), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n851), .B(new_n871), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n872), .A2(KEYINPUT39), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(KEYINPUT39), .ZN(new_n874));
  XNOR2_X1  g449(.A(KEYINPUT106), .B(G860), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n862), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n877), .A2(new_n875), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT37), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n876), .A2(new_n879), .ZN(G145));
  INV_X1    g455(.A(KEYINPUT40), .ZN(new_n881));
  INV_X1    g456(.A(G160), .ZN(new_n882));
  OR2_X1    g457(.A1(G162), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n655), .ZN(new_n884));
  NAND2_X1  g459(.A1(G162), .A2(new_n882), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n884), .B1(new_n883), .B2(new_n885), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n823), .A2(KEYINPUT108), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(new_n784), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n889), .A2(new_n784), .ZN(new_n892));
  NOR3_X1   g467(.A1(new_n891), .A2(new_n771), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n771), .B1(new_n891), .B2(new_n892), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n502), .A2(KEYINPUT107), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n501), .A2(new_n498), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT107), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n897), .A2(new_n898), .A3(new_n497), .A4(new_n496), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n894), .A2(new_n895), .A3(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n900), .ZN(new_n902));
  INV_X1    g477(.A(new_n892), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n772), .B1(new_n903), .B2(new_n890), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n902), .B1(new_n904), .B2(new_n893), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n901), .A2(new_n905), .ZN(new_n906));
  XOR2_X1   g481(.A(new_n750), .B(new_n644), .Z(new_n907));
  NAND2_X1  g482(.A1(new_n484), .A2(G142), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT109), .ZN(new_n909));
  OR3_X1    g484(.A1(new_n909), .A2(new_n472), .A3(G118), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n909), .B1(new_n472), .B2(G118), .ZN(new_n911));
  OR2_X1    g486(.A1(G106), .A2(G2105), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n910), .A2(G2104), .A3(new_n911), .A4(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n490), .A2(G130), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n908), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n907), .B(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n906), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT111), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n888), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n916), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n901), .A2(new_n920), .A3(new_n905), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT110), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT110), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n901), .A2(new_n905), .A3(new_n923), .A4(new_n920), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n920), .B1(new_n901), .B2(new_n905), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT111), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n919), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(G37), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n926), .B1(new_n922), .B2(new_n924), .ZN(new_n930));
  INV_X1    g505(.A(new_n888), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n881), .B1(new_n928), .B2(new_n932), .ZN(new_n933));
  OR2_X1    g508(.A1(new_n930), .A2(new_n931), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n919), .A2(new_n925), .A3(new_n927), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n934), .A2(KEYINPUT40), .A3(new_n929), .A4(new_n935), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n933), .A2(new_n936), .ZN(G395));
  OAI21_X1  g512(.A(KEYINPUT113), .B1(new_n628), .B2(G299), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n628), .A2(G299), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n627), .A2(new_n626), .ZN(new_n940));
  INV_X1    g515(.A(new_n615), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n620), .A2(new_n621), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n616), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n941), .B1(new_n943), .B2(G651), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n940), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT113), .ZN(new_n946));
  INV_X1    g521(.A(G65), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n947), .B1(new_n618), .B2(new_n619), .ZN(new_n948));
  INV_X1    g523(.A(new_n577), .ZN(new_n949));
  OAI21_X1  g524(.A(G651), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n580), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n578), .A2(KEYINPUT82), .A3(G651), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n945), .A2(new_n946), .A3(new_n953), .A4(new_n572), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n938), .A2(new_n939), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT41), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n632), .A2(new_n945), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n956), .B1(new_n628), .B2(G299), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n955), .A2(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT112), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n871), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n862), .A2(new_n637), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n869), .A2(new_n557), .A3(new_n856), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT112), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n640), .A2(new_n961), .A3(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n640), .B1(new_n965), .B2(new_n961), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n959), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n961), .A2(new_n965), .ZN(new_n970));
  INV_X1    g545(.A(new_n640), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n945), .B(G299), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(new_n973), .A3(new_n966), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n969), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT42), .ZN(new_n976));
  AOI22_X1  g551(.A1(new_n514), .A2(G85), .B1(G47), .B2(new_n523), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT114), .B1(new_n977), .B2(new_n610), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT114), .ZN(new_n979));
  NOR2_X1   g554(.A1(G290), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n727), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(G290), .A2(new_n979), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n977), .A2(KEYINPUT114), .A3(new_n610), .ZN(new_n983));
  NAND3_X1  g558(.A1(G305), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(G166), .B1(new_n719), .B2(new_n720), .ZN(new_n986));
  INV_X1    g561(.A(new_n720), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n987), .A2(G303), .A3(new_n718), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n985), .A2(new_n989), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n981), .A2(new_n984), .A3(new_n986), .A4(new_n988), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT42), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n969), .A2(new_n993), .A3(new_n974), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n976), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n992), .B1(new_n976), .B2(new_n994), .ZN(new_n996));
  OAI21_X1  g571(.A(G868), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(G868), .B2(new_n877), .ZN(G295));
  OAI21_X1  g573(.A(new_n997), .B1(G868), .B2(new_n877), .ZN(G331));
  AND2_X1   g574(.A1(new_n990), .A2(new_n991), .ZN(new_n1000));
  NAND2_X1  g575(.A1(G301), .A2(G168), .ZN(new_n1001));
  INV_X1    g576(.A(G89), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n587), .A2(new_n1002), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n534), .B(new_n541), .C1(new_n1003), .C2(new_n532), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1005), .B1(new_n863), .B2(new_n870), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1005), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1007), .A2(new_n962), .A3(new_n963), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n973), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1000), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n955), .A2(new_n956), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n957), .A2(new_n958), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1009), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n1012), .A2(new_n1015), .A3(KEYINPUT115), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1009), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n973), .B1(new_n1008), .B2(new_n1006), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1021), .A2(new_n992), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1017), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  OR2_X1    g598(.A1(new_n1016), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT43), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1011), .B1(new_n959), .B2(new_n1009), .ZN(new_n1026));
  AOI21_X1  g601(.A(G37), .B1(new_n1026), .B2(new_n992), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1024), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1010), .B1(new_n1009), .B2(new_n956), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n938), .A2(new_n958), .A3(new_n954), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1029), .B1(new_n1009), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(G37), .B1(new_n1031), .B2(new_n992), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n1024), .A2(new_n1032), .ZN(new_n1033));
  OAI211_X1 g608(.A(KEYINPUT44), .B(new_n1028), .C1(new_n1033), .C2(new_n1025), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT116), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1027), .B1(new_n1016), .B2(new_n1023), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT43), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1032), .B(new_n1025), .C1(new_n1023), .C2(new_n1016), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT44), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1035), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  AOI211_X1 g616(.A(KEYINPUT116), .B(KEYINPUT44), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1034), .B1(new_n1041), .B2(new_n1042), .ZN(G397));
  INV_X1    g618(.A(G1384), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n900), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT45), .ZN(new_n1046));
  INV_X1    g621(.A(G40), .ZN(new_n1047));
  AOI211_X1 g622(.A(new_n1047), .B(new_n475), .C1(new_n479), .C2(new_n482), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1045), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n771), .B(G2067), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1050), .B1(new_n1052), .B2(new_n783), .ZN(new_n1053));
  INV_X1    g628(.A(G1996), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1050), .A2(new_n1054), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1055), .A2(KEYINPUT46), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1055), .A2(KEYINPUT46), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1053), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  XOR2_X1   g633(.A(new_n1058), .B(KEYINPUT47), .Z(new_n1059));
  XNOR2_X1  g634(.A(new_n783), .B(new_n1054), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1051), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n751), .A2(new_n753), .ZN(new_n1062));
  OAI22_X1  g637(.A1(new_n1061), .A2(new_n1062), .B1(G2067), .B2(new_n772), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n1050), .ZN(new_n1064));
  XOR2_X1   g639(.A(new_n750), .B(new_n753), .Z(new_n1065));
  OAI21_X1  g640(.A(new_n1050), .B1(new_n1061), .B2(new_n1065), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n1049), .A2(G1986), .A3(G290), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1066), .B1(KEYINPUT48), .B2(new_n1067), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n1067), .A2(KEYINPUT48), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1064), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1059), .A2(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g646(.A(KEYINPUT118), .B(G8), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n475), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n478), .A2(KEYINPUT70), .ZN(new_n1075));
  NOR3_X1   g650(.A1(new_n481), .A2(new_n480), .A3(new_n472), .ZN(new_n1076));
  OAI211_X1 g651(.A(G40), .B(new_n1074), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n502), .A2(new_n1044), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1073), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT119), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1081), .B(new_n1073), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(G1981), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n727), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n601), .A2(new_n592), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(G1981), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT49), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1085), .A2(new_n1087), .A3(KEYINPUT49), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1090), .A2(new_n1083), .A3(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(G288), .A2(G1976), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1085), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1083), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n721), .A2(G1976), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1083), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT120), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1098), .A2(new_n1099), .A3(KEYINPUT52), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1080), .A2(new_n1082), .B1(new_n721), .B2(G1976), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT52), .ZN(new_n1102));
  OAI21_X1  g677(.A(KEYINPUT120), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(G1976), .ZN(new_n1104));
  AOI21_X1  g679(.A(KEYINPUT52), .B1(G288), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1100), .A2(new_n1103), .A3(new_n1092), .A4(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT55), .ZN(new_n1108));
  INV_X1    g683(.A(G8), .ZN(new_n1109));
  NOR3_X1   g684(.A1(G166), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1111));
  OR2_X1    g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1046), .A2(G1384), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n896), .A2(new_n899), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1078), .A2(new_n1046), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1114), .A2(new_n1048), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(G1971), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1078), .A2(KEYINPUT50), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT50), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n502), .A2(new_n1120), .A3(new_n1044), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1119), .A2(new_n1048), .A3(new_n841), .A4(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1118), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1112), .A2(G8), .A3(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1096), .B1(new_n1107), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT62), .ZN(new_n1126));
  NOR2_X1   g701(.A1(G168), .A2(new_n1072), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT51), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n502), .A2(new_n1113), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1115), .A2(new_n1048), .A3(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1119), .A2(new_n1048), .A3(new_n1121), .ZN(new_n1133));
  OAI22_X1  g708(.A1(new_n1132), .A2(G1966), .B1(G2084), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1130), .B1(new_n1134), .B2(new_n1073), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1133), .ZN(new_n1136));
  INV_X1    g711(.A(G2084), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1115), .A2(new_n1048), .A3(new_n1131), .ZN(new_n1138));
  INV_X1    g713(.A(G1966), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1136), .A2(new_n1137), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1128), .B1(new_n1140), .B2(new_n1109), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1135), .B1(new_n1141), .B2(KEYINPUT51), .ZN(new_n1142));
  NOR3_X1   g717(.A1(new_n1140), .A2(KEYINPUT125), .A3(new_n1128), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT125), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1144), .B1(new_n1134), .B2(new_n1127), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1126), .B1(new_n1142), .B2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1127), .B1(new_n1134), .B2(G8), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1140), .A2(new_n1072), .ZN(new_n1149));
  OAI22_X1  g724(.A1(new_n1148), .A2(new_n1129), .B1(new_n1149), .B2(new_n1130), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1145), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1134), .A2(new_n1144), .A3(new_n1127), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1150), .A2(new_n1153), .A3(KEYINPUT62), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1147), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1077), .B1(new_n1046), .B2(new_n1078), .ZN(new_n1156));
  AOI21_X1  g731(.A(G1971), .B1(new_n1156), .B2(new_n1114), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1122), .ZN(new_n1158));
  OAI21_X1  g733(.A(KEYINPUT121), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT121), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1118), .A2(new_n1160), .A3(new_n1122), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1159), .A2(new_n1073), .A3(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n1124), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT53), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1166), .B1(new_n1116), .B2(G2078), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1133), .A2(new_n791), .ZN(new_n1168));
  AND2_X1   g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(G2078), .ZN(new_n1170));
  AOI21_X1  g745(.A(KEYINPUT126), .B1(new_n1132), .B2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1132), .A2(KEYINPUT126), .A3(new_n1170), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(KEYINPUT53), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1169), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(G171), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n1165), .A2(new_n1175), .A3(new_n1107), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1125), .B1(new_n1155), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1107), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1149), .A2(G168), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1112), .B1(G8), .B2(new_n1123), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1178), .A2(KEYINPUT63), .A3(new_n1124), .A4(new_n1181), .ZN(new_n1182));
  NOR3_X1   g757(.A1(new_n1165), .A2(new_n1107), .A3(new_n1179), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1182), .B1(new_n1183), .B2(KEYINPUT63), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1177), .A2(new_n1184), .ZN(new_n1185));
  XOR2_X1   g760(.A(KEYINPUT56), .B(G2072), .Z(new_n1186));
  OAI22_X1  g761(.A1(new_n1136), .A2(G1956), .B1(new_n1116), .B2(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g762(.A(G299), .B(KEYINPUT57), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1192), .A2(KEYINPUT122), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT122), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1187), .A2(new_n1188), .A3(new_n1194), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1191), .A2(new_n1193), .A3(new_n1195), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1156), .A2(new_n1054), .A3(new_n1114), .ZN(new_n1197));
  XNOR2_X1  g772(.A(KEYINPUT123), .B(KEYINPUT58), .ZN(new_n1198));
  XNOR2_X1  g773(.A(new_n1198), .B(G1341), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1199), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n637), .B1(new_n1197), .B2(new_n1200), .ZN(new_n1201));
  AND2_X1   g776(.A1(new_n1201), .A2(KEYINPUT59), .ZN(new_n1202));
  NOR3_X1   g777(.A1(new_n1077), .A2(new_n1078), .A3(G2067), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n1203), .B1(new_n1133), .B2(new_n834), .ZN(new_n1204));
  INV_X1    g779(.A(KEYINPUT60), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1204), .A2(new_n1205), .A3(new_n628), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1206), .B1(new_n1201), .B2(KEYINPUT59), .ZN(new_n1207));
  NOR2_X1   g782(.A1(new_n1202), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g783(.A(new_n1192), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1190), .B1(new_n1209), .B2(new_n1189), .ZN(new_n1210));
  AND2_X1   g785(.A1(new_n1204), .A2(new_n945), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n1204), .A2(new_n945), .ZN(new_n1212));
  OAI21_X1  g787(.A(KEYINPUT60), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  NAND4_X1  g788(.A1(new_n1196), .A2(new_n1208), .A3(new_n1210), .A4(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1193), .A2(new_n1195), .ZN(new_n1215));
  OAI22_X1  g790(.A1(new_n1215), .A2(new_n1212), .B1(new_n1188), .B2(new_n1187), .ZN(new_n1216));
  NAND3_X1  g791(.A1(new_n1214), .A2(KEYINPUT124), .A3(new_n1216), .ZN(new_n1217));
  INV_X1    g792(.A(new_n1217), .ZN(new_n1218));
  AOI21_X1  g793(.A(KEYINPUT124), .B1(new_n1214), .B2(new_n1216), .ZN(new_n1219));
  NOR2_X1   g794(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g795(.A(KEYINPUT127), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1150), .A2(new_n1153), .ZN(new_n1222));
  INV_X1    g797(.A(KEYINPUT54), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1224));
  NAND3_X1  g799(.A1(new_n1170), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1225));
  NOR3_X1   g800(.A1(new_n475), .A2(new_n478), .A3(new_n1225), .ZN(new_n1226));
  NAND3_X1  g801(.A1(new_n1224), .A2(new_n1114), .A3(new_n1226), .ZN(new_n1227));
  NAND3_X1  g802(.A1(new_n1227), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1228));
  AOI21_X1  g803(.A(new_n1223), .B1(new_n1228), .B2(G171), .ZN(new_n1229));
  OAI211_X1 g804(.A(new_n1169), .B(G301), .C1(new_n1171), .C2(new_n1173), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  AND3_X1   g806(.A1(new_n1112), .A2(G8), .A3(new_n1123), .ZN(new_n1232));
  AOI21_X1  g807(.A(new_n1232), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1233));
  NAND4_X1  g808(.A1(new_n1222), .A2(new_n1178), .A3(new_n1231), .A4(new_n1233), .ZN(new_n1234));
  NAND3_X1  g809(.A1(new_n1169), .A2(G301), .A3(new_n1227), .ZN(new_n1235));
  AOI21_X1  g810(.A(KEYINPUT54), .B1(new_n1175), .B2(new_n1235), .ZN(new_n1236));
  OAI21_X1  g811(.A(new_n1221), .B1(new_n1234), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g812(.A(new_n1236), .ZN(new_n1238));
  NOR2_X1   g813(.A1(new_n1165), .A2(new_n1107), .ZN(new_n1239));
  AOI22_X1  g814(.A1(new_n1150), .A2(new_n1153), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1240));
  NAND4_X1  g815(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .A4(KEYINPUT127), .ZN(new_n1241));
  NAND2_X1  g816(.A1(new_n1237), .A2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g817(.A(new_n1185), .B1(new_n1220), .B2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g818(.A(new_n755), .B1(new_n977), .B2(new_n610), .ZN(new_n1244));
  AOI21_X1  g819(.A(new_n1067), .B1(new_n1050), .B2(new_n1244), .ZN(new_n1245));
  XNOR2_X1  g820(.A(new_n1245), .B(KEYINPUT117), .ZN(new_n1246));
  NAND2_X1  g821(.A1(new_n1246), .A2(new_n1066), .ZN(new_n1247));
  OAI21_X1  g822(.A(new_n1071), .B1(new_n1243), .B2(new_n1247), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g823(.A1(new_n934), .A2(new_n929), .A3(new_n935), .ZN(new_n1250));
  OAI21_X1  g824(.A(new_n463), .B1(new_n674), .B2(new_n675), .ZN(new_n1251));
  NOR2_X1   g825(.A1(G227), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g826(.A(new_n1252), .ZN(new_n1253));
  AOI21_X1  g827(.A(new_n1253), .B1(new_n714), .B2(new_n715), .ZN(new_n1254));
  AND3_X1   g828(.A1(new_n1250), .A2(new_n1254), .A3(new_n1039), .ZN(G308));
  NAND3_X1  g829(.A1(new_n1250), .A2(new_n1254), .A3(new_n1039), .ZN(G225));
endmodule


