

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597;

  XNOR2_X1 U326 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U327 ( .A(n336), .B(n335), .ZN(n340) );
  NOR2_X1 U328 ( .A1(n472), .A2(n498), .ZN(n473) );
  XNOR2_X1 U329 ( .A(n463), .B(KEYINPUT119), .ZN(n464) );
  NOR2_X1 U330 ( .A1(n462), .A2(n461), .ZN(n465) );
  XNOR2_X1 U331 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U332 ( .A(n322), .B(n321), .ZN(n323) );
  NOR2_X1 U333 ( .A1(n550), .A2(n500), .ZN(n578) );
  XOR2_X1 U334 ( .A(n393), .B(n392), .Z(n574) );
  NOR2_X1 U335 ( .A1(n550), .A2(n467), .ZN(n561) );
  XOR2_X1 U336 ( .A(n381), .B(n423), .Z(n294) );
  XOR2_X1 U337 ( .A(n421), .B(n420), .Z(n295) );
  XOR2_X1 U338 ( .A(G218GAT), .B(G106GAT), .Z(n296) );
  XOR2_X1 U339 ( .A(G204GAT), .B(KEYINPUT99), .Z(n297) );
  NOR2_X1 U340 ( .A1(n591), .A2(n454), .ZN(n455) );
  INV_X1 U341 ( .A(KEYINPUT94), .ZN(n321) );
  XNOR2_X1 U342 ( .A(KEYINPUT47), .B(KEYINPUT116), .ZN(n459) );
  INV_X1 U343 ( .A(KEYINPUT102), .ZN(n479) );
  INV_X1 U344 ( .A(KEYINPUT48), .ZN(n463) );
  XOR2_X1 U345 ( .A(G22GAT), .B(G155GAT), .Z(n395) );
  INV_X1 U346 ( .A(n395), .ZN(n333) );
  XNOR2_X1 U347 ( .A(n377), .B(n296), .ZN(n378) );
  XNOR2_X1 U348 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U349 ( .A(n494), .B(KEYINPUT123), .ZN(n495) );
  XNOR2_X1 U350 ( .A(n379), .B(n378), .ZN(n383) );
  XNOR2_X1 U351 ( .A(n396), .B(n297), .ZN(n362) );
  XNOR2_X1 U352 ( .A(n466), .B(KEYINPUT120), .ZN(n564) );
  XNOR2_X1 U353 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U354 ( .A(n426), .B(n425), .Z(n588) );
  XNOR2_X1 U355 ( .A(n413), .B(n412), .ZN(n591) );
  INV_X1 U356 ( .A(G134GAT), .ZN(n468) );
  INV_X1 U357 ( .A(G43GAT), .ZN(n504) );
  XOR2_X1 U358 ( .A(n367), .B(n366), .Z(n548) );
  XNOR2_X1 U359 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n508) );
  XNOR2_X1 U360 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U361 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U362 ( .A(n509), .B(n508), .ZN(G1351GAT) );
  XNOR2_X1 U363 ( .A(n507), .B(n506), .ZN(G1330GAT) );
  XOR2_X1 U364 ( .A(KEYINPUT87), .B(KEYINPUT88), .Z(n299) );
  XNOR2_X1 U365 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n298) );
  XNOR2_X1 U366 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U367 ( .A(G113GAT), .B(n300), .Z(n346) );
  XOR2_X1 U368 ( .A(KEYINPUT89), .B(KEYINPUT20), .Z(n302) );
  XNOR2_X1 U369 ( .A(G183GAT), .B(KEYINPUT90), .ZN(n301) );
  XNOR2_X1 U370 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U371 ( .A(G71GAT), .B(G176GAT), .Z(n304) );
  XNOR2_X1 U372 ( .A(KEYINPUT92), .B(KEYINPUT65), .ZN(n303) );
  XNOR2_X1 U373 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U374 ( .A(n306), .B(n305), .Z(n317) );
  XOR2_X1 U375 ( .A(KEYINPUT17), .B(KEYINPUT91), .Z(n308) );
  XNOR2_X1 U376 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n307) );
  XNOR2_X1 U377 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U378 ( .A(G169GAT), .B(n309), .Z(n365) );
  XOR2_X1 U379 ( .A(G15GAT), .B(G127GAT), .Z(n406) );
  XOR2_X1 U380 ( .A(G134GAT), .B(G190GAT), .Z(n311) );
  XNOR2_X1 U381 ( .A(G43GAT), .B(G99GAT), .ZN(n310) );
  XNOR2_X1 U382 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U383 ( .A(n406), .B(n312), .Z(n314) );
  NAND2_X1 U384 ( .A1(G227GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U385 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U386 ( .A(n365), .B(n315), .ZN(n316) );
  XNOR2_X1 U387 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U388 ( .A(n346), .B(n318), .ZN(n550) );
  XOR2_X1 U389 ( .A(KEYINPUT97), .B(KEYINPUT22), .Z(n320) );
  XNOR2_X1 U390 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n319) );
  XNOR2_X1 U391 ( .A(n320), .B(n319), .ZN(n324) );
  NAND2_X1 U392 ( .A1(G228GAT), .A2(G233GAT), .ZN(n322) );
  XOR2_X1 U393 ( .A(n325), .B(KEYINPUT93), .Z(n331) );
  XNOR2_X1 U394 ( .A(G148GAT), .B(KEYINPUT76), .ZN(n326) );
  XNOR2_X1 U395 ( .A(n326), .B(KEYINPUT77), .ZN(n327) );
  XOR2_X1 U396 ( .A(n327), .B(G204GAT), .Z(n329) );
  XNOR2_X1 U397 ( .A(G78GAT), .B(G106GAT), .ZN(n328) );
  XNOR2_X1 U398 ( .A(n329), .B(n328), .ZN(n424) );
  XNOR2_X1 U399 ( .A(n424), .B(KEYINPUT96), .ZN(n330) );
  XNOR2_X1 U400 ( .A(n331), .B(n330), .ZN(n336) );
  XOR2_X1 U401 ( .A(G50GAT), .B(G162GAT), .Z(n372) );
  XNOR2_X1 U402 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n332) );
  XNOR2_X1 U403 ( .A(n332), .B(KEYINPUT2), .ZN(n342) );
  XNOR2_X1 U404 ( .A(n372), .B(n342), .ZN(n334) );
  XOR2_X1 U405 ( .A(KEYINPUT21), .B(G218GAT), .Z(n338) );
  XNOR2_X1 U406 ( .A(KEYINPUT95), .B(G211GAT), .ZN(n337) );
  XNOR2_X1 U407 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U408 ( .A(G197GAT), .B(n339), .ZN(n366) );
  XNOR2_X1 U409 ( .A(n340), .B(n366), .ZN(n498) );
  XNOR2_X1 U410 ( .A(n498), .B(KEYINPUT28), .ZN(n341) );
  XNOR2_X1 U411 ( .A(n341), .B(KEYINPUT67), .ZN(n553) );
  XOR2_X1 U412 ( .A(G134GAT), .B(KEYINPUT80), .Z(n377) );
  XOR2_X1 U413 ( .A(n377), .B(G85GAT), .Z(n344) );
  XNOR2_X1 U414 ( .A(G162GAT), .B(n342), .ZN(n343) );
  XNOR2_X1 U415 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U416 ( .A(n346), .B(n345), .ZN(n359) );
  XOR2_X1 U417 ( .A(G155GAT), .B(G148GAT), .Z(n348) );
  XNOR2_X1 U418 ( .A(G29GAT), .B(G127GAT), .ZN(n347) );
  XNOR2_X1 U419 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U420 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n350) );
  XNOR2_X1 U421 ( .A(G1GAT), .B(G57GAT), .ZN(n349) );
  XNOR2_X1 U422 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U423 ( .A(n352), .B(n351), .Z(n357) );
  XOR2_X1 U424 ( .A(KEYINPUT98), .B(KEYINPUT1), .Z(n354) );
  NAND2_X1 U425 ( .A1(G225GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U426 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U427 ( .A(KEYINPUT6), .B(n355), .ZN(n356) );
  XNOR2_X1 U428 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U429 ( .A(n359), .B(n358), .ZN(n546) );
  XOR2_X1 U430 ( .A(G36GAT), .B(G190GAT), .Z(n381) );
  XNOR2_X1 U431 ( .A(G176GAT), .B(G92GAT), .ZN(n360) );
  XNOR2_X1 U432 ( .A(n360), .B(G64GAT), .ZN(n423) );
  NAND2_X1 U433 ( .A1(G226GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U434 ( .A(n294), .B(n361), .ZN(n363) );
  XOR2_X1 U435 ( .A(G8GAT), .B(G183GAT), .Z(n396) );
  XNOR2_X1 U436 ( .A(n365), .B(n364), .ZN(n367) );
  XNOR2_X1 U437 ( .A(KEYINPUT27), .B(n548), .ZN(n476) );
  NOR2_X1 U438 ( .A1(n546), .A2(n476), .ZN(n368) );
  XOR2_X1 U439 ( .A(KEYINPUT100), .B(n368), .Z(n484) );
  XOR2_X1 U440 ( .A(KEYINPUT79), .B(KEYINPUT10), .Z(n370) );
  XNOR2_X1 U441 ( .A(G92GAT), .B(KEYINPUT11), .ZN(n369) );
  XNOR2_X1 U442 ( .A(n370), .B(n369), .ZN(n373) );
  INV_X1 U443 ( .A(n373), .ZN(n371) );
  NAND2_X1 U444 ( .A1(n371), .A2(n372), .ZN(n376) );
  INV_X1 U445 ( .A(n372), .ZN(n374) );
  NAND2_X1 U446 ( .A1(n374), .A2(n373), .ZN(n375) );
  NAND2_X1 U447 ( .A1(n376), .A2(n375), .ZN(n379) );
  XNOR2_X1 U448 ( .A(G99GAT), .B(G85GAT), .ZN(n380) );
  XNOR2_X1 U449 ( .A(n380), .B(KEYINPUT78), .ZN(n419) );
  XNOR2_X1 U450 ( .A(n381), .B(n419), .ZN(n382) );
  XNOR2_X1 U451 ( .A(n383), .B(n382), .ZN(n387) );
  XOR2_X1 U452 ( .A(KEYINPUT9), .B(KEYINPUT81), .Z(n385) );
  NAND2_X1 U453 ( .A1(G232GAT), .A2(G233GAT), .ZN(n384) );
  XOR2_X1 U454 ( .A(n385), .B(n384), .Z(n386) );
  XNOR2_X1 U455 ( .A(n387), .B(n386), .ZN(n393) );
  INV_X1 U456 ( .A(KEYINPUT71), .ZN(n391) );
  XOR2_X1 U457 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n389) );
  XNOR2_X1 U458 ( .A(G43GAT), .B(G29GAT), .ZN(n388) );
  XNOR2_X1 U459 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U460 ( .A(n391), .B(n390), .ZN(n443) );
  XNOR2_X1 U461 ( .A(n443), .B(KEYINPUT64), .ZN(n392) );
  INV_X1 U462 ( .A(n574), .ZN(n457) );
  INV_X1 U463 ( .A(KEYINPUT36), .ZN(n394) );
  XNOR2_X1 U464 ( .A(n457), .B(n394), .ZN(n593) );
  XOR2_X1 U465 ( .A(n396), .B(n395), .Z(n398) );
  NAND2_X1 U466 ( .A1(G231GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U467 ( .A(n398), .B(n397), .ZN(n402) );
  XOR2_X1 U468 ( .A(KEYINPUT84), .B(KEYINPUT12), .Z(n400) );
  XNOR2_X1 U469 ( .A(KEYINPUT83), .B(KEYINPUT15), .ZN(n399) );
  XNOR2_X1 U470 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U471 ( .A(n402), .B(n401), .Z(n408) );
  XOR2_X1 U472 ( .A(G64GAT), .B(G78GAT), .Z(n404) );
  XNOR2_X1 U473 ( .A(G1GAT), .B(G211GAT), .ZN(n403) );
  XNOR2_X1 U474 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U475 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U476 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U477 ( .A(n409), .B(KEYINPUT82), .Z(n413) );
  XOR2_X1 U478 ( .A(G57GAT), .B(KEYINPUT13), .Z(n411) );
  XNOR2_X1 U479 ( .A(G71GAT), .B(KEYINPUT75), .ZN(n410) );
  XNOR2_X1 U480 ( .A(n411), .B(n410), .ZN(n422) );
  XNOR2_X1 U481 ( .A(n422), .B(KEYINPUT14), .ZN(n412) );
  NAND2_X1 U482 ( .A1(n593), .A2(n591), .ZN(n415) );
  XOR2_X1 U483 ( .A(KEYINPUT66), .B(KEYINPUT45), .Z(n414) );
  XNOR2_X1 U484 ( .A(n415), .B(n414), .ZN(n427) );
  XOR2_X1 U485 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n421) );
  XOR2_X1 U486 ( .A(KEYINPUT31), .B(G120GAT), .Z(n417) );
  NAND2_X1 U487 ( .A1(G230GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U488 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U489 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U490 ( .A(n295), .B(n422), .ZN(n426) );
  XNOR2_X1 U491 ( .A(n424), .B(n423), .ZN(n425) );
  INV_X1 U492 ( .A(n588), .ZN(n489) );
  NAND2_X1 U493 ( .A1(n427), .A2(n489), .ZN(n429) );
  INV_X1 U494 ( .A(KEYINPUT117), .ZN(n428) );
  XNOR2_X1 U495 ( .A(n429), .B(n428), .ZN(n450) );
  XOR2_X1 U496 ( .A(G197GAT), .B(G15GAT), .Z(n431) );
  XNOR2_X1 U497 ( .A(G169GAT), .B(G113GAT), .ZN(n430) );
  XNOR2_X1 U498 ( .A(n431), .B(n430), .ZN(n433) );
  XOR2_X1 U499 ( .A(G36GAT), .B(G50GAT), .Z(n432) );
  XNOR2_X1 U500 ( .A(n433), .B(n432), .ZN(n447) );
  XOR2_X1 U501 ( .A(KEYINPUT74), .B(G8GAT), .Z(n435) );
  XNOR2_X1 U502 ( .A(G141GAT), .B(G22GAT), .ZN(n434) );
  XNOR2_X1 U503 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U504 ( .A(KEYINPUT70), .B(G1GAT), .Z(n437) );
  XNOR2_X1 U505 ( .A(KEYINPUT73), .B(KEYINPUT68), .ZN(n436) );
  XNOR2_X1 U506 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U507 ( .A(n439), .B(n438), .Z(n445) );
  XOR2_X1 U508 ( .A(KEYINPUT72), .B(KEYINPUT30), .Z(n441) );
  XNOR2_X1 U509 ( .A(KEYINPUT69), .B(KEYINPUT29), .ZN(n440) );
  XNOR2_X1 U510 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U511 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U512 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U513 ( .A(n447), .B(n446), .ZN(n449) );
  NAND2_X1 U514 ( .A1(G229GAT), .A2(G233GAT), .ZN(n448) );
  XOR2_X1 U515 ( .A(n449), .B(n448), .Z(n534) );
  INV_X1 U516 ( .A(n534), .ZN(n583) );
  NOR2_X1 U517 ( .A1(n450), .A2(n583), .ZN(n451) );
  XNOR2_X1 U518 ( .A(KEYINPUT118), .B(n451), .ZN(n462) );
  INV_X1 U519 ( .A(KEYINPUT115), .ZN(n456) );
  INV_X1 U520 ( .A(KEYINPUT41), .ZN(n452) );
  XNOR2_X1 U521 ( .A(n588), .B(n452), .ZN(n567) );
  NAND2_X1 U522 ( .A1(n583), .A2(n567), .ZN(n453) );
  XOR2_X1 U523 ( .A(KEYINPUT46), .B(n453), .Z(n454) );
  XNOR2_X1 U524 ( .A(n456), .B(n455), .ZN(n458) );
  NAND2_X1 U525 ( .A1(n458), .A2(n457), .ZN(n460) );
  XNOR2_X1 U526 ( .A(n465), .B(n464), .ZN(n493) );
  NOR2_X1 U527 ( .A1(n484), .A2(n493), .ZN(n466) );
  NAND2_X1 U528 ( .A1(n553), .A2(n564), .ZN(n467) );
  NAND2_X1 U529 ( .A1(n561), .A2(n574), .ZN(n471) );
  XOR2_X1 U530 ( .A(KEYINPUT121), .B(KEYINPUT51), .Z(n469) );
  XNOR2_X1 U531 ( .A(n471), .B(n470), .ZN(G1343GAT) );
  NOR2_X1 U532 ( .A1(n548), .A2(n550), .ZN(n472) );
  XOR2_X1 U533 ( .A(KEYINPUT25), .B(n473), .Z(n478) );
  XOR2_X1 U534 ( .A(KEYINPUT101), .B(KEYINPUT26), .Z(n475) );
  NAND2_X1 U535 ( .A1(n498), .A2(n550), .ZN(n474) );
  XNOR2_X1 U536 ( .A(n475), .B(n474), .ZN(n582) );
  NOR2_X1 U537 ( .A1(n582), .A2(n476), .ZN(n477) );
  NOR2_X1 U538 ( .A1(n478), .A2(n477), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n480), .B(n479), .ZN(n481) );
  NAND2_X1 U540 ( .A1(n481), .A2(n546), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n482), .B(KEYINPUT103), .ZN(n486) );
  NAND2_X1 U542 ( .A1(n553), .A2(n550), .ZN(n483) );
  NOR2_X1 U543 ( .A1(n484), .A2(n483), .ZN(n485) );
  NOR2_X1 U544 ( .A1(n486), .A2(n485), .ZN(n515) );
  NOR2_X1 U545 ( .A1(n591), .A2(n515), .ZN(n487) );
  NAND2_X1 U546 ( .A1(n487), .A2(n593), .ZN(n488) );
  XOR2_X1 U547 ( .A(KEYINPUT37), .B(n488), .Z(n545) );
  NAND2_X1 U548 ( .A1(n583), .A2(n489), .ZN(n518) );
  NOR2_X1 U549 ( .A1(n545), .A2(n518), .ZN(n490) );
  XOR2_X1 U550 ( .A(KEYINPUT38), .B(n490), .Z(n531) );
  NOR2_X1 U551 ( .A1(n531), .A2(n546), .ZN(n492) );
  XNOR2_X1 U552 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n492), .B(n491), .ZN(G1328GAT) );
  XNOR2_X1 U554 ( .A(KEYINPUT112), .B(n567), .ZN(n558) );
  NOR2_X1 U555 ( .A1(n548), .A2(n493), .ZN(n496) );
  INV_X1 U556 ( .A(KEYINPUT54), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n496), .B(n495), .ZN(n497) );
  NAND2_X1 U558 ( .A1(n497), .A2(n546), .ZN(n581) );
  NOR2_X1 U559 ( .A1(n498), .A2(n581), .ZN(n499) );
  XNOR2_X1 U560 ( .A(n499), .B(KEYINPUT55), .ZN(n500) );
  NAND2_X1 U561 ( .A1(n558), .A2(n578), .ZN(n503) );
  XOR2_X1 U562 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n501) );
  XNOR2_X1 U563 ( .A(n501), .B(G176GAT), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n503), .B(n502), .ZN(G1349GAT) );
  NOR2_X1 U565 ( .A1(n531), .A2(n550), .ZN(n507) );
  XNOR2_X1 U566 ( .A(KEYINPUT40), .B(KEYINPUT110), .ZN(n505) );
  NAND2_X1 U567 ( .A1(n574), .A2(n578), .ZN(n509) );
  XOR2_X1 U568 ( .A(KEYINPUT106), .B(KEYINPUT34), .Z(n511) );
  XNOR2_X1 U569 ( .A(G1GAT), .B(KEYINPUT105), .ZN(n510) );
  XNOR2_X1 U570 ( .A(n511), .B(n510), .ZN(n521) );
  NAND2_X1 U571 ( .A1(n457), .A2(n591), .ZN(n514) );
  XNOR2_X1 U572 ( .A(KEYINPUT16), .B(KEYINPUT86), .ZN(n512) );
  XNOR2_X1 U573 ( .A(n512), .B(KEYINPUT85), .ZN(n513) );
  XNOR2_X1 U574 ( .A(n514), .B(n513), .ZN(n517) );
  INV_X1 U575 ( .A(n515), .ZN(n516) );
  NAND2_X1 U576 ( .A1(n517), .A2(n516), .ZN(n535) );
  NOR2_X1 U577 ( .A1(n518), .A2(n535), .ZN(n519) );
  XOR2_X1 U578 ( .A(KEYINPUT104), .B(n519), .Z(n526) );
  NOR2_X1 U579 ( .A1(n546), .A2(n526), .ZN(n520) );
  XOR2_X1 U580 ( .A(n521), .B(n520), .Z(G1324GAT) );
  XNOR2_X1 U581 ( .A(G8GAT), .B(KEYINPUT107), .ZN(n523) );
  NOR2_X1 U582 ( .A1(n548), .A2(n526), .ZN(n522) );
  XNOR2_X1 U583 ( .A(n523), .B(n522), .ZN(G1325GAT) );
  NOR2_X1 U584 ( .A1(n526), .A2(n550), .ZN(n525) );
  XNOR2_X1 U585 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n524) );
  XNOR2_X1 U586 ( .A(n525), .B(n524), .ZN(G1326GAT) );
  NOR2_X1 U587 ( .A1(n553), .A2(n526), .ZN(n527) );
  XOR2_X1 U588 ( .A(KEYINPUT108), .B(n527), .Z(n528) );
  XNOR2_X1 U589 ( .A(G22GAT), .B(n528), .ZN(G1327GAT) );
  XNOR2_X1 U590 ( .A(G36GAT), .B(KEYINPUT109), .ZN(n530) );
  NOR2_X1 U591 ( .A1(n548), .A2(n531), .ZN(n529) );
  XNOR2_X1 U592 ( .A(n530), .B(n529), .ZN(G1329GAT) );
  XNOR2_X1 U593 ( .A(G50GAT), .B(KEYINPUT111), .ZN(n533) );
  NOR2_X1 U594 ( .A1(n553), .A2(n531), .ZN(n532) );
  XNOR2_X1 U595 ( .A(n533), .B(n532), .ZN(G1331GAT) );
  NAND2_X1 U596 ( .A1(n558), .A2(n534), .ZN(n544) );
  OR2_X1 U597 ( .A1(n535), .A2(n544), .ZN(n540) );
  NOR2_X1 U598 ( .A1(n546), .A2(n540), .ZN(n536) );
  XOR2_X1 U599 ( .A(n536), .B(KEYINPUT42), .Z(n537) );
  XNOR2_X1 U600 ( .A(G57GAT), .B(n537), .ZN(G1332GAT) );
  NOR2_X1 U601 ( .A1(n548), .A2(n540), .ZN(n538) );
  XOR2_X1 U602 ( .A(G64GAT), .B(n538), .Z(G1333GAT) );
  NOR2_X1 U603 ( .A1(n550), .A2(n540), .ZN(n539) );
  XOR2_X1 U604 ( .A(G71GAT), .B(n539), .Z(G1334GAT) );
  NOR2_X1 U605 ( .A1(n553), .A2(n540), .ZN(n542) );
  XNOR2_X1 U606 ( .A(KEYINPUT113), .B(KEYINPUT43), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U608 ( .A(G78GAT), .B(n543), .Z(G1335GAT) );
  OR2_X1 U609 ( .A1(n545), .A2(n544), .ZN(n552) );
  NOR2_X1 U610 ( .A1(n546), .A2(n552), .ZN(n547) );
  XOR2_X1 U611 ( .A(G85GAT), .B(n547), .Z(G1336GAT) );
  NOR2_X1 U612 ( .A1(n548), .A2(n552), .ZN(n549) );
  XOR2_X1 U613 ( .A(G92GAT), .B(n549), .Z(G1337GAT) );
  NOR2_X1 U614 ( .A1(n550), .A2(n552), .ZN(n551) );
  XOR2_X1 U615 ( .A(G99GAT), .B(n551), .Z(G1338GAT) );
  NOR2_X1 U616 ( .A1(n553), .A2(n552), .ZN(n555) );
  XNOR2_X1 U617 ( .A(KEYINPUT114), .B(KEYINPUT44), .ZN(n554) );
  XNOR2_X1 U618 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U619 ( .A(G106GAT), .B(n556), .Z(G1339GAT) );
  NAND2_X1 U620 ( .A1(n583), .A2(n561), .ZN(n557) );
  XNOR2_X1 U621 ( .A(G113GAT), .B(n557), .ZN(G1340GAT) );
  XOR2_X1 U622 ( .A(G120GAT), .B(KEYINPUT49), .Z(n560) );
  NAND2_X1 U623 ( .A1(n561), .A2(n558), .ZN(n559) );
  XNOR2_X1 U624 ( .A(n560), .B(n559), .ZN(G1341GAT) );
  NAND2_X1 U625 ( .A1(n561), .A2(n591), .ZN(n562) );
  XNOR2_X1 U626 ( .A(n562), .B(KEYINPUT50), .ZN(n563) );
  XNOR2_X1 U627 ( .A(G127GAT), .B(n563), .ZN(G1342GAT) );
  INV_X1 U628 ( .A(n564), .ZN(n565) );
  NOR2_X1 U629 ( .A1(n582), .A2(n565), .ZN(n573) );
  NAND2_X1 U630 ( .A1(n583), .A2(n573), .ZN(n566) );
  XNOR2_X1 U631 ( .A(G141GAT), .B(n566), .ZN(G1344GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n569) );
  NAND2_X1 U633 ( .A1(n573), .A2(n567), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(G148GAT), .B(n570), .ZN(G1345GAT) );
  NAND2_X1 U636 ( .A1(n573), .A2(n591), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(KEYINPUT122), .ZN(n572) );
  XNOR2_X1 U638 ( .A(G155GAT), .B(n572), .ZN(G1346GAT) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U641 ( .A(G169GAT), .B(KEYINPUT124), .ZN(n577) );
  NAND2_X1 U642 ( .A1(n583), .A2(n578), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(G1348GAT) );
  XOR2_X1 U644 ( .A(G183GAT), .B(KEYINPUT125), .Z(n580) );
  NAND2_X1 U645 ( .A1(n578), .A2(n591), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(G1350GAT) );
  XNOR2_X1 U647 ( .A(KEYINPUT126), .B(KEYINPUT59), .ZN(n587) );
  XOR2_X1 U648 ( .A(G197GAT), .B(KEYINPUT60), .Z(n585) );
  NOR2_X1 U649 ( .A1(n582), .A2(n581), .ZN(n594) );
  NAND2_X1 U650 ( .A1(n594), .A2(n583), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(G1352GAT) );
  XOR2_X1 U653 ( .A(G204GAT), .B(KEYINPUT61), .Z(n590) );
  NAND2_X1 U654 ( .A1(n594), .A2(n588), .ZN(n589) );
  XNOR2_X1 U655 ( .A(n590), .B(n589), .ZN(G1353GAT) );
  NAND2_X1 U656 ( .A1(n594), .A2(n591), .ZN(n592) );
  XNOR2_X1 U657 ( .A(n592), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U658 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n596) );
  NAND2_X1 U659 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U660 ( .A(n596), .B(n595), .ZN(n597) );
  XNOR2_X1 U661 ( .A(G218GAT), .B(n597), .ZN(G1355GAT) );
endmodule

