//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 1 1 0 1 0 0 1 1 0 0 1 0 0 1 1 1 1 0 0 1 0 1 0 1 0 1 0 0 1 0 1 1 0 0 0 0 1 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:55 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  XOR2_X1   g0009(.A(KEYINPUT64), .B(G77), .Z(new_n210));
  XOR2_X1   g0010(.A(KEYINPUT65), .B(G244), .Z(new_n211));
  AOI22_X1  g0011(.A1(new_n210), .A2(new_n211), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G226), .ZN(new_n213));
  INV_X1    g0013(.A(G107), .ZN(new_n214));
  INV_X1    g0014(.A(G264), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n212), .B1(new_n202), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G58), .ZN(new_n220));
  INV_X1    g0020(.A(G232), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G68), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NOR4_X1   g0025(.A1(new_n216), .A2(new_n219), .A3(new_n222), .A4(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G97), .A2(G257), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n209), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT1), .Z(new_n229));
  NOR2_X1   g0029(.A1(new_n208), .A2(G13), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n230), .B(G250), .C1(G257), .C2(G264), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT0), .Z(new_n232));
  INV_X1    g0032(.A(new_n201), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(G50), .ZN(new_n234));
  INV_X1    g0034(.A(G20), .ZN(new_n235));
  NAND2_X1  g0035(.A1(G1), .A2(G13), .ZN(new_n236));
  NOR3_X1   g0036(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  NOR3_X1   g0037(.A1(new_n229), .A2(new_n232), .A3(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT2), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G250), .B(G257), .Z(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G68), .B(G77), .Z(new_n250));
  XNOR2_X1  g0050(.A(G50), .B(G58), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  NAND2_X1  g0053(.A1(new_n203), .A2(G20), .ZN(new_n254));
  INV_X1    g0054(.A(G150), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n235), .A2(G33), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT8), .B(G58), .ZN(new_n259));
  OAI221_X1 g0059(.A(new_n254), .B1(new_n255), .B2(new_n257), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n236), .B1(new_n208), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G20), .ZN(new_n264));
  INV_X1    g0064(.A(G13), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n260), .A2(new_n262), .B1(new_n202), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT66), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n264), .B(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G50), .ZN(new_n270));
  XOR2_X1   g0070(.A(new_n270), .B(KEYINPUT67), .Z(new_n271));
  NOR2_X1   g0071(.A1(new_n266), .A2(new_n262), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n267), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT9), .ZN(new_n275));
  AND2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n274), .A2(new_n275), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT3), .B(G33), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G222), .A2(G1698), .ZN(new_n279));
  INV_X1    g0079(.A(G1698), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(G223), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n278), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n236), .B1(G33), .B2(G41), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n282), .B(new_n283), .C1(new_n210), .C2(new_n278), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n263), .B1(G41), .B2(G45), .ZN(new_n285));
  INV_X1    g0085(.A(G274), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n283), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n285), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n284), .B(new_n288), .C1(new_n213), .C2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G190), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NOR3_X1   g0093(.A1(new_n276), .A2(new_n277), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT70), .ZN(new_n295));
  AOI21_X1  g0095(.A(KEYINPUT10), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n291), .A2(G200), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n294), .B(new_n297), .C1(new_n295), .C2(KEYINPUT10), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n291), .A2(new_n301), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n291), .A2(G179), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n274), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n299), .A2(new_n300), .A3(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT13), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n221), .A2(G1698), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n278), .B(new_n307), .C1(G226), .C2(G1698), .ZN(new_n308));
  NAND2_X1  g0108(.A1(G33), .A2(G97), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n289), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n310), .A2(new_n287), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n290), .A2(new_n224), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n306), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  NOR4_X1   g0114(.A1(new_n310), .A2(new_n312), .A3(KEYINPUT13), .A4(new_n287), .ZN(new_n315));
  OAI21_X1  g0115(.A(G169), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT14), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n314), .A2(new_n315), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G179), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT14), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n320), .B(G169), .C1(new_n314), .C2(new_n315), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n317), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n223), .A2(G20), .ZN(new_n323));
  INV_X1    g0123(.A(G77), .ZN(new_n324));
  OAI221_X1 g0124(.A(new_n323), .B1(new_n258), .B2(new_n324), .C1(new_n257), .C2(new_n202), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n325), .A2(new_n262), .ZN(new_n326));
  OR2_X1    g0126(.A1(new_n326), .A2(KEYINPUT11), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(KEYINPUT11), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n266), .A2(new_n223), .ZN(new_n329));
  XNOR2_X1  g0129(.A(new_n329), .B(KEYINPUT12), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n269), .A2(new_n272), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G68), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n327), .A2(new_n328), .A3(new_n330), .A4(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n318), .A2(G190), .ZN(new_n334));
  OAI21_X1  g0134(.A(G200), .B1(new_n314), .B2(new_n315), .ZN(new_n335));
  INV_X1    g0135(.A(new_n333), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n322), .A2(new_n333), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n220), .A2(new_n223), .ZN(new_n340));
  OAI21_X1  g0140(.A(G20), .B1(new_n340), .B2(new_n201), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n256), .A2(G159), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT3), .ZN(new_n345));
  OAI21_X1  g0145(.A(KEYINPUT71), .B1(new_n345), .B2(G33), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(G33), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n345), .A2(KEYINPUT71), .A3(G33), .ZN(new_n349));
  AOI21_X1  g0149(.A(G20), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT7), .ZN(new_n351));
  OAI21_X1  g0151(.A(G68), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI211_X1 g0152(.A(KEYINPUT7), .B(G20), .C1(new_n348), .C2(new_n349), .ZN(new_n353));
  OAI211_X1 g0153(.A(KEYINPUT16), .B(new_n344), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT16), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n351), .B1(new_n278), .B2(G20), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n347), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n358), .A2(KEYINPUT7), .A3(new_n235), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n223), .B1(new_n356), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n355), .B1(new_n360), .B2(new_n343), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n354), .A2(new_n262), .A3(new_n361), .ZN(new_n362));
  OR2_X1    g0162(.A1(G223), .A2(G1698), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n213), .A2(G1698), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n348), .A2(new_n349), .A3(new_n363), .A4(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(G33), .A2(G87), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n289), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n288), .B1(new_n290), .B2(new_n221), .ZN(new_n368));
  OAI21_X1  g0168(.A(G200), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n266), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n259), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(new_n331), .B2(new_n259), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n367), .A2(new_n368), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(G190), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n362), .A2(new_n369), .A3(new_n372), .A4(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT72), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT17), .ZN(new_n378));
  OR2_X1    g0178(.A1(new_n377), .A2(KEYINPUT17), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(KEYINPUT17), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n375), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n362), .A2(new_n372), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n373), .A2(G179), .ZN(new_n383));
  OAI21_X1  g0183(.A(G169), .B1(new_n367), .B2(new_n368), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(KEYINPUT18), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n382), .A2(KEYINPUT18), .A3(new_n385), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n378), .B(new_n381), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n224), .A2(G1698), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(G232), .B2(G1698), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n289), .B1(new_n278), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(G107), .B2(new_n278), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n289), .A2(new_n211), .A3(new_n285), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n392), .A2(new_n288), .A3(new_n393), .ZN(new_n394));
  OR2_X1    g0194(.A1(new_n394), .A2(G179), .ZN(new_n395));
  INV_X1    g0195(.A(new_n259), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n396), .A2(new_n256), .B1(new_n210), .B2(G20), .ZN(new_n397));
  XNOR2_X1  g0197(.A(KEYINPUT15), .B(G87), .ZN(new_n398));
  XNOR2_X1  g0198(.A(new_n398), .B(KEYINPUT69), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n397), .B1(new_n399), .B2(new_n258), .ZN(new_n400));
  INV_X1    g0200(.A(new_n210), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n400), .A2(new_n262), .B1(new_n401), .B2(new_n266), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n331), .A2(G77), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n394), .A2(new_n301), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n395), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  OR2_X1    g0207(.A1(new_n388), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n394), .A2(new_n292), .ZN(new_n409));
  XNOR2_X1  g0209(.A(new_n409), .B(KEYINPUT68), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n394), .A2(G200), .ZN(new_n411));
  INV_X1    g0211(.A(new_n404), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NOR4_X1   g0214(.A1(new_n305), .A2(new_n339), .A3(new_n408), .A4(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT22), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n235), .A2(G87), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n416), .B1(new_n358), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n348), .A2(new_n349), .ZN(new_n419));
  OR3_X1    g0219(.A1(new_n419), .A2(new_n416), .A3(new_n417), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT23), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n421), .B1(G20), .B2(new_n214), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n421), .A2(new_n214), .A3(G20), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT81), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n421), .A2(new_n214), .A3(KEYINPUT81), .A4(G20), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n422), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT82), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n235), .A2(G33), .A3(G116), .ZN(new_n429));
  AND3_X1   g0229(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n428), .B1(new_n427), .B2(new_n429), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n418), .B(new_n420), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT24), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n427), .A2(new_n429), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT82), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n438), .A2(KEYINPUT24), .A3(new_n418), .A4(new_n420), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n434), .A2(new_n439), .A3(new_n262), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n272), .B1(G1), .B2(new_n261), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(G107), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n266), .A2(new_n214), .ZN(new_n444));
  XOR2_X1   g0244(.A(new_n444), .B(KEYINPUT25), .Z(new_n445));
  NAND3_X1  g0245(.A1(new_n440), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n218), .A2(new_n280), .ZN(new_n447));
  INV_X1    g0247(.A(G257), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(G1698), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n348), .A2(new_n349), .A3(new_n447), .A4(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G33), .A2(G294), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n289), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n263), .A2(G45), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(KEYINPUT5), .A2(G41), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(KEYINPUT5), .A2(G41), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n454), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n289), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n459), .A2(new_n215), .ZN(new_n460));
  INV_X1    g0260(.A(new_n457), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n453), .B1(new_n461), .B2(new_n455), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G274), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n452), .A2(new_n460), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(KEYINPUT83), .A3(G169), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT83), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n468), .B1(new_n465), .B2(new_n301), .ZN(new_n469));
  INV_X1    g0269(.A(G179), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n467), .B(new_n469), .C1(new_n470), .C2(new_n466), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n446), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n465), .A2(new_n292), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n473), .B1(new_n465), .B2(G200), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n440), .A2(new_n474), .A3(new_n443), .A4(new_n445), .ZN(new_n475));
  AND2_X1   g0275(.A1(new_n475), .A2(KEYINPUT84), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n475), .A2(KEYINPUT84), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n472), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT75), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n462), .A2(new_n283), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n481), .A2(G257), .B1(G274), .B2(new_n462), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G283), .ZN(new_n483));
  AND2_X1   g0283(.A1(G250), .A2(G1698), .ZN(new_n484));
  INV_X1    g0284(.A(G244), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(G1698), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n484), .B1(new_n486), .B2(KEYINPUT4), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n483), .B1(new_n487), .B2(new_n358), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT4), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT71), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n490), .B1(KEYINPUT3), .B2(new_n261), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n349), .B(new_n486), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n488), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  OAI211_X1 g0294(.A(G179), .B(new_n482), .C1(new_n494), .C2(new_n289), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(new_n489), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n280), .A2(G244), .ZN(new_n497));
  OAI22_X1  g0297(.A1(new_n497), .A2(new_n489), .B1(new_n218), .B2(new_n280), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n498), .A2(new_n278), .B1(G33), .B2(G283), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n289), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n463), .B1(new_n459), .B2(new_n448), .ZN(new_n501));
  OAI21_X1  g0301(.A(G169), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n495), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n370), .A2(G97), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n442), .A2(G97), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n214), .B1(new_n356), .B2(new_n359), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n256), .A2(G77), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT6), .ZN(new_n510));
  INV_X1    g0310(.A(G97), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n511), .A2(new_n214), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n510), .B1(new_n512), .B2(new_n205), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n214), .A2(KEYINPUT6), .A3(G97), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n235), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR3_X1   g0315(.A1(new_n507), .A2(new_n509), .A3(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n262), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n505), .B(new_n506), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n503), .A2(KEYINPUT74), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(KEYINPUT74), .B1(new_n503), .B2(new_n518), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT73), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT7), .B1(new_n358), .B2(new_n235), .ZN(new_n524));
  AOI211_X1 g0324(.A(new_n351), .B(G20), .C1(new_n347), .C2(new_n357), .ZN(new_n525));
  OAI21_X1  g0325(.A(G107), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n515), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n526), .A2(new_n527), .A3(new_n508), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n504), .B1(new_n528), .B2(new_n262), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n529), .A2(KEYINPUT73), .A3(new_n506), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n500), .A2(new_n501), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n292), .ZN(new_n532));
  INV_X1    g0332(.A(G200), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n500), .B2(new_n501), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n523), .A2(new_n530), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n480), .B1(new_n521), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n532), .A2(new_n534), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n518), .A2(new_n522), .ZN(new_n538));
  AOI21_X1  g0338(.A(KEYINPUT73), .B1(new_n529), .B2(new_n506), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n540), .B(KEYINPUT75), .C1(new_n520), .C2(new_n519), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n224), .A2(new_n280), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n485), .A2(G1698), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n348), .A2(new_n349), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(G33), .A2(G116), .ZN(new_n545));
  AND3_X1   g0345(.A1(new_n544), .A2(KEYINPUT77), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(KEYINPUT77), .B1(new_n544), .B2(new_n545), .ZN(new_n547));
  NOR3_X1   g0347(.A1(new_n546), .A2(new_n547), .A3(new_n289), .ZN(new_n548));
  OR2_X1    g0348(.A1(new_n454), .A2(KEYINPUT76), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n454), .A2(KEYINPUT76), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n549), .A2(new_n289), .A3(G250), .A4(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n454), .A2(G274), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(G200), .B1(new_n548), .B2(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n348), .A2(new_n235), .A3(G68), .A4(new_n349), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT19), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n235), .B1(new_n309), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(G87), .B2(new_n206), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n556), .B1(new_n258), .B2(new_n511), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n555), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n262), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n399), .A2(new_n266), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n561), .B(new_n562), .C1(new_n217), .C2(new_n441), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n544), .A2(new_n545), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT77), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n544), .A2(KEYINPUT77), .A3(new_n545), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n567), .A2(new_n283), .A3(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n553), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n554), .B(new_n564), .C1(new_n292), .C2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n569), .A2(new_n470), .A3(new_n570), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n561), .B(new_n562), .C1(new_n399), .C2(new_n441), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n548), .A2(new_n553), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n573), .B(new_n574), .C1(new_n575), .C2(G169), .ZN(new_n576));
  AND2_X1   g0376(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n536), .A2(KEYINPUT78), .A3(new_n541), .A4(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT80), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT79), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n448), .A2(new_n280), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n215), .A2(G1698), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n348), .A2(new_n349), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n358), .A2(G303), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n580), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n583), .A2(new_n580), .A3(new_n584), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n586), .A2(new_n283), .A3(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(G270), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n463), .B1(new_n459), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n301), .B1(new_n588), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n587), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n593), .A2(new_n585), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n590), .B1(new_n594), .B2(new_n283), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n592), .A2(KEYINPUT21), .B1(new_n595), .B2(G179), .ZN(new_n596));
  INV_X1    g0396(.A(G116), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n266), .A2(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n483), .B(new_n235), .C1(G33), .C2(new_n511), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n599), .B(new_n262), .C1(new_n235), .C2(G116), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT20), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n600), .A2(new_n601), .ZN(new_n603));
  OAI221_X1 g0403(.A(new_n598), .B1(new_n441), .B2(new_n597), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n579), .B1(new_n596), .B2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT21), .ZN(new_n607));
  NOR3_X1   g0407(.A1(new_n595), .A2(new_n607), .A3(new_n301), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n588), .A2(new_n591), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n609), .A2(new_n470), .ZN(new_n610));
  OAI211_X1 g0410(.A(KEYINPUT80), .B(new_n604), .C1(new_n608), .C2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n592), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n607), .B1(new_n612), .B2(new_n605), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n609), .A2(G200), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n614), .B(new_n605), .C1(new_n292), .C2(new_n609), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n606), .A2(new_n611), .A3(new_n613), .A4(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n536), .A2(new_n577), .A3(new_n541), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT78), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AND4_X1   g0419(.A1(new_n415), .A2(new_n479), .A3(new_n578), .A4(new_n619), .ZN(G372));
  INV_X1    g0420(.A(new_n576), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n577), .A2(new_n521), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n621), .B1(new_n622), .B2(KEYINPUT26), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n571), .A2(new_n292), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n533), .B1(new_n569), .B2(new_n570), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n625), .A2(new_n563), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT85), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n624), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(KEYINPUT85), .B1(new_n625), .B2(new_n563), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n621), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT26), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n523), .A2(new_n530), .A3(new_n503), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(KEYINPUT86), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT86), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n523), .A2(new_n530), .A3(new_n634), .A4(new_n503), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n630), .A2(new_n631), .A3(new_n633), .A4(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n521), .A2(new_n535), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n637), .B(new_n630), .C1(new_n476), .C2(new_n477), .ZN(new_n638));
  INV_X1    g0438(.A(new_n472), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n613), .B1(new_n596), .B2(new_n605), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n623), .B(new_n636), .C1(new_n638), .C2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n415), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n304), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n299), .A2(new_n300), .ZN(new_n645));
  OR2_X1    g0445(.A1(new_n387), .A2(new_n386), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n337), .A2(new_n334), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n322), .A2(new_n333), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n647), .B1(new_n649), .B2(new_n407), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n378), .A2(new_n381), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n646), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n644), .B1(new_n645), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n643), .A2(new_n653), .ZN(G369));
  NAND3_X1  g0454(.A1(new_n606), .A2(new_n611), .A3(new_n613), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n265), .A2(G20), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  OR3_X1    g0457(.A1(new_n657), .A2(KEYINPUT27), .A3(G1), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT27), .B1(new_n657), .B2(G1), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(G213), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g0460(.A(KEYINPUT87), .B(G343), .Z(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n655), .A2(new_n664), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n665), .A2(new_n478), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT88), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n639), .A2(new_n664), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n667), .B1(new_n666), .B2(new_n668), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n446), .A2(new_n663), .ZN(new_n674));
  AOI22_X1  g0474(.A1(new_n479), .A2(new_n674), .B1(new_n639), .B2(new_n663), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n605), .A2(new_n664), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n640), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n616), .B2(new_n676), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(G330), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n673), .A2(new_n681), .ZN(G399));
  NAND3_X1  g0482(.A1(new_n205), .A2(new_n217), .A3(new_n597), .ZN(new_n683));
  XOR2_X1   g0483(.A(new_n683), .B(KEYINPUT89), .Z(new_n684));
  INV_X1    g0484(.A(new_n230), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(G41), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n684), .A2(G1), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(new_n234), .B2(new_n687), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT28), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n572), .A2(new_n576), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n691), .A2(new_n520), .A3(new_n519), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n621), .B1(new_n692), .B2(new_n631), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n626), .A2(new_n627), .ZN(new_n694));
  INV_X1    g0494(.A(new_n624), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(new_n695), .A3(new_n629), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n696), .A2(new_n576), .A3(new_n633), .A4(new_n635), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(KEYINPUT26), .ZN(new_n698));
  AND4_X1   g0498(.A1(new_n472), .A2(new_n606), .A3(new_n611), .A4(new_n613), .ZN(new_n699));
  OAI211_X1 g0499(.A(new_n693), .B(new_n698), .C1(new_n638), .C2(new_n699), .ZN(new_n700));
  AND3_X1   g0500(.A1(new_n700), .A2(KEYINPUT29), .A3(new_n664), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT29), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n642), .A2(new_n664), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(G330), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n619), .A2(new_n479), .A3(new_n578), .A4(new_n664), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n452), .A2(new_n460), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n569), .A2(new_n707), .A3(new_n570), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT90), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n610), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n575), .A2(KEYINPUT90), .A3(new_n707), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n711), .A2(KEYINPUT30), .A3(new_n531), .A4(new_n712), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n712), .A2(new_n610), .A3(new_n531), .A4(new_n710), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT30), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n465), .A2(new_n531), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n717), .A2(new_n609), .A3(new_n470), .A4(new_n571), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n713), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n719), .A2(KEYINPUT31), .A3(new_n663), .ZN(new_n720));
  AOI21_X1  g0520(.A(KEYINPUT31), .B1(new_n719), .B2(new_n663), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n705), .B1(new_n706), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n704), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n690), .B1(new_n724), .B2(G1), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT91), .ZN(G364));
  AOI21_X1  g0526(.A(new_n263), .B1(new_n656), .B2(G45), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n686), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n292), .A2(G200), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(new_n470), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G20), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(new_n511), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n235), .A2(new_n470), .A3(KEYINPUT92), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT92), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n737), .B1(G20), .B2(G179), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(new_n731), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n533), .A2(G190), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI22_X1  g0545(.A1(G58), .A2(new_n742), .B1(new_n745), .B2(G68), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n292), .A2(new_n533), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n739), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G190), .A2(G200), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n740), .A2(new_n751), .ZN(new_n752));
  OAI221_X1 g0552(.A(new_n746), .B1(new_n202), .B2(new_n750), .C1(new_n401), .C2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n235), .A2(G179), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n747), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n217), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n358), .ZN(new_n757));
  AOI211_X1 g0557(.A(new_n735), .B(new_n753), .C1(KEYINPUT94), .C2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n754), .A2(new_n751), .ZN(new_n759));
  OR2_X1    g0559(.A1(new_n759), .A2(KEYINPUT93), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(KEYINPUT93), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G159), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT32), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n743), .A2(new_n754), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G107), .ZN(new_n768));
  OR2_X1    g0568(.A1(new_n757), .A2(KEYINPUT94), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n758), .A2(new_n765), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT95), .ZN(new_n771));
  XNOR2_X1  g0571(.A(KEYINPUT33), .B(G317), .ZN(new_n772));
  AOI22_X1  g0572(.A1(G322), .A2(new_n742), .B1(new_n745), .B2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(G311), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n773), .B1(new_n774), .B2(new_n752), .ZN(new_n775));
  INV_X1    g0575(.A(new_n762), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n776), .A2(G329), .ZN(new_n777));
  INV_X1    g0577(.A(G294), .ZN(new_n778));
  INV_X1    g0578(.A(G303), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n734), .A2(new_n778), .B1(new_n755), .B2(new_n779), .ZN(new_n780));
  NOR4_X1   g0580(.A1(new_n775), .A2(new_n278), .A3(new_n777), .A4(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G283), .ZN(new_n782));
  INV_X1    g0582(.A(G326), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n749), .B(KEYINPUT96), .ZN(new_n784));
  OAI221_X1 g0584(.A(new_n781), .B1(new_n782), .B2(new_n766), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n771), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n236), .B1(G20), .B2(new_n301), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n730), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(G355), .A2(new_n278), .A3(new_n230), .ZN(new_n789));
  INV_X1    g0589(.A(new_n419), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n685), .ZN(new_n791));
  INV_X1    g0591(.A(G45), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n791), .B1(new_n252), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n234), .A2(G45), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n789), .B1(G116), .B2(new_n230), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(G13), .A2(G33), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(G20), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n787), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n798), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n788), .B(new_n800), .C1(new_n678), .C2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n729), .B1(new_n678), .B2(G330), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(G330), .B2(new_n678), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(G396));
  NOR2_X1   g0606(.A1(new_n406), .A2(new_n663), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n413), .B1(new_n412), .B2(new_n664), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n807), .B1(new_n808), .B2(new_n406), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n703), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n642), .A2(new_n664), .A3(new_n809), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(new_n723), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(new_n730), .ZN(new_n815));
  AOI22_X1  g0615(.A1(G143), .A2(new_n742), .B1(new_n745), .B2(G150), .ZN(new_n816));
  INV_X1    g0616(.A(G137), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n816), .B1(new_n817), .B2(new_n750), .C1(new_n763), .C2(new_n752), .ZN(new_n818));
  XOR2_X1   g0618(.A(new_n818), .B(KEYINPUT34), .Z(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(G132), .B2(new_n776), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n766), .A2(new_n223), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n733), .A2(G58), .ZN(new_n823));
  INV_X1    g0623(.A(new_n755), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(G50), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n820), .A2(new_n822), .A3(new_n823), .A4(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n767), .A2(G87), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n358), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n776), .A2(G311), .B1(new_n749), .B2(G303), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n214), .B2(new_n755), .ZN(new_n830));
  INV_X1    g0630(.A(new_n752), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n735), .B(new_n830), .C1(G116), .C2(new_n831), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n832), .B1(new_n782), .B2(new_n744), .C1(new_n778), .C2(new_n741), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n826), .A2(new_n419), .B1(new_n828), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(new_n787), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n787), .A2(new_n796), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n324), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n730), .B1(new_n810), .B2(new_n796), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n835), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n815), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(G384));
  NAND2_X1  g0641(.A1(new_n513), .A2(new_n514), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n597), .B1(new_n842), .B2(KEYINPUT35), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n236), .A2(new_n235), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n843), .B(new_n844), .C1(KEYINPUT35), .C2(new_n842), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT36), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n234), .A2(new_n340), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n847), .A2(new_n401), .B1(G50), .B2(new_n223), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n848), .A2(G1), .A3(new_n265), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(KEYINPUT97), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n706), .A2(new_n722), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n344), .B1(new_n352), .B2(new_n353), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n355), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n854), .A2(new_n262), .A3(new_n354), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n660), .B1(new_n855), .B2(new_n372), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n388), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n385), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n858), .A2(new_n660), .B1(new_n855), .B2(new_n372), .ZN(new_n859));
  OAI21_X1  g0659(.A(KEYINPUT37), .B1(new_n859), .B2(new_n376), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n382), .A2(new_n385), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT101), .ZN(new_n862));
  INV_X1    g0662(.A(new_n660), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n862), .B1(new_n382), .B2(new_n863), .ZN(new_n864));
  AOI211_X1 g0664(.A(KEYINPUT101), .B(new_n660), .C1(new_n362), .C2(new_n372), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n861), .B(new_n375), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n860), .B1(new_n866), .B2(KEYINPUT37), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n857), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT38), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n857), .A2(new_n867), .A3(KEYINPUT38), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n333), .A2(new_n663), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT99), .ZN(new_n874));
  OR2_X1    g0674(.A1(new_n873), .A2(KEYINPUT99), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n648), .A2(new_n647), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(KEYINPUT100), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT100), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n338), .A2(new_n878), .A3(new_n874), .A4(new_n875), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n877), .A2(new_n879), .B1(new_n649), .B2(new_n663), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n852), .A2(new_n809), .A3(new_n872), .A4(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT40), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT104), .ZN(new_n885));
  XOR2_X1   g0685(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n886));
  AOI21_X1  g0686(.A(new_n660), .B1(new_n362), .B2(new_n372), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n887), .B(new_n862), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT37), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n888), .A2(new_n889), .A3(new_n861), .A4(new_n375), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n866), .A2(KEYINPUT37), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n888), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n388), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n886), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n857), .A2(new_n867), .A3(KEYINPUT38), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n885), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n890), .A2(new_n891), .B1(new_n388), .B2(new_n893), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n871), .B(KEYINPUT104), .C1(new_n898), .C2(new_n886), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n810), .B1(new_n706), .B2(new_n722), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n900), .A2(new_n901), .A3(KEYINPUT40), .A4(new_n881), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n884), .A2(G330), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n723), .A2(new_n415), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n905), .B(KEYINPUT105), .Z(new_n906));
  AOI211_X1 g0706(.A(new_n810), .B(new_n880), .C1(new_n706), .C2(new_n722), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n883), .B1(new_n897), .B2(new_n899), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n883), .A2(new_n882), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(new_n415), .A3(new_n852), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT103), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n892), .A2(new_n894), .ZN(new_n913));
  INV_X1    g0713(.A(new_n886), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(KEYINPUT39), .B1(new_n872), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n895), .A2(new_n896), .ZN(new_n917));
  NOR2_X1   g0717(.A1(KEYINPUT103), .A2(KEYINPUT39), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n648), .A2(new_n663), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n646), .A2(new_n863), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n807), .B(KEYINPUT98), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n880), .B1(new_n812), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n923), .B1(new_n926), .B2(new_n872), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n922), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n704), .A2(new_n415), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n653), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n928), .B(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n911), .B(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n656), .A2(new_n263), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n851), .B1(new_n932), .B2(new_n933), .ZN(G367));
  XNOR2_X1  g0734(.A(new_n686), .B(KEYINPUT41), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n675), .A2(new_n665), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n666), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n680), .B1(new_n937), .B2(new_n679), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n724), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n523), .A2(new_n530), .A3(new_n663), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n637), .A2(new_n940), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n632), .A2(new_n664), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n673), .A2(new_n943), .ZN(new_n944));
  XOR2_X1   g0744(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n945));
  XNOR2_X1  g0745(.A(new_n944), .B(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n943), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n672), .A2(new_n947), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT44), .Z(new_n949));
  AOI21_X1  g0749(.A(new_n939), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n724), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n935), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n727), .ZN(new_n953));
  OR3_X1    g0753(.A1(new_n666), .A2(KEYINPUT42), .A3(new_n941), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n947), .A2(new_n472), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n664), .B1(new_n955), .B2(new_n521), .ZN(new_n956));
  OAI21_X1  g0756(.A(KEYINPUT42), .B1(new_n666), .B2(new_n941), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n954), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n630), .B1(new_n564), .B2(new_n664), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n621), .A2(new_n563), .A3(new_n663), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(KEYINPUT43), .Z(new_n962));
  AND2_X1   g0762(.A1(new_n958), .A2(new_n962), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n963), .A2(KEYINPUT106), .ZN(new_n964));
  OR3_X1    g0764(.A1(new_n958), .A2(KEYINPUT43), .A3(new_n961), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(KEYINPUT106), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n681), .A2(new_n947), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n967), .B(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n953), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n762), .A2(new_n817), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n278), .B1(new_n401), .B2(new_n766), .C1(new_n752), .C2(new_n202), .ZN(new_n974));
  AOI211_X1 g0774(.A(new_n973), .B(new_n974), .C1(G58), .C2(new_n824), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n742), .A2(G150), .ZN(new_n976));
  INV_X1    g0776(.A(G143), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n784), .A2(new_n977), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n745), .A2(G159), .B1(G68), .B2(new_n733), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n975), .A2(new_n976), .A3(new_n978), .A4(new_n979), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n744), .A2(new_n778), .B1(new_n214), .B2(new_n734), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n790), .B(new_n981), .C1(G283), .C2(new_n831), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n784), .A2(new_n774), .ZN(new_n983));
  OAI21_X1  g0783(.A(KEYINPUT108), .B1(new_n755), .B2(new_n597), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n741), .A2(new_n779), .B1(KEYINPUT46), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n984), .A2(KEYINPUT46), .B1(G97), .B2(new_n767), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n982), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(KEYINPUT109), .B(G317), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n776), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n980), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT47), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n787), .ZN(new_n993));
  INV_X1    g0793(.A(new_n791), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n799), .B1(new_n230), .B2(new_n399), .C1(new_n994), .C2(new_n245), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n993), .A2(new_n729), .A3(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n961), .A2(new_n801), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n972), .A2(new_n999), .ZN(G387));
  NOR2_X1   g0800(.A1(new_n399), .A2(new_n734), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n790), .B1(new_n744), .B2(new_n259), .C1(new_n750), .C2(new_n763), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n1001), .B(new_n1002), .C1(G150), .C2(new_n776), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n831), .A2(G68), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n210), .A2(new_n824), .B1(new_n767), .B2(G97), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n742), .A2(G50), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n779), .A2(new_n752), .B1(new_n744), .B2(new_n774), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(new_n742), .B2(new_n989), .ZN(new_n1009));
  INV_X1    g0809(.A(G322), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1009), .B1(new_n1010), .B2(new_n784), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT48), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1012), .B1(new_n782), .B2(new_n734), .C1(new_n778), .C2(new_n755), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT49), .Z(new_n1014));
  OAI221_X1 g0814(.A(new_n419), .B1(new_n597), .B2(new_n766), .C1(new_n762), .C2(new_n783), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT111), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1007), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n787), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n684), .B(new_n792), .C1(new_n223), .C2(new_n324), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT110), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n396), .A2(new_n202), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT50), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n791), .B1(new_n792), .B2(new_n242), .C1(new_n1020), .C2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n278), .A2(new_n230), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1023), .B1(G107), .B2(new_n230), .C1(new_n684), .C2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n799), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1018), .A2(new_n729), .A3(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n675), .B2(new_n798), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(new_n728), .B2(new_n938), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n724), .A2(new_n938), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1030), .A2(new_n686), .A3(new_n939), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1029), .A2(new_n1031), .ZN(G393));
  NAND2_X1  g0832(.A1(new_n946), .A2(new_n949), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n680), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n946), .A2(new_n949), .A3(new_n681), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n950), .B1(new_n1036), .B2(new_n939), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n686), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1034), .A2(new_n728), .A3(new_n1035), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n947), .A2(new_n798), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n768), .B1(new_n597), .B2(new_n734), .C1(new_n744), .C2(new_n779), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n742), .A2(G311), .B1(new_n749), .B2(G317), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT52), .Z(new_n1043));
  AOI21_X1  g0843(.A(new_n278), .B1(new_n776), .B2(G322), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1043), .B(new_n1044), .C1(new_n778), .C2(new_n752), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1041), .B(new_n1045), .C1(G283), .C2(new_n824), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n742), .A2(G159), .B1(new_n749), .B2(G150), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT51), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n734), .A2(new_n324), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n827), .B1(new_n762), .B2(new_n977), .C1(new_n202), .C2(new_n744), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n790), .B1(new_n223), .B2(new_n755), .C1(new_n752), .C2(new_n259), .ZN(new_n1051));
  NOR4_X1   g0851(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n787), .B1(new_n1046), .B2(new_n1052), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n799), .B1(new_n511), .B2(new_n230), .C1(new_n994), .C2(new_n249), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1040), .A2(new_n1053), .A3(new_n729), .A4(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1039), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1038), .A2(new_n1057), .ZN(G390));
  NAND3_X1  g0858(.A1(new_n916), .A2(new_n796), .A3(new_n919), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n836), .A2(new_n259), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n755), .A2(new_n255), .ZN(new_n1061));
  XOR2_X1   g0861(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n1062));
  XNOR2_X1  g0862(.A(new_n1061), .B(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n278), .B1(new_n766), .B2(new_n202), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(new_n776), .B2(G125), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT113), .Z(new_n1066));
  XOR2_X1   g0866(.A(KEYINPUT54), .B(G143), .Z(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n817), .A2(new_n744), .B1(new_n752), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(G128), .B2(new_n749), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1066), .B(new_n1070), .C1(new_n763), .C2(new_n734), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n1063), .B(new_n1071), .C1(G132), .C2(new_n742), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1049), .B1(new_n776), .B2(G294), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n511), .B2(new_n752), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n822), .B1(new_n741), .B2(new_n597), .C1(new_n750), .C2(new_n782), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1076), .B(new_n358), .C1(new_n214), .C2(new_n744), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1077), .A2(new_n756), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n787), .B1(new_n1072), .B2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1059), .A2(new_n729), .A3(new_n1060), .A4(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n700), .A2(new_n664), .A3(new_n809), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n925), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n881), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n921), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1083), .A2(new_n900), .A3(new_n1084), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n916), .B(new_n919), .C1(new_n926), .C2(new_n921), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n723), .A2(new_n809), .A3(new_n881), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1085), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1080), .B1(new_n1092), .B2(new_n727), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n812), .A2(new_n925), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n723), .A2(new_n809), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n880), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1094), .B1(new_n1096), .B2(new_n1088), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT112), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n881), .B1(new_n723), .B2(new_n809), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1098), .B1(new_n1089), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1082), .B1(new_n1096), .B2(KEYINPUT112), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1097), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n929), .A2(new_n904), .A3(new_n653), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1091), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1088), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n687), .B1(new_n1104), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(KEYINPUT112), .B1(new_n1096), .B2(new_n1088), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n925), .B(new_n1081), .C1(new_n1099), .C2(new_n1098), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1089), .A2(new_n1099), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n1109), .A2(new_n1110), .B1(new_n1111), .B2(new_n1094), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1103), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n1092), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1093), .B1(new_n1108), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(G378));
  INV_X1    g0917(.A(KEYINPUT57), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n305), .A2(new_n274), .A3(new_n863), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n274), .A2(new_n863), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n299), .A2(new_n300), .A3(new_n304), .A4(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1119), .A2(new_n1121), .A3(new_n1123), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n903), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n928), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n884), .A2(new_n902), .A3(G330), .A4(new_n1130), .ZN(new_n1131));
  AND3_X1   g0931(.A1(new_n1128), .A2(new_n1129), .A3(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1129), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1103), .B1(new_n1107), .B2(new_n1112), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1118), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1130), .B1(new_n909), .B2(G330), .ZN(new_n1137));
  AND4_X1   g0937(.A1(G330), .A2(new_n884), .A3(new_n902), .A4(new_n1130), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n928), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1128), .A2(new_n1129), .A3(new_n1131), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1113), .B1(new_n1102), .B2(new_n1092), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1141), .A2(new_n1142), .A3(KEYINPUT57), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1136), .A2(new_n686), .A3(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n730), .B1(new_n1127), .B2(new_n796), .ZN(new_n1145));
  INV_X1    g0945(.A(G41), .ZN(new_n1146));
  AOI21_X1  g0946(.A(G50), .B1(new_n419), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(G33), .B2(G41), .ZN(new_n1148));
  INV_X1    g0948(.A(G132), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n744), .A2(new_n1149), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n749), .A2(G125), .B1(G150), .B2(new_n733), .ZN(new_n1151));
  XOR2_X1   g0951(.A(new_n1151), .B(KEYINPUT116), .Z(new_n1152));
  AOI211_X1 g0952(.A(new_n1150), .B(new_n1152), .C1(new_n824), .C2(new_n1067), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n742), .A2(G128), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1153), .B(new_n1154), .C1(new_n817), .C2(new_n752), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT59), .ZN(new_n1156));
  AOI211_X1 g0956(.A(G33), .B(G41), .C1(new_n767), .C2(G159), .ZN(new_n1157));
  INV_X1    g0957(.A(G124), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1157), .B1(new_n1158), .B2(new_n762), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1159), .B(KEYINPUT117), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1148), .B1(new_n1156), .B2(new_n1160), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n419), .B(new_n1146), .C1(new_n401), .C2(new_n755), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT115), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n399), .A2(new_n752), .B1(new_n741), .B2(new_n214), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n744), .A2(new_n511), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n734), .A2(new_n223), .B1(new_n220), .B2(new_n766), .ZN(new_n1166));
  NOR4_X1   g0966(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n1167), .B1(new_n597), .B2(new_n750), .C1(new_n782), .C2(new_n762), .ZN(new_n1168));
  XOR2_X1   g0968(.A(new_n1168), .B(KEYINPUT58), .Z(new_n1169));
  OAI21_X1  g0969(.A(new_n787), .B1(new_n1161), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n836), .A2(new_n202), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1145), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT118), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(new_n728), .B2(new_n1141), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1144), .A2(new_n1174), .ZN(G375));
  AOI21_X1  g0975(.A(new_n419), .B1(G50), .B2(new_n733), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(G137), .A2(new_n742), .B1(new_n745), .B2(new_n1067), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n1149), .B2(new_n750), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1176), .B1(new_n255), .B2(new_n752), .C1(new_n1178), .C2(KEYINPUT121), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1178), .A2(KEYINPUT121), .B1(G58), .B2(new_n767), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n763), .B2(new_n755), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1179), .B(new_n1181), .C1(G128), .C2(new_n776), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n214), .A2(new_n752), .B1(new_n744), .B2(new_n597), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1183), .B(KEYINPUT119), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n511), .B2(new_n755), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n358), .B1(new_n750), .B2(new_n778), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1001), .B1(G283), .B2(new_n742), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1186), .B1(new_n1188), .B2(KEYINPUT120), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1189), .B1(KEYINPUT120), .B2(new_n1188), .C1(new_n779), .C2(new_n762), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1185), .B(new_n1190), .C1(G77), .C2(new_n767), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n787), .B1(new_n1182), .B2(new_n1191), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1192), .B(new_n729), .C1(new_n881), .C2(new_n797), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n223), .B2(new_n836), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n1112), .B2(new_n728), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n935), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1195), .B1(new_n1196), .B2(new_n1104), .ZN(G381));
  AOI21_X1  g0997(.A(new_n1056), .B1(new_n1037), .B2(new_n686), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1198), .A2(new_n972), .A3(new_n999), .ZN(new_n1199));
  NOR3_X1   g0999(.A1(new_n1199), .A2(G396), .A3(G393), .ZN(new_n1200));
  OR2_X1    g1000(.A1(G381), .A2(G384), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(G375), .A2(G378), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1200), .A2(new_n1202), .A3(new_n1203), .ZN(G407));
  NAND2_X1  g1004(.A1(new_n662), .A2(G213), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1203), .A2(new_n1206), .ZN(new_n1207));
  OR2_X1    g1007(.A1(new_n1207), .A2(KEYINPUT122), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(KEYINPUT122), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(G407), .A2(new_n1208), .A3(G213), .A4(new_n1209), .ZN(G409));
  AOI21_X1  g1010(.A(KEYINPUT124), .B1(new_n972), .B2(new_n999), .ZN(new_n1211));
  OAI21_X1  g1011(.A(G390), .B1(new_n1211), .B2(KEYINPUT125), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT125), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n970), .B1(new_n727), .B2(new_n952), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1214), .A2(new_n998), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1198), .B(new_n1213), .C1(new_n1215), .C2(KEYINPUT124), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1212), .A2(new_n1216), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(G393), .B(new_n805), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(G387), .B2(KEYINPUT125), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1217), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(G390), .A2(G387), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1221), .A2(new_n1199), .A3(new_n1218), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1220), .A2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1116), .B1(new_n1144), .B2(new_n1174), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1141), .A2(new_n1142), .A3(new_n935), .ZN(new_n1225));
  AND3_X1   g1025(.A1(new_n1116), .A2(new_n1174), .A3(new_n1225), .ZN(new_n1226));
  NOR3_X1   g1026(.A1(new_n1224), .A2(new_n1226), .A3(new_n1206), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT60), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1228), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1102), .A2(KEYINPUT60), .A3(new_n1103), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1229), .A2(new_n1230), .A3(new_n686), .A4(new_n1114), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n1195), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n840), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT63), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1231), .A2(G384), .A3(new_n1195), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  NOR3_X1   g1037(.A1(new_n1234), .A2(new_n1235), .A3(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(KEYINPUT61), .B1(new_n1227), .B2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT123), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n1224), .B2(new_n1226), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1116), .A2(new_n1174), .A3(new_n1225), .ZN(new_n1242));
  XOR2_X1   g1042(.A(new_n1172), .B(KEYINPUT118), .Z(new_n1243));
  NAND2_X1  g1043(.A1(new_n1141), .A2(new_n728), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n687), .B1(new_n1246), .B2(new_n1118), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1245), .B1(new_n1247), .B2(new_n1143), .ZN(new_n1248));
  OAI211_X1 g1048(.A(KEYINPUT123), .B(new_n1242), .C1(new_n1248), .C2(new_n1116), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1241), .A2(new_n1205), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1206), .A2(G2897), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n1234), .B2(new_n1237), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1233), .A2(G2897), .A3(new_n1206), .A4(new_n1236), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1235), .B1(new_n1250), .B2(new_n1254), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1234), .A2(new_n1237), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1241), .A2(new_n1205), .A3(new_n1256), .A4(new_n1249), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1223), .B(new_n1239), .C1(new_n1255), .C2(new_n1258), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1221), .A2(new_n1199), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n1218), .A2(new_n1260), .B1(new_n1217), .B2(new_n1219), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1233), .A2(KEYINPUT62), .A3(new_n1236), .ZN(new_n1262));
  NOR4_X1   g1062(.A1(new_n1224), .A2(new_n1262), .A3(new_n1226), .A4(new_n1206), .ZN(new_n1263));
  XOR2_X1   g1063(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1264));
  AOI21_X1  g1064(.A(new_n1263), .B1(new_n1257), .B2(new_n1264), .ZN(new_n1265));
  XOR2_X1   g1065(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n1266));
  INV_X1    g1066(.A(new_n1254), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1266), .B1(new_n1267), .B2(new_n1227), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1261), .B1(new_n1265), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1259), .A2(new_n1269), .ZN(G405));
  OR2_X1    g1070(.A1(new_n1203), .A2(new_n1224), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1271), .A2(new_n1256), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1271), .A2(new_n1256), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1273), .A2(new_n1261), .A3(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1274), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1223), .B1(new_n1276), .B2(new_n1272), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1275), .A2(new_n1277), .ZN(G402));
endmodule


