//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 0 0 0 0 0 1 0 0 0 0 0 1 1 1 0 1 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 1 1 0 1 0 1 0 0 1 0 0 0 1 0 0 0 0 1 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n578, new_n579, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n630, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1200;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT65), .B(G452), .ZN(G409));
  XNOR2_X1  g003(.A(KEYINPUT66), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT67), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT69), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT69), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(G2105), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n461), .A2(new_n463), .A3(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT70), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT70), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n471), .A2(new_n468), .A3(G2104), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n466), .A2(new_n467), .A3(new_n470), .A4(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G137), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n465), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT71), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT71), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n477), .B(new_n465), .C1(new_n473), .C2(new_n474), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g054(.A(KEYINPUT3), .B(G2104), .ZN(new_n480));
  AOI22_X1  g055(.A1(new_n480), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(new_n467), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n479), .A2(new_n482), .ZN(G160));
  NAND4_X1  g058(.A1(new_n466), .A2(G2105), .A3(new_n470), .A4(new_n472), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n467), .A2(G112), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n473), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n489), .B1(G136), .B2(new_n490), .ZN(new_n491));
  XOR2_X1   g066(.A(new_n491), .B(KEYINPUT72), .Z(G162));
  INV_X1    g067(.A(G126), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n467), .A2(G114), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  OAI22_X1  g070(.A1(new_n484), .A2(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n469), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n499), .A2(new_n467), .A3(G138), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  AND2_X1   g076(.A1(new_n467), .A2(G138), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n466), .A2(new_n470), .A3(new_n472), .A4(new_n502), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n501), .B1(new_n503), .B2(KEYINPUT4), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n496), .A2(new_n504), .ZN(G164));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(KEYINPUT73), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT73), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n510), .A2(KEYINPUT6), .A3(G651), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n506), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G50), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT74), .ZN(new_n514));
  XNOR2_X1  g089(.A(new_n513), .B(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n509), .A2(new_n511), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT5), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(new_n506), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AND3_X1   g095(.A1(new_n516), .A2(KEYINPUT75), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g096(.A(KEYINPUT75), .B1(new_n516), .B2(new_n520), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G88), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n520), .A2(G62), .ZN(new_n525));
  AND2_X1   g100(.A1(G75), .A2(G543), .ZN(new_n526));
  OAI21_X1  g101(.A(G651), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n515), .A2(new_n524), .A3(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XOR2_X1   g105(.A(new_n530), .B(KEYINPUT7), .Z(new_n531));
  XOR2_X1   g106(.A(KEYINPUT78), .B(G89), .Z(new_n532));
  AOI21_X1  g107(.A(new_n531), .B1(new_n523), .B2(new_n532), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n533), .A2(KEYINPUT79), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(KEYINPUT79), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n516), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT77), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n512), .A2(KEYINPUT77), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT76), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n518), .A2(new_n541), .A3(new_n519), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n541), .B1(new_n518), .B2(new_n519), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AND2_X1   g120(.A1(G63), .A2(G651), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n540), .A2(G51), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n534), .A2(new_n535), .A3(new_n547), .ZN(G286));
  INV_X1    g123(.A(G286), .ZN(G168));
  NAND2_X1  g124(.A1(G77), .A2(G543), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n520), .A2(KEYINPUT76), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(new_n542), .ZN(new_n552));
  INV_X1    g127(.A(G64), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n550), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n508), .B1(new_n554), .B2(KEYINPUT80), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n555), .B1(KEYINPUT80), .B2(new_n554), .ZN(new_n556));
  AOI22_X1  g131(.A1(G90), .A2(new_n523), .B1(new_n540), .B2(G52), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(G301));
  INV_X1    g133(.A(G301), .ZN(G171));
  AOI22_X1  g134(.A1(new_n545), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n560), .A2(new_n508), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n512), .B(new_n537), .ZN(new_n563));
  INV_X1    g138(.A(G43), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n516), .A2(new_n520), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT75), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n516), .A2(KEYINPUT75), .A3(new_n520), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(G81), .ZN(new_n570));
  OAI22_X1  g145(.A1(new_n563), .A2(new_n564), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AND2_X1   g146(.A1(new_n571), .A2(KEYINPUT81), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n571), .A2(KEYINPUT81), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n562), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G860), .ZN(G153));
  NAND4_X1  g151(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g152(.A1(G1), .A2(G3), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT8), .ZN(new_n579));
  NAND4_X1  g154(.A1(G319), .A2(G483), .A3(G661), .A4(new_n579), .ZN(G188));
  NAND2_X1  g155(.A1(new_n512), .A2(G53), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT9), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n523), .A2(G91), .ZN(new_n583));
  AND2_X1   g158(.A1(new_n520), .A2(G65), .ZN(new_n584));
  AND2_X1   g159(.A1(G78), .A2(G543), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n582), .A2(new_n583), .A3(new_n586), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n587), .A2(KEYINPUT82), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(KEYINPUT82), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G299));
  INV_X1    g166(.A(G74), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n592), .B1(new_n543), .B2(new_n544), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n593), .A2(G651), .B1(G49), .B2(new_n512), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n567), .A2(G87), .A3(new_n568), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(G288));
  NAND2_X1  g171(.A1(G73), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT83), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n597), .B(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(G61), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n600), .B1(new_n518), .B2(new_n519), .ZN(new_n601));
  OAI21_X1  g176(.A(G651), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n512), .A2(G48), .ZN(new_n603));
  AND2_X1   g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n567), .A2(G86), .A3(new_n568), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(G305));
  AOI22_X1  g181(.A1(G85), .A2(new_n523), .B1(new_n540), .B2(G47), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT84), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n545), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n609), .A2(new_n508), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n608), .A2(new_n610), .ZN(G290));
  NAND2_X1  g186(.A1(G301), .A2(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n523), .A2(G92), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT10), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n563), .A2(KEYINPUT85), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT85), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n540), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n615), .A2(new_n617), .A3(G54), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n520), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT86), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n508), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(new_n620), .B2(new_n619), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n614), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n612), .B1(new_n624), .B2(G868), .ZN(G321));
  XNOR2_X1  g200(.A(G321), .B(KEYINPUT87), .ZN(G284));
  NAND2_X1  g201(.A1(G286), .A2(G868), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(new_n590), .B2(G868), .ZN(G297));
  OAI21_X1  g203(.A(new_n627), .B1(new_n590), .B2(G868), .ZN(G280));
  INV_X1    g204(.A(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n624), .B1(new_n630), .B2(G860), .ZN(G148));
  NAND2_X1  g206(.A1(new_n624), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G868), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(G868), .B2(new_n575), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g210(.A1(new_n464), .A2(new_n480), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT12), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  INV_X1    g213(.A(G2100), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n490), .A2(G135), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n485), .A2(G123), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n467), .A2(G111), .ZN(new_n643));
  OAI21_X1  g218(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n641), .B(new_n642), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT88), .B(G2096), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n640), .A2(new_n647), .ZN(G156));
  INV_X1    g223(.A(KEYINPUT14), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2427), .B(G2438), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2430), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT15), .B(G2435), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n649), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(new_n652), .B2(new_n651), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2451), .B(G2454), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT16), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n654), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2443), .B(G2446), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  AND3_X1   g237(.A1(new_n661), .A2(G14), .A3(new_n662), .ZN(G401));
  INV_X1    g238(.A(KEYINPUT18), .ZN(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(KEYINPUT17), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n665), .A2(new_n666), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n664), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(new_n639), .ZN(new_n671));
  XOR2_X1   g246(.A(G2072), .B(G2078), .Z(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(new_n667), .B2(KEYINPUT18), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(G2096), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n671), .B(new_n674), .ZN(G227));
  XNOR2_X1  g250(.A(G1956), .B(G2474), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT89), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1961), .B(G1966), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT20), .Z(new_n684));
  NOR2_X1   g259(.A1(new_n677), .A2(new_n679), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n686), .A2(new_n682), .A3(new_n680), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n684), .B(new_n687), .C1(new_n682), .C2(new_n686), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1991), .B(G1996), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1981), .B(G1986), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(G229));
  NOR2_X1   g269(.A1(G4), .A2(G16), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT94), .ZN(new_n696));
  INV_X1    g271(.A(new_n624), .ZN(new_n697));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(G1348), .Z(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(G5), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(G171), .B2(new_n698), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n702), .A2(G1961), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT24), .ZN(new_n704));
  INV_X1    g279(.A(G34), .ZN(new_n705));
  AOI21_X1  g280(.A(G29), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(new_n704), .B2(new_n705), .ZN(new_n707));
  INV_X1    g282(.A(G29), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(G160), .B2(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n703), .B1(G2084), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G2084), .B2(new_n709), .ZN(new_n711));
  NOR2_X1   g286(.A1(G29), .A2(G35), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(G162), .B2(G29), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT29), .Z(new_n714));
  INV_X1    g289(.A(G2090), .ZN(new_n715));
  AOI211_X1 g290(.A(new_n700), .B(new_n711), .C1(new_n714), .C2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n708), .A2(G33), .ZN(new_n717));
  AOI22_X1  g292(.A1(new_n480), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT96), .ZN(new_n719));
  OAI21_X1  g294(.A(G2105), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n719), .B2(new_n718), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT25), .Z(new_n723));
  INV_X1    g298(.A(G139), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n473), .B2(new_n724), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n717), .B1(new_n727), .B2(new_n708), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n728), .A2(G2072), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT97), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT30), .B(G28), .ZN(new_n731));
  OR2_X1    g306(.A1(KEYINPUT31), .A2(G11), .ZN(new_n732));
  NAND2_X1  g307(.A1(KEYINPUT31), .A2(G11), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n731), .A2(new_n708), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n645), .B2(new_n708), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n735), .A2(KEYINPUT99), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n735), .A2(KEYINPUT99), .ZN(new_n737));
  AOI211_X1 g312(.A(new_n736), .B(new_n737), .C1(new_n728), .C2(G2072), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n708), .A2(G26), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT28), .ZN(new_n740));
  OR2_X1    g315(.A1(G104), .A2(G2105), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n741), .B(G2104), .C1(G116), .C2(new_n467), .ZN(new_n742));
  INV_X1    g317(.A(G140), .ZN(new_n743));
  INV_X1    g318(.A(G128), .ZN(new_n744));
  OAI221_X1 g319(.A(new_n742), .B1(new_n473), .B2(new_n743), .C1(new_n744), .C2(new_n484), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n740), .B1(new_n746), .B2(new_n708), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G2067), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n708), .A2(G27), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G164), .B2(new_n708), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G2078), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n702), .A2(G1961), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n730), .A2(new_n738), .A3(new_n752), .A4(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(G168), .A2(new_n698), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n698), .B2(G21), .ZN(new_n756));
  INV_X1    g331(.A(G1966), .ZN(new_n757));
  AND2_X1   g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(G16), .A2(G19), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n575), .B2(G16), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT95), .B(G1341), .Z(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(G29), .A2(G32), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n490), .A2(G141), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n485), .A2(G129), .ZN(new_n765));
  NAND3_X1  g340(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT26), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n766), .A2(new_n767), .ZN(new_n769));
  AOI22_X1  g344(.A1(G105), .A2(new_n464), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n764), .A2(new_n765), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n771), .A2(KEYINPUT98), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT98), .ZN(new_n773));
  NAND4_X1  g348(.A1(new_n764), .A2(new_n765), .A3(new_n773), .A4(new_n770), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n763), .B1(new_n776), .B2(G29), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT27), .B(G1996), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n756), .B2(new_n757), .ZN(new_n780));
  NOR4_X1   g355(.A1(new_n754), .A2(new_n758), .A3(new_n762), .A4(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT101), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n698), .A2(G20), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT23), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n590), .B2(new_n698), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT100), .ZN(new_n786));
  INV_X1    g361(.A(G1956), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n786), .A2(new_n787), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n788), .B(new_n789), .C1(new_n714), .C2(new_n715), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n716), .B(new_n781), .C1(new_n782), .C2(new_n790), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n790), .A2(new_n782), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n698), .A2(G22), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G166), .B2(new_n698), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT92), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1971), .ZN(new_n798));
  MUX2_X1   g373(.A(G6), .B(G305), .S(G16), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT32), .ZN(new_n800));
  INV_X1    g375(.A(G1981), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(G16), .A2(G23), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT91), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n512), .A2(G49), .ZN(new_n805));
  AOI21_X1  g380(.A(G74), .B1(new_n551), .B2(new_n542), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n805), .B1(new_n806), .B2(new_n508), .ZN(new_n807));
  INV_X1    g382(.A(G87), .ZN(new_n808));
  NOR3_X1   g383(.A1(new_n521), .A2(new_n522), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n804), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n594), .A2(KEYINPUT91), .A3(new_n595), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n803), .B1(new_n812), .B2(G16), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT33), .B(G1976), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n802), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n798), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT34), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT93), .ZN(new_n820));
  INV_X1    g395(.A(G290), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G16), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G16), .B2(G24), .ZN(new_n823));
  INV_X1    g398(.A(G1986), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  NOR2_X1   g401(.A1(G25), .A2(G29), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n490), .A2(G131), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n485), .A2(G119), .ZN(new_n829));
  OR2_X1    g404(.A1(G95), .A2(G2105), .ZN(new_n830));
  OAI211_X1 g405(.A(new_n830), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n828), .A2(new_n829), .A3(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n827), .B1(new_n833), .B2(G29), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT90), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT35), .B(G1991), .Z(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n826), .A2(new_n837), .ZN(new_n838));
  AOI211_X1 g413(.A(new_n825), .B(new_n838), .C1(new_n817), .C2(new_n818), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n820), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(KEYINPUT36), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT36), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n820), .A2(new_n842), .A3(new_n839), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n794), .B1(new_n841), .B2(new_n843), .ZN(G311));
  INV_X1    g419(.A(new_n843), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n842), .B1(new_n820), .B2(new_n839), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n793), .B1(new_n845), .B2(new_n846), .ZN(G150));
  NAND2_X1  g422(.A1(new_n624), .A2(G559), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT38), .ZN(new_n849));
  AOI22_X1  g424(.A1(new_n545), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n850), .A2(new_n508), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n540), .A2(G55), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n523), .A2(G93), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n574), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n854), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n856), .B(new_n562), .C1(new_n572), .C2(new_n573), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n849), .B(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT39), .ZN(new_n860));
  AOI21_X1  g435(.A(G860), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(new_n860), .B2(new_n859), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n854), .A2(G860), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(KEYINPUT37), .Z(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(KEYINPUT102), .Z(G145));
  XOR2_X1   g441(.A(G164), .B(new_n745), .Z(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n727), .B1(new_n868), .B2(new_n771), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n869), .B1(new_n771), .B2(new_n868), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT104), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n776), .A2(KEYINPUT103), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT103), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n775), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(new_n867), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n872), .A2(new_n868), .A3(new_n874), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n871), .B1(new_n878), .B2(new_n727), .ZN(new_n879));
  AOI211_X1 g454(.A(KEYINPUT104), .B(new_n726), .C1(new_n876), .C2(new_n877), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n870), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n485), .A2(G130), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n467), .A2(G118), .ZN(new_n883));
  OAI21_X1  g458(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n885), .B1(G142), .B2(new_n490), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n637), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n832), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n881), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT105), .ZN(new_n890));
  INV_X1    g465(.A(new_n888), .ZN(new_n891));
  OAI211_X1 g466(.A(new_n891), .B(new_n870), .C1(new_n879), .C2(new_n880), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n889), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(G160), .B(new_n645), .ZN(new_n894));
  XNOR2_X1  g469(.A(G162), .B(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n881), .A2(KEYINPUT105), .A3(new_n888), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n893), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n895), .B1(new_n881), .B2(new_n888), .ZN(new_n898));
  AOI21_X1  g473(.A(G37), .B1(new_n898), .B2(new_n892), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g476(.A(new_n858), .B(new_n632), .ZN(new_n902));
  AOI21_X1  g477(.A(KEYINPUT106), .B1(new_n588), .B2(new_n589), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n903), .A2(new_n697), .ZN(new_n904));
  NAND2_X1  g479(.A1(G299), .A2(KEYINPUT106), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(G299), .A2(KEYINPUT106), .A3(new_n697), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n902), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT41), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n906), .A2(KEYINPUT41), .A3(new_n907), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n909), .B1(new_n913), .B2(new_n902), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT42), .ZN(new_n915));
  XNOR2_X1  g490(.A(G290), .B(G305), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n812), .B(G303), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n916), .B(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT42), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n919), .B(new_n909), .C1(new_n913), .C2(new_n902), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n915), .A2(new_n918), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n918), .B1(new_n915), .B2(new_n920), .ZN(new_n922));
  OAI21_X1  g497(.A(G868), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n923), .B1(G868), .B2(new_n856), .ZN(G295));
  OAI21_X1  g499(.A(new_n923), .B1(G868), .B2(new_n856), .ZN(G331));
  INV_X1    g500(.A(KEYINPUT107), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n855), .A2(new_n857), .A3(G301), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(G301), .B1(new_n855), .B2(new_n857), .ZN(new_n929));
  OAI21_X1  g504(.A(G286), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n858), .A2(G171), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n931), .A2(G168), .A3(new_n927), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n911), .A2(new_n930), .A3(new_n912), .A4(new_n932), .ZN(new_n933));
  NOR3_X1   g508(.A1(new_n928), .A2(new_n929), .A3(G286), .ZN(new_n934));
  AOI21_X1  g509(.A(G168), .B1(new_n931), .B2(new_n927), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n907), .B(new_n906), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(new_n918), .ZN(new_n938));
  INV_X1    g513(.A(G37), .ZN(new_n939));
  INV_X1    g514(.A(new_n918), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n936), .A2(new_n933), .A3(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n938), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n926), .B1(new_n942), .B2(KEYINPUT43), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n944));
  AOI21_X1  g519(.A(G37), .B1(new_n937), .B2(new_n918), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n945), .A2(new_n946), .A3(new_n941), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n946), .B1(new_n945), .B2(new_n941), .ZN(new_n949));
  OAI22_X1  g524(.A1(new_n943), .A2(new_n944), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n949), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n951), .A2(new_n947), .A3(new_n926), .A4(KEYINPUT44), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(G397));
  INV_X1    g528(.A(G1384), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n954), .B1(new_n496), .B2(new_n504), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT45), .ZN(new_n958));
  OAI211_X1 g533(.A(KEYINPUT108), .B(new_n954), .C1(new_n496), .C2(new_n504), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G40), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n482), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n476), .A2(new_n478), .A3(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  OR3_X1    g540(.A1(new_n965), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT46), .B1(new_n965), .B2(G1996), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n745), .B(G2067), .ZN(new_n968));
  OR2_X1    g543(.A1(new_n968), .A2(new_n771), .ZN(new_n969));
  AOI22_X1  g544(.A1(new_n966), .A2(new_n967), .B1(new_n964), .B2(new_n969), .ZN(new_n970));
  XOR2_X1   g545(.A(new_n970), .B(KEYINPUT47), .Z(new_n971));
  NAND2_X1  g546(.A1(new_n821), .A2(new_n824), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n972), .B(KEYINPUT109), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n964), .ZN(new_n974));
  XOR2_X1   g549(.A(new_n974), .B(KEYINPUT48), .Z(new_n975));
  NAND2_X1  g550(.A1(new_n964), .A2(new_n968), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n976), .A2(KEYINPUT110), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n976), .A2(KEYINPUT110), .ZN(new_n978));
  INV_X1    g553(.A(G1996), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n771), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n980), .B1(new_n775), .B2(new_n979), .ZN(new_n981));
  AOI211_X1 g556(.A(new_n977), .B(new_n978), .C1(new_n964), .C2(new_n981), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n833), .A2(new_n836), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n833), .A2(new_n836), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n964), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n982), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n971), .B1(new_n975), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G2067), .ZN(new_n988));
  AOI22_X1  g563(.A1(new_n982), .A2(new_n983), .B1(new_n988), .B2(new_n746), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n965), .B1(new_n989), .B2(KEYINPUT127), .ZN(new_n990));
  OR2_X1    g565(.A1(new_n989), .A2(KEYINPUT127), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n987), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n476), .A2(new_n478), .A3(new_n962), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n955), .A2(KEYINPUT50), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n993), .A2(new_n994), .A3(KEYINPUT118), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT50), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n996), .B(new_n954), .C1(new_n496), .C2(new_n504), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT118), .B1(new_n993), .B2(new_n994), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n787), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  XOR2_X1   g575(.A(new_n587), .B(KEYINPUT57), .Z(new_n1001));
  NAND2_X1  g576(.A1(new_n955), .A2(new_n958), .ZN(new_n1002));
  OAI211_X1 g577(.A(KEYINPUT45), .B(new_n954), .C1(new_n496), .C2(new_n504), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n993), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g579(.A(KEYINPUT56), .B(G2072), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1000), .A2(new_n1001), .A3(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n963), .A2(new_n955), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(new_n988), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n994), .A2(new_n1012), .A3(new_n997), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n955), .A2(KEYINPUT113), .A3(KEYINPUT50), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n963), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1011), .B1(new_n1015), .B2(G1348), .ZN(new_n1016));
  AND2_X1   g591(.A1(new_n1016), .A2(new_n624), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1001), .B1(new_n1000), .B2(new_n1008), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1009), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT120), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  OAI211_X1 g596(.A(KEYINPUT120), .B(new_n1009), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT61), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n1000), .A2(new_n1001), .A3(new_n1008), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1023), .B1(new_n1024), .B2(new_n1018), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT60), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1026), .B1(new_n614), .B2(new_n623), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1011), .B(new_n1027), .C1(new_n1015), .C2(G1348), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n624), .A2(KEYINPUT60), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n1028), .B(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1001), .ZN(new_n1031));
  INV_X1    g606(.A(new_n997), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n963), .B1(KEYINPUT50), .B2(new_n955), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1032), .B1(new_n1033), .B2(KEYINPUT118), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n993), .A2(new_n994), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT118), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(G1956), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1031), .B1(new_n1038), .B2(new_n1007), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1039), .A2(KEYINPUT61), .A3(new_n1009), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1025), .A2(new_n1030), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT59), .ZN(new_n1042));
  XOR2_X1   g617(.A(KEYINPUT58), .B(G1341), .Z(new_n1043));
  OAI21_X1  g618(.A(new_n1043), .B1(new_n963), .B2(new_n955), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT121), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n993), .A2(new_n1002), .A3(new_n979), .A4(new_n1003), .ZN(new_n1047));
  OAI211_X1 g622(.A(KEYINPUT121), .B(new_n1043), .C1(new_n963), .C2(new_n955), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT122), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT122), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1046), .A2(new_n1051), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1042), .B1(new_n1053), .B2(new_n575), .ZN(new_n1054));
  AOI211_X1 g629(.A(KEYINPUT59), .B(new_n574), .C1(new_n1050), .C2(new_n1052), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1021), .B(new_n1022), .C1(new_n1041), .C2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT51), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1059));
  INV_X1    g634(.A(G2084), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1059), .A2(new_n1060), .A3(new_n993), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT123), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1004), .A2(new_n757), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1062), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1065));
  OAI21_X1  g640(.A(G8), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(G286), .A2(G8), .ZN(new_n1067));
  XNOR2_X1  g642(.A(new_n1067), .B(KEYINPUT124), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1058), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G8), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1070), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1067), .ZN(new_n1072));
  NOR3_X1   g647(.A1(new_n1071), .A2(new_n1072), .A3(KEYINPUT51), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1074));
  OAI22_X1  g649(.A1(new_n1069), .A2(new_n1073), .B1(new_n1074), .B2(new_n1067), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1015), .A2(G1961), .ZN(new_n1076));
  INV_X1    g651(.A(G2078), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n993), .A2(new_n1002), .A3(new_n1077), .A4(new_n1003), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1079), .A2(G2078), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n476), .A2(new_n962), .A3(new_n478), .A4(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n494), .A2(new_n495), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1083), .B1(new_n485), .B2(G126), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n503), .A2(KEYINPUT4), .ZN(new_n1085));
  INV_X1    g660(.A(new_n501), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(G1384), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1082), .B1(KEYINPUT45), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n960), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1080), .A2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(G171), .B1(new_n1076), .B2(new_n1091), .ZN(new_n1092));
  AOI22_X1  g667(.A1(new_n1079), .A2(new_n1078), .B1(new_n1089), .B2(new_n1002), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1093), .B(G301), .C1(G1961), .C2(new_n1015), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1092), .A2(KEYINPUT54), .A3(new_n1094), .ZN(new_n1095));
  XNOR2_X1  g670(.A(KEYINPUT114), .B(G2090), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1037), .A2(new_n997), .A3(new_n995), .A4(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT112), .B(G1971), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1004), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(G8), .ZN(new_n1101));
  AND3_X1   g676(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT115), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1106), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1107));
  NAND2_X1  g682(.A1(G303), .A2(G8), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT55), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1110), .A2(KEYINPUT115), .A3(new_n1111), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1107), .A2(new_n1112), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1015), .A2(new_n1096), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n1004), .A2(new_n1098), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1113), .B(G8), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(G86), .ZN(new_n1117));
  NOR3_X1   g692(.A1(new_n521), .A2(new_n522), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(G48), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n602), .B1(new_n1119), .B2(new_n536), .ZN(new_n1120));
  OAI21_X1  g695(.A(G1981), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n604), .A2(new_n605), .A3(new_n801), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1121), .A2(KEYINPUT49), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT116), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1121), .A2(new_n1122), .A3(KEYINPUT116), .A4(KEYINPUT49), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(G8), .B1(new_n963), .B2(new_n955), .ZN(new_n1128));
  AOI21_X1  g703(.A(KEYINPUT49), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1088), .A2(new_n476), .A3(new_n478), .A4(new_n962), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n810), .A2(new_n811), .A3(G1976), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1131), .A2(new_n1132), .A3(G8), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n1127), .A2(new_n1130), .B1(new_n1133), .B2(KEYINPUT52), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1128), .ZN(new_n1135));
  INV_X1    g710(.A(G1976), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT52), .B1(G288), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1135), .A2(new_n1137), .A3(new_n1132), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1134), .A2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1095), .A2(new_n1105), .A3(new_n1116), .A4(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT54), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1089), .A2(new_n1002), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1080), .A2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(G171), .B1(new_n1076), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT125), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  OAI211_X1 g721(.A(KEYINPUT125), .B(G171), .C1(new_n1076), .C2(new_n1143), .ZN(new_n1147));
  OR2_X1    g722(.A1(new_n1076), .A2(new_n1091), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1146), .B(new_n1147), .C1(G171), .C2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1140), .B1(new_n1141), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1057), .A2(new_n1075), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1115), .B1(new_n1015), .B2(new_n1096), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1107), .A2(new_n1112), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1152), .A2(new_n1070), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT117), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1155), .B1(new_n1134), .B2(new_n1138), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1127), .A2(new_n1130), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1133), .A2(KEYINPUT52), .ZN(new_n1158));
  AND4_X1   g733(.A1(new_n1155), .A2(new_n1157), .A3(new_n1138), .A4(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1154), .B1(new_n1156), .B2(new_n1159), .ZN(new_n1160));
  AOI211_X1 g735(.A(G1976), .B(G288), .C1(new_n1127), .C2(new_n1130), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1122), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1135), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1104), .B1(new_n1152), .B2(new_n1070), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1165), .B1(new_n1159), .B2(new_n1156), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT119), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1165), .B(KEYINPUT119), .C1(new_n1156), .C2(new_n1159), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1071), .A2(G168), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT63), .ZN(new_n1171));
  NOR3_X1   g746(.A1(new_n1154), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1168), .A2(new_n1169), .A3(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1105), .A2(new_n1116), .A3(new_n1139), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1171), .B1(new_n1174), .B2(new_n1170), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1164), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  AND3_X1   g751(.A1(new_n1151), .A2(KEYINPUT126), .A3(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(KEYINPUT126), .B1(new_n1151), .B2(new_n1176), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1174), .B1(new_n1147), .B2(new_n1146), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1074), .A2(new_n1067), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(KEYINPUT123), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1070), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1068), .ZN(new_n1185));
  OAI21_X1  g760(.A(KEYINPUT51), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1073), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1180), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT62), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1179), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1075), .A2(KEYINPUT62), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NOR3_X1   g767(.A1(new_n1177), .A2(new_n1178), .A3(new_n1192), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n821), .A2(new_n824), .ZN(new_n1194));
  OR2_X1    g769(.A1(new_n973), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n986), .B1(new_n1195), .B2(new_n964), .ZN(new_n1196));
  XOR2_X1   g771(.A(new_n1196), .B(KEYINPUT111), .Z(new_n1197));
  OAI21_X1  g772(.A(new_n992), .B1(new_n1193), .B2(new_n1197), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g773(.A1(G229), .A2(new_n458), .A3(G401), .A4(G227), .ZN(new_n1200));
  OAI211_X1 g774(.A(new_n900), .B(new_n1200), .C1(new_n948), .C2(new_n949), .ZN(G225));
  INV_X1    g775(.A(G225), .ZN(G308));
endmodule


